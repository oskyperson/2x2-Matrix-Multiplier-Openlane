magic
tech sky130A
magscale 1 2
timestamp 1747094377
<< viali >>
rect 20269 43401 20303 43435
rect 20821 43401 20855 43435
rect 21557 43401 21591 43435
rect 22753 43401 22787 43435
rect 24041 43401 24075 43435
rect 20085 43265 20119 43299
rect 21005 43265 21039 43299
rect 21097 43265 21131 43299
rect 21281 43265 21315 43299
rect 21373 43265 21407 43299
rect 22937 43265 22971 43299
rect 24225 43265 24259 43299
rect 26433 43197 26467 43231
rect 34345 43197 34379 43231
rect 21189 43061 21223 43095
rect 25881 43061 25915 43095
rect 33793 43061 33827 43095
rect 32400 42857 32434 42891
rect 33885 42857 33919 42891
rect 19901 42721 19935 42755
rect 20637 42721 20671 42755
rect 25789 42721 25823 42755
rect 26617 42721 26651 42755
rect 27077 42721 27111 42755
rect 29561 42721 29595 42755
rect 31309 42721 31343 42755
rect 31953 42721 31987 42755
rect 19717 42653 19751 42687
rect 20453 42653 20487 42687
rect 20913 42653 20947 42687
rect 21465 42653 21499 42687
rect 21741 42653 21775 42687
rect 24225 42653 24259 42687
rect 25605 42653 25639 42687
rect 32137 42653 32171 42687
rect 33977 42653 34011 42687
rect 34713 42653 34747 42687
rect 22017 42585 22051 42619
rect 23581 42585 23615 42619
rect 27353 42585 27387 42619
rect 29837 42585 29871 42619
rect 34069 42585 34103 42619
rect 34253 42585 34287 42619
rect 19257 42517 19291 42551
rect 19625 42517 19659 42551
rect 20085 42517 20119 42551
rect 20545 42517 20579 42551
rect 23489 42517 23523 42551
rect 25237 42517 25271 42551
rect 25697 42517 25731 42551
rect 26065 42517 26099 42551
rect 26433 42517 26467 42551
rect 26525 42517 26559 42551
rect 28825 42517 28859 42551
rect 31401 42517 31435 42551
rect 33977 42517 34011 42551
rect 35357 42517 35391 42551
rect 21189 42313 21223 42347
rect 26065 42313 26099 42347
rect 26801 42313 26835 42347
rect 27629 42313 27663 42347
rect 29929 42313 29963 42347
rect 30297 42313 30331 42347
rect 33149 42313 33183 42347
rect 33517 42313 33551 42347
rect 33977 42313 34011 42347
rect 19717 42245 19751 42279
rect 21281 42245 21315 42279
rect 24593 42245 24627 42279
rect 31125 42245 31159 42279
rect 32965 42245 32999 42279
rect 19441 42177 19475 42211
rect 21465 42177 21499 42211
rect 22201 42177 22235 42211
rect 24317 42177 24351 42211
rect 26985 42177 27019 42211
rect 27169 42177 27203 42211
rect 27997 42177 28031 42211
rect 28457 42177 28491 42211
rect 29009 42177 29043 42211
rect 30941 42177 30975 42211
rect 31217 42177 31251 42211
rect 31401 42177 31435 42211
rect 31493 42177 31527 42211
rect 31585 42177 31619 42211
rect 31769 42177 31803 42211
rect 32873 42177 32907 42211
rect 33057 42177 33091 42211
rect 22477 42109 22511 42143
rect 26249 42109 26283 42143
rect 28089 42109 28123 42143
rect 28181 42109 28215 42143
rect 30389 42109 30423 42143
rect 30481 42109 30515 42143
rect 30757 42109 30791 42143
rect 33609 42109 33643 42143
rect 33701 42109 33735 42143
rect 35449 42109 35483 42143
rect 35725 42109 35759 42143
rect 38301 42109 38335 42143
rect 38853 42109 38887 42143
rect 21649 41973 21683 42007
rect 23949 41973 23983 42007
rect 27077 41973 27111 42007
rect 31217 41973 31251 42007
rect 31677 41973 31711 42007
rect 37749 41973 37783 42007
rect 39497 41973 39531 42007
rect 21097 41769 21131 41803
rect 22661 41769 22695 41803
rect 26525 41769 26559 41803
rect 31493 41769 31527 41803
rect 34069 41769 34103 41803
rect 34713 41769 34747 41803
rect 24685 41701 24719 41735
rect 28457 41701 28491 41735
rect 31585 41701 31619 41735
rect 34437 41701 34471 41735
rect 16865 41633 16899 41667
rect 19533 41633 19567 41667
rect 21005 41633 21039 41667
rect 23213 41633 23247 41667
rect 24041 41633 24075 41667
rect 24777 41633 24811 41667
rect 25053 41633 25087 41667
rect 29745 41633 29779 41667
rect 33057 41633 33091 41667
rect 33149 41633 33183 41667
rect 35357 41633 35391 41667
rect 39681 41633 39715 41667
rect 19257 41565 19291 41599
rect 21649 41565 21683 41599
rect 21833 41565 21867 41599
rect 21925 41565 21959 41599
rect 22569 41565 22603 41599
rect 23029 41565 23063 41599
rect 24409 41565 24443 41599
rect 24685 41565 24719 41599
rect 26985 41565 27019 41599
rect 28181 41565 28215 41599
rect 28549 41565 28583 41599
rect 28825 41565 28859 41599
rect 29009 41565 29043 41599
rect 31585 41565 31619 41599
rect 31677 41565 31711 41599
rect 31861 41565 31895 41599
rect 32965 41565 32999 41599
rect 33241 41565 33275 41599
rect 33701 41565 33735 41599
rect 34161 41565 34195 41599
rect 34253 41565 34287 41599
rect 37473 41565 37507 41599
rect 17141 41497 17175 41531
rect 22109 41497 22143 41531
rect 22293 41497 22327 41531
rect 22477 41497 22511 41531
rect 23121 41497 23155 41531
rect 24501 41497 24535 41531
rect 26801 41497 26835 41531
rect 28457 41497 28491 41531
rect 28733 41497 28767 41531
rect 29193 41497 29227 41531
rect 30021 41497 30055 41531
rect 33885 41497 33919 41531
rect 34437 41497 34471 41531
rect 35081 41497 35115 41531
rect 37565 41497 37599 41531
rect 37749 41497 37783 41531
rect 39405 41497 39439 41531
rect 18613 41429 18647 41463
rect 21833 41429 21867 41463
rect 22569 41429 22603 41463
rect 23489 41429 23523 41463
rect 26617 41429 26651 41463
rect 28273 41429 28307 41463
rect 28641 41429 28675 41463
rect 29377 41429 29411 41463
rect 32781 41429 32815 41463
rect 35173 41429 35207 41463
rect 37473 41429 37507 41463
rect 37933 41429 37967 41463
rect 17509 41225 17543 41259
rect 22477 41225 22511 41259
rect 23489 41225 23523 41259
rect 27997 41225 28031 41259
rect 34345 41225 34379 41259
rect 35173 41225 35207 41259
rect 37657 41225 37691 41259
rect 39221 41225 39255 41259
rect 39589 41225 39623 41259
rect 23857 41157 23891 41191
rect 25973 41157 26007 41191
rect 26433 41157 26467 41191
rect 31861 41157 31895 41191
rect 34713 41157 34747 41191
rect 35633 41157 35667 41191
rect 36829 41157 36863 41191
rect 40049 41157 40083 41191
rect 16129 41089 16163 41123
rect 17877 41089 17911 41123
rect 20269 41089 20303 41123
rect 20545 41089 20579 41123
rect 21096 41089 21130 41123
rect 21189 41089 21223 41123
rect 21281 41089 21315 41123
rect 21465 41089 21499 41123
rect 21557 41089 21591 41123
rect 22845 41089 22879 41123
rect 23673 41089 23707 41123
rect 23949 41089 23983 41123
rect 24133 41089 24167 41123
rect 25789 41089 25823 41123
rect 26065 41089 26099 41123
rect 26157 41089 26191 41123
rect 26249 41089 26283 41123
rect 27813 41089 27847 41123
rect 27997 41089 28031 41123
rect 28273 41089 28307 41123
rect 28549 41089 28583 41123
rect 28733 41089 28767 41123
rect 29101 41089 29135 41123
rect 30113 41089 30147 41123
rect 30941 41089 30975 41123
rect 31585 41089 31619 41123
rect 31769 41089 31803 41123
rect 31953 41089 31987 41123
rect 32321 41089 32355 41123
rect 33149 41089 33183 41123
rect 33333 41089 33367 41123
rect 33517 41089 33551 41123
rect 33609 41089 33643 41123
rect 35541 41089 35575 41123
rect 37013 41089 37047 41123
rect 37105 41089 37139 41123
rect 38117 41089 38151 41123
rect 38301 41089 38335 41123
rect 38761 41089 38795 41123
rect 40233 41089 40267 41123
rect 16037 41021 16071 41055
rect 16865 41021 16899 41055
rect 17969 41021 18003 41055
rect 18061 41021 18095 41055
rect 22937 41021 22971 41055
rect 23121 41021 23155 41055
rect 28365 41021 28399 41055
rect 28457 41021 28491 41055
rect 32413 41021 32447 41055
rect 34805 41021 34839 41055
rect 34897 41021 34931 41055
rect 35725 41021 35759 41055
rect 37749 41021 37783 41055
rect 37841 41021 37875 41055
rect 38209 41021 38243 41055
rect 38853 41021 38887 41055
rect 39037 41021 39071 41055
rect 39681 41021 39715 41055
rect 39773 41021 39807 41055
rect 16497 40953 16531 40987
rect 20361 40953 20395 40987
rect 20453 40953 20487 40987
rect 20821 40953 20855 40987
rect 21281 40953 21315 40987
rect 24041 40953 24075 40987
rect 28089 40953 28123 40987
rect 33425 40953 33459 40987
rect 38393 40953 38427 40987
rect 17417 40885 17451 40919
rect 20729 40885 20763 40919
rect 26065 40885 26099 40919
rect 26433 40885 26467 40919
rect 31033 40885 31067 40919
rect 32597 40885 32631 40919
rect 33793 40885 33827 40919
rect 36829 40885 36863 40919
rect 37289 40885 37323 40919
rect 40417 40885 40451 40919
rect 17141 40681 17175 40715
rect 17785 40681 17819 40715
rect 18613 40681 18647 40715
rect 24961 40681 24995 40715
rect 30113 40681 30147 40715
rect 36264 40681 36298 40715
rect 37749 40681 37783 40715
rect 19441 40613 19475 40647
rect 21189 40613 21223 40647
rect 26065 40613 26099 40647
rect 28733 40613 28767 40647
rect 31033 40613 31067 40647
rect 31125 40613 31159 40647
rect 33057 40613 33091 40647
rect 18337 40545 18371 40579
rect 21097 40545 21131 40579
rect 21465 40545 21499 40579
rect 25329 40545 25363 40579
rect 28457 40545 28491 40579
rect 30665 40545 30699 40579
rect 31493 40545 31527 40579
rect 32873 40545 32907 40579
rect 36001 40545 36035 40579
rect 15393 40477 15427 40511
rect 18797 40477 18831 40511
rect 18889 40477 18923 40511
rect 19257 40477 19291 40511
rect 19441 40477 19475 40511
rect 20545 40477 20579 40511
rect 20729 40477 20763 40511
rect 20821 40477 20855 40511
rect 21005 40477 21039 40511
rect 21281 40477 21315 40511
rect 22783 40477 22817 40511
rect 22937 40477 22971 40511
rect 25145 40477 25179 40511
rect 25237 40477 25271 40511
rect 25421 40477 25455 40511
rect 25605 40477 25639 40511
rect 26433 40477 26467 40511
rect 27445 40477 27479 40511
rect 27629 40477 27663 40511
rect 27996 40477 28030 40511
rect 28089 40477 28123 40511
rect 28365 40477 28399 40511
rect 28825 40477 28859 40511
rect 29009 40477 29043 40511
rect 29101 40477 29135 40511
rect 29193 40477 29227 40511
rect 29285 40477 29319 40511
rect 30481 40477 30515 40511
rect 32781 40477 32815 40511
rect 33271 40477 33305 40511
rect 33425 40477 33459 40511
rect 39221 40477 39255 40511
rect 15669 40409 15703 40443
rect 18613 40409 18647 40443
rect 19533 40409 19567 40443
rect 20269 40409 20303 40443
rect 18153 40341 18187 40375
rect 18245 40341 18279 40375
rect 20637 40341 20671 40375
rect 22569 40341 22603 40375
rect 25973 40341 26007 40375
rect 27537 40341 27571 40375
rect 27721 40341 27755 40375
rect 30573 40341 30607 40375
rect 32413 40341 32447 40375
rect 16681 40137 16715 40171
rect 17049 40137 17083 40171
rect 17141 40137 17175 40171
rect 17509 40137 17543 40171
rect 17877 40137 17911 40171
rect 23305 40137 23339 40171
rect 36461 40137 36495 40171
rect 39313 40137 39347 40171
rect 39773 40137 39807 40171
rect 17969 40069 18003 40103
rect 23397 40069 23431 40103
rect 32413 40069 32447 40103
rect 36921 40069 36955 40103
rect 38301 40069 38335 40103
rect 39681 40069 39715 40103
rect 18521 40001 18555 40035
rect 19625 40001 19659 40035
rect 20729 40001 20763 40035
rect 22017 40001 22051 40035
rect 22937 40001 22971 40035
rect 24225 40001 24259 40035
rect 24593 40001 24627 40035
rect 24777 40001 24811 40035
rect 25053 40001 25087 40035
rect 25145 40001 25179 40035
rect 25329 40001 25363 40035
rect 25513 40001 25547 40035
rect 25973 40001 26007 40035
rect 27997 40001 28031 40035
rect 31033 40001 31067 40035
rect 32137 40001 32171 40035
rect 32229 40001 32263 40035
rect 17325 39933 17359 39967
rect 18061 39933 18095 39967
rect 18613 39933 18647 39967
rect 20821 39933 20855 39967
rect 21925 39933 21959 39967
rect 23029 39933 23063 39967
rect 26065 39933 26099 39967
rect 26801 39933 26835 39967
rect 27905 39933 27939 39967
rect 39129 39933 39163 39967
rect 39865 39933 39899 39967
rect 21097 39865 21131 39899
rect 25237 39865 25271 39899
rect 28365 39865 28399 39899
rect 30849 39865 30883 39899
rect 36553 39865 36587 39899
rect 18889 39797 18923 39831
rect 22385 39797 22419 39831
rect 22937 39797 22971 39831
rect 24777 39797 24811 39831
rect 32413 39797 32447 39831
rect 30021 39593 30055 39627
rect 30849 39593 30883 39627
rect 32137 39593 32171 39627
rect 32873 39593 32907 39627
rect 35633 39593 35667 39627
rect 34529 39525 34563 39559
rect 39405 39525 39439 39559
rect 18797 39457 18831 39491
rect 22937 39457 22971 39491
rect 24869 39457 24903 39491
rect 25605 39457 25639 39491
rect 30665 39457 30699 39491
rect 31493 39457 31527 39491
rect 32505 39457 32539 39491
rect 32689 39457 32723 39491
rect 35265 39457 35299 39491
rect 40417 39457 40451 39491
rect 18705 39389 18739 39423
rect 22661 39389 22695 39423
rect 22753 39389 22787 39423
rect 22845 39389 22879 39423
rect 24041 39389 24075 39423
rect 24777 39389 24811 39423
rect 25237 39389 25271 39423
rect 25330 39389 25364 39423
rect 31769 39389 31803 39423
rect 32413 39389 32447 39423
rect 32597 39389 32631 39423
rect 32873 39389 32907 39423
rect 32965 39389 32999 39423
rect 34253 39389 34287 39423
rect 34345 39389 34379 39423
rect 34897 39389 34931 39423
rect 34989 39389 35023 39423
rect 35633 39389 35667 39423
rect 35817 39389 35851 39423
rect 37289 39389 37323 39423
rect 37473 39389 37507 39423
rect 39681 39389 39715 39423
rect 41245 39389 41279 39423
rect 42165 39389 42199 39423
rect 30389 39321 30423 39355
rect 31309 39321 31343 39355
rect 31953 39321 31987 39355
rect 34529 39321 34563 39355
rect 35357 39321 35391 39355
rect 39405 39321 39439 39355
rect 40233 39321 40267 39355
rect 40693 39321 40727 39355
rect 19073 39253 19107 39287
rect 22477 39253 22511 39287
rect 25145 39253 25179 39287
rect 30481 39253 30515 39287
rect 31217 39253 31251 39287
rect 32229 39253 32263 39287
rect 33241 39253 33275 39287
rect 34713 39253 34747 39287
rect 35449 39253 35483 39287
rect 37381 39253 37415 39287
rect 39589 39253 39623 39287
rect 39865 39253 39899 39287
rect 40325 39253 40359 39287
rect 41521 39253 41555 39287
rect 17141 39049 17175 39083
rect 17509 39049 17543 39083
rect 25053 39049 25087 39083
rect 29101 39049 29135 39083
rect 40969 39049 41003 39083
rect 41429 39049 41463 39083
rect 17049 38981 17083 39015
rect 20237 38981 20271 39015
rect 20453 38981 20487 39015
rect 21281 38981 21315 39015
rect 22109 38981 22143 39015
rect 25605 38981 25639 39015
rect 28641 38981 28675 39015
rect 30205 38981 30239 39015
rect 39497 38981 39531 39015
rect 14749 38913 14783 38947
rect 18521 38913 18555 38947
rect 19625 38913 19659 38947
rect 19718 38913 19752 38947
rect 20821 38913 20855 38947
rect 21465 38913 21499 38947
rect 21649 38913 21683 38947
rect 21833 38913 21867 38947
rect 21925 38913 21959 38947
rect 22201 38913 22235 38947
rect 24777 38913 24811 38947
rect 24961 38913 24995 38947
rect 25053 38913 25087 38947
rect 25145 38913 25179 38947
rect 25237 38913 25271 38947
rect 25421 38913 25455 38947
rect 25789 38913 25823 38947
rect 28089 38913 28123 38947
rect 28365 38913 28399 38947
rect 28549 38913 28583 38947
rect 28917 38913 28951 38947
rect 30113 38913 30147 38947
rect 30297 38913 30331 38947
rect 30757 38913 30791 38947
rect 31309 38913 31343 38947
rect 32137 38913 32171 38947
rect 33977 38913 34011 38947
rect 36185 38913 36219 38947
rect 36461 38913 36495 38947
rect 36645 38913 36679 38947
rect 37657 38913 37691 38947
rect 38117 38913 38151 38947
rect 38209 38913 38243 38947
rect 38393 38913 38427 38947
rect 38791 38913 38825 38947
rect 38945 38913 38979 38947
rect 15025 38845 15059 38879
rect 16865 38845 16899 38879
rect 18153 38845 18187 38879
rect 18429 38845 18463 38879
rect 19993 38845 20027 38879
rect 22477 38845 22511 38879
rect 24593 38845 24627 38879
rect 28733 38845 28767 38879
rect 30849 38845 30883 38879
rect 32413 38845 32447 38879
rect 36093 38845 36127 38879
rect 36553 38845 36587 38879
rect 37749 38845 37783 38879
rect 38577 38845 38611 38879
rect 39221 38845 39255 38879
rect 41521 38845 41555 38879
rect 41613 38845 41647 38879
rect 20637 38777 20671 38811
rect 23949 38777 23983 38811
rect 25421 38777 25455 38811
rect 35725 38777 35759 38811
rect 37289 38777 37323 38811
rect 38301 38777 38335 38811
rect 16497 38709 16531 38743
rect 17601 38709 17635 38743
rect 18889 38709 18923 38743
rect 20085 38709 20119 38743
rect 20269 38709 20303 38743
rect 22109 38709 22143 38743
rect 24041 38709 24075 38743
rect 25973 38709 26007 38743
rect 28227 38709 28261 38743
rect 28457 38709 28491 38743
rect 28641 38709 28675 38743
rect 30481 38709 30515 38743
rect 31125 38709 31159 38743
rect 33885 38709 33919 38743
rect 34240 38709 34274 38743
rect 35909 38709 35943 38743
rect 37933 38709 37967 38743
rect 41061 38709 41095 38743
rect 16681 38505 16715 38539
rect 22477 38505 22511 38539
rect 24869 38505 24903 38539
rect 26065 38505 26099 38539
rect 32137 38505 32171 38539
rect 34161 38505 34195 38539
rect 35265 38505 35299 38539
rect 39865 38505 39899 38539
rect 42165 38505 42199 38539
rect 16589 38437 16623 38471
rect 19717 38437 19751 38471
rect 20269 38437 20303 38471
rect 22017 38437 22051 38471
rect 26985 38437 27019 38471
rect 38209 38437 38243 38471
rect 39405 38437 39439 38471
rect 17325 38369 17359 38403
rect 19625 38369 19659 38403
rect 21005 38369 21039 38403
rect 21557 38369 21591 38403
rect 22661 38369 22695 38403
rect 23121 38369 23155 38403
rect 25329 38369 25363 38403
rect 27353 38369 27387 38403
rect 27537 38369 27571 38403
rect 28181 38369 28215 38403
rect 28641 38369 28675 38403
rect 32321 38369 32355 38403
rect 32689 38369 32723 38403
rect 35357 38369 35391 38403
rect 37105 38369 37139 38403
rect 38301 38369 38335 38403
rect 40417 38369 40451 38403
rect 40693 38369 40727 38403
rect 14841 38301 14875 38335
rect 17509 38301 17543 38335
rect 19533 38301 19567 38335
rect 19809 38301 19843 38335
rect 20545 38301 20579 38335
rect 21649 38301 21683 38335
rect 21741 38301 21775 38335
rect 21833 38301 21867 38335
rect 22017 38301 22051 38335
rect 22293 38301 22327 38335
rect 22753 38301 22787 38335
rect 24409 38301 24443 38335
rect 24593 38301 24627 38335
rect 24777 38301 24811 38335
rect 24961 38301 24995 38335
rect 25237 38301 25271 38335
rect 25881 38301 25915 38335
rect 26709 38301 26743 38335
rect 26985 38301 27019 38335
rect 27261 38301 27295 38335
rect 27445 38301 27479 38335
rect 28089 38301 28123 38335
rect 28733 38301 28767 38335
rect 32413 38301 32447 38335
rect 32781 38301 32815 38335
rect 34805 38301 34839 38335
rect 34897 38301 34931 38335
rect 34989 38301 35023 38335
rect 35081 38301 35115 38335
rect 37749 38301 37783 38335
rect 38117 38301 38151 38335
rect 38393 38301 38427 38335
rect 38577 38301 38611 38335
rect 39405 38301 39439 38335
rect 39497 38301 39531 38335
rect 39681 38301 39715 38335
rect 40049 38301 40083 38335
rect 15117 38233 15151 38267
rect 17049 38233 17083 38267
rect 18429 38233 18463 38267
rect 18797 38233 18831 38267
rect 20269 38233 20303 38267
rect 20453 38233 20487 38267
rect 20637 38233 20671 38267
rect 20821 38233 20855 38267
rect 22201 38233 22235 38267
rect 23029 38233 23063 38267
rect 24501 38233 24535 38267
rect 25697 38233 25731 38267
rect 26801 38233 26835 38267
rect 34345 38233 34379 38267
rect 34529 38233 34563 38267
rect 35633 38233 35667 38267
rect 40233 38233 40267 38267
rect 17141 38165 17175 38199
rect 17693 38165 17727 38199
rect 19349 38165 19383 38199
rect 21373 38165 21407 38199
rect 25605 38165 25639 38199
rect 27077 38165 27111 38199
rect 28457 38165 28491 38199
rect 29101 38165 29135 38199
rect 37197 38165 37231 38199
rect 37933 38165 37967 38199
rect 15669 37961 15703 37995
rect 16037 37961 16071 37995
rect 16681 37961 16715 37995
rect 28273 37961 28307 37995
rect 29561 37961 29595 37995
rect 35633 37961 35667 37995
rect 36001 37961 36035 37995
rect 39957 37961 39991 37995
rect 40325 37961 40359 37995
rect 41153 37961 41187 37995
rect 17417 37893 17451 37927
rect 17785 37893 17819 37927
rect 18429 37893 18463 37927
rect 19073 37893 19107 37927
rect 21557 37893 21591 37927
rect 40693 37893 40727 37927
rect 41613 37893 41647 37927
rect 16129 37825 16163 37859
rect 18337 37825 18371 37859
rect 21189 37825 21223 37859
rect 21281 37825 21315 37859
rect 25421 37825 25455 37859
rect 27169 37825 27203 37859
rect 27261 37825 27295 37859
rect 28089 37825 28123 37859
rect 28549 37825 28583 37859
rect 29469 37825 29503 37859
rect 29929 37825 29963 37859
rect 33793 37825 33827 37859
rect 36093 37825 36127 37859
rect 37841 37825 37875 37859
rect 39957 37825 39991 37859
rect 40141 37825 40175 37859
rect 40785 37825 40819 37859
rect 41521 37825 41555 37859
rect 13369 37757 13403 37791
rect 13645 37757 13679 37791
rect 16313 37757 16347 37791
rect 17233 37757 17267 37791
rect 18521 37757 18555 37791
rect 18797 37757 18831 37791
rect 21649 37757 21683 37791
rect 22477 37757 22511 37791
rect 23029 37757 23063 37791
rect 27537 37757 27571 37791
rect 27629 37757 27663 37791
rect 28273 37757 28307 37791
rect 29653 37757 29687 37791
rect 30481 37757 30515 37791
rect 36185 37757 36219 37791
rect 37933 37757 37967 37791
rect 38117 37757 38151 37791
rect 38577 37757 38611 37791
rect 40877 37757 40911 37791
rect 41705 37757 41739 37791
rect 15117 37689 15151 37723
rect 28457 37689 28491 37723
rect 37473 37689 37507 37723
rect 38301 37689 38335 37723
rect 17969 37621 18003 37655
rect 20545 37621 20579 37655
rect 21005 37621 21039 37655
rect 25329 37621 25363 37655
rect 26985 37621 27019 37655
rect 27813 37621 27847 37655
rect 29101 37621 29135 37655
rect 16221 37417 16255 37451
rect 17049 37417 17083 37451
rect 19257 37417 19291 37451
rect 22385 37417 22419 37451
rect 15669 37281 15703 37315
rect 16497 37281 16531 37315
rect 17601 37281 17635 37315
rect 20637 37281 20671 37315
rect 20913 37281 20947 37315
rect 23029 37281 23063 37315
rect 24869 37281 24903 37315
rect 24961 37281 24995 37315
rect 26249 37281 26283 37315
rect 26525 37281 26559 37315
rect 32045 37281 32079 37315
rect 33701 37281 33735 37315
rect 34161 37281 34195 37315
rect 13277 37213 13311 37247
rect 14841 37213 14875 37247
rect 17325 37213 17359 37247
rect 19809 37213 19843 37247
rect 20269 37213 20303 37247
rect 25789 37213 25823 37247
rect 30849 37213 30883 37247
rect 31033 37213 31067 37247
rect 31309 37213 31343 37247
rect 31493 37213 31527 37247
rect 32137 37213 32171 37247
rect 35081 37213 35115 37247
rect 35265 37213 35299 37247
rect 37381 37213 37415 37247
rect 37565 37213 37599 37247
rect 42165 37213 42199 37247
rect 14105 37145 14139 37179
rect 15761 37145 15795 37179
rect 16681 37145 16715 37179
rect 20361 37145 20395 37179
rect 23121 37145 23155 37179
rect 32873 37145 32907 37179
rect 33977 37145 34011 37179
rect 15853 37077 15887 37111
rect 16589 37077 16623 37111
rect 19073 37077 19107 37111
rect 23213 37077 23247 37111
rect 23581 37077 23615 37111
rect 24409 37077 24443 37111
rect 24777 37077 24811 37111
rect 25237 37077 25271 37111
rect 27997 37077 28031 37111
rect 30941 37077 30975 37111
rect 31401 37077 31435 37111
rect 32505 37077 32539 37111
rect 35265 37077 35299 37111
rect 37473 37077 37507 37111
rect 41521 37077 41555 37111
rect 20361 36873 20395 36907
rect 23213 36873 23247 36907
rect 25053 36873 25087 36907
rect 25973 36873 26007 36907
rect 31309 36873 31343 36907
rect 31953 36873 31987 36907
rect 35357 36873 35391 36907
rect 37289 36873 37323 36907
rect 40233 36873 40267 36907
rect 41061 36873 41095 36907
rect 7297 36805 7331 36839
rect 19165 36805 19199 36839
rect 23581 36805 23615 36839
rect 30573 36805 30607 36839
rect 39589 36805 39623 36839
rect 40049 36805 40083 36839
rect 8125 36737 8159 36771
rect 15945 36737 15979 36771
rect 17509 36737 17543 36771
rect 17693 36737 17727 36771
rect 17785 36737 17819 36771
rect 18705 36737 18739 36771
rect 18797 36737 18831 36771
rect 18981 36737 19015 36771
rect 19441 36737 19475 36771
rect 19533 36737 19567 36771
rect 19809 36737 19843 36771
rect 20269 36737 20303 36771
rect 20729 36737 20763 36771
rect 23305 36737 23339 36771
rect 25881 36737 25915 36771
rect 26985 36737 27019 36771
rect 28549 36737 28583 36771
rect 30481 36737 30515 36771
rect 30665 36737 30699 36771
rect 30849 36737 30883 36771
rect 30941 36737 30975 36771
rect 31125 36737 31159 36771
rect 31585 36737 31619 36771
rect 32137 36737 32171 36771
rect 34897 36737 34931 36771
rect 35541 36737 35575 36771
rect 35817 36737 35851 36771
rect 36369 36737 36403 36771
rect 37473 36737 37507 36771
rect 37657 36737 37691 36771
rect 37749 36737 37783 36771
rect 37933 36737 37967 36771
rect 38025 36737 38059 36771
rect 38118 36737 38152 36771
rect 39497 36737 39531 36771
rect 39681 36737 39715 36771
rect 39773 36737 39807 36771
rect 39865 36737 39899 36771
rect 40141 36737 40175 36771
rect 40325 36737 40359 36771
rect 40417 36737 40451 36771
rect 3801 36669 3835 36703
rect 4077 36669 4111 36703
rect 15577 36669 15611 36703
rect 16221 36669 16255 36703
rect 17233 36669 17267 36703
rect 20821 36669 20855 36703
rect 21005 36669 21039 36703
rect 22661 36669 22695 36703
rect 26157 36669 26191 36703
rect 27537 36669 27571 36703
rect 28825 36669 28859 36703
rect 31493 36669 31527 36703
rect 32413 36669 32447 36703
rect 33885 36669 33919 36703
rect 34529 36669 34563 36703
rect 34805 36669 34839 36703
rect 35633 36669 35667 36703
rect 36461 36669 36495 36703
rect 41153 36669 41187 36703
rect 41245 36669 41279 36703
rect 42073 36669 42107 36703
rect 16129 36601 16163 36635
rect 31033 36601 31067 36635
rect 35265 36601 35299 36635
rect 35725 36601 35759 36635
rect 36001 36601 36035 36635
rect 37565 36601 37599 36635
rect 5549 36533 5583 36567
rect 15025 36533 15059 36567
rect 15761 36533 15795 36567
rect 16681 36533 16715 36567
rect 17969 36533 18003 36567
rect 19257 36533 19291 36567
rect 19717 36533 19751 36567
rect 20177 36533 20211 36567
rect 25513 36533 25547 36567
rect 30297 36533 30331 36567
rect 33977 36533 34011 36567
rect 38209 36533 38243 36567
rect 40049 36533 40083 36567
rect 40693 36533 40727 36567
rect 41521 36533 41555 36567
rect 3893 36329 3927 36363
rect 13829 36329 13863 36363
rect 16773 36329 16807 36363
rect 19901 36329 19935 36363
rect 20545 36329 20579 36363
rect 30757 36329 30791 36363
rect 30941 36329 30975 36363
rect 31493 36329 31527 36363
rect 32229 36329 32263 36363
rect 34437 36329 34471 36363
rect 35173 36329 35207 36363
rect 36645 36329 36679 36363
rect 37197 36329 37231 36363
rect 39037 36329 39071 36363
rect 39957 36329 39991 36363
rect 42165 36329 42199 36363
rect 4537 36261 4571 36295
rect 29009 36261 29043 36295
rect 34345 36261 34379 36295
rect 37565 36261 37599 36295
rect 39681 36261 39715 36295
rect 10701 36193 10735 36227
rect 12081 36193 12115 36227
rect 17601 36193 17635 36227
rect 21189 36193 21223 36227
rect 21925 36193 21959 36227
rect 23397 36193 23431 36227
rect 30665 36193 30699 36227
rect 32689 36193 32723 36227
rect 32873 36193 32907 36227
rect 34785 36193 34819 36227
rect 35357 36193 35391 36227
rect 37013 36193 37047 36227
rect 40693 36193 40727 36227
rect 4077 36125 4111 36159
rect 4445 36125 4479 36159
rect 4813 36125 4847 36159
rect 4905 36125 4939 36159
rect 5089 36125 5123 36159
rect 5825 36125 5859 36159
rect 6009 36125 6043 36159
rect 6193 36125 6227 36159
rect 6561 36125 6595 36159
rect 6837 36125 6871 36159
rect 8677 36125 8711 36159
rect 14105 36125 14139 36159
rect 15025 36125 15059 36159
rect 16865 36125 16899 36159
rect 16958 36125 16992 36159
rect 17325 36125 17359 36159
rect 19257 36125 19291 36159
rect 23673 36125 23707 36159
rect 25053 36125 25087 36159
rect 27261 36125 27295 36159
rect 29193 36125 29227 36159
rect 29377 36125 29411 36159
rect 30113 36125 30147 36159
rect 30297 36125 30331 36159
rect 31217 36125 31251 36159
rect 31309 36125 31343 36159
rect 32597 36125 32631 36159
rect 33057 36125 33091 36159
rect 33241 36125 33275 36159
rect 33517 36125 33551 36159
rect 34989 36125 35023 36159
rect 35081 36125 35115 36159
rect 36921 36125 36955 36159
rect 37381 36125 37415 36159
rect 37473 36125 37507 36159
rect 37657 36125 37691 36159
rect 37841 36125 37875 36159
rect 38117 36125 38151 36159
rect 38669 36125 38703 36159
rect 39037 36125 39071 36159
rect 39313 36125 39347 36159
rect 40417 36125 40451 36159
rect 4169 36057 4203 36091
rect 4261 36057 4295 36091
rect 4537 36057 4571 36091
rect 6377 36057 6411 36091
rect 8401 36057 8435 36091
rect 10425 36057 10459 36091
rect 12357 36057 12391 36091
rect 15301 36057 15335 36091
rect 25329 36057 25363 36091
rect 27537 36057 27571 36091
rect 29285 36057 29319 36091
rect 30481 36057 30515 36091
rect 31125 36057 31159 36091
rect 31493 36057 31527 36091
rect 33333 36057 33367 36091
rect 33977 36057 34011 36091
rect 34713 36057 34747 36091
rect 38393 36057 38427 36091
rect 38577 36057 38611 36091
rect 39129 36057 39163 36091
rect 39497 36057 39531 36091
rect 40141 36057 40175 36091
rect 40325 36057 40359 36091
rect 4721 35989 4755 36023
rect 4997 35989 5031 36023
rect 6745 35989 6779 36023
rect 6929 35989 6963 36023
rect 8953 35989 8987 36023
rect 14749 35989 14783 36023
rect 17233 35989 17267 36023
rect 19073 35989 19107 36023
rect 20913 35989 20947 36023
rect 21005 35989 21039 36023
rect 26801 35989 26835 36023
rect 29561 35989 29595 36023
rect 30915 35989 30949 36023
rect 33149 35989 33183 36023
rect 33701 35989 33735 36023
rect 34897 35989 34931 36023
rect 35357 35989 35391 36023
rect 37939 35989 37973 36023
rect 38025 35989 38059 36023
rect 38209 35989 38243 36023
rect 38853 35989 38887 36023
rect 8401 35785 8435 35819
rect 9965 35785 9999 35819
rect 13323 35785 13357 35819
rect 16221 35785 16255 35819
rect 17233 35785 17267 35819
rect 18797 35785 18831 35819
rect 22845 35785 22879 35819
rect 22937 35785 22971 35819
rect 23397 35785 23431 35819
rect 27997 35785 28031 35819
rect 28457 35785 28491 35819
rect 31677 35785 31711 35819
rect 34621 35785 34655 35819
rect 39313 35785 39347 35819
rect 41337 35785 41371 35819
rect 5549 35717 5583 35751
rect 5641 35717 5675 35751
rect 6377 35717 6411 35751
rect 8769 35717 8803 35751
rect 8907 35717 8941 35751
rect 9873 35717 9907 35751
rect 10241 35717 10275 35751
rect 14013 35717 14047 35751
rect 14749 35717 14783 35751
rect 18521 35717 18555 35751
rect 20913 35717 20947 35751
rect 22477 35717 22511 35751
rect 28365 35717 28399 35751
rect 30205 35717 30239 35751
rect 30849 35717 30883 35751
rect 31769 35717 31803 35751
rect 34529 35717 34563 35751
rect 34713 35717 34747 35751
rect 35541 35717 35575 35751
rect 2697 35649 2731 35683
rect 4721 35649 4755 35683
rect 4905 35649 4939 35683
rect 4997 35649 5031 35683
rect 5365 35649 5399 35683
rect 5733 35649 5767 35683
rect 7297 35649 7331 35683
rect 8585 35649 8619 35683
rect 8677 35649 8711 35683
rect 9045 35649 9079 35683
rect 10149 35649 10183 35683
rect 10333 35649 10367 35683
rect 10517 35649 10551 35683
rect 10609 35649 10643 35683
rect 10793 35649 10827 35683
rect 10885 35649 10919 35683
rect 10977 35649 11011 35683
rect 11161 35649 11195 35683
rect 11529 35649 11563 35683
rect 13645 35649 13679 35683
rect 13829 35649 13863 35683
rect 13921 35649 13955 35683
rect 14197 35649 14231 35683
rect 14473 35649 14507 35683
rect 17325 35649 17359 35683
rect 17785 35649 17819 35683
rect 21557 35649 21591 35683
rect 23305 35649 23339 35683
rect 24409 35649 24443 35683
rect 33241 35649 33275 35683
rect 33701 35649 33735 35683
rect 34437 35649 34471 35683
rect 35081 35649 35115 35683
rect 35173 35649 35207 35683
rect 35449 35649 35483 35683
rect 35725 35649 35759 35683
rect 35909 35649 35943 35683
rect 36277 35649 36311 35683
rect 38025 35649 38059 35683
rect 38577 35649 38611 35683
rect 39129 35649 39163 35683
rect 39313 35649 39347 35683
rect 39497 35649 39531 35683
rect 39589 35649 39623 35683
rect 2973 35581 3007 35615
rect 4813 35581 4847 35615
rect 6929 35581 6963 35615
rect 9321 35581 9355 35615
rect 11897 35581 11931 35615
rect 14381 35581 14415 35615
rect 17049 35581 17083 35615
rect 19349 35581 19383 35615
rect 19901 35581 19935 35615
rect 20453 35581 20487 35615
rect 21005 35581 21039 35615
rect 21189 35581 21223 35615
rect 22293 35581 22327 35615
rect 22385 35581 22419 35615
rect 23581 35581 23615 35615
rect 24685 35581 24719 35615
rect 26157 35581 26191 35615
rect 27537 35581 27571 35615
rect 28641 35581 28675 35615
rect 30297 35581 30331 35615
rect 30481 35581 30515 35615
rect 31401 35581 31435 35615
rect 33333 35581 33367 35615
rect 33517 35581 33551 35615
rect 34345 35581 34379 35615
rect 36001 35581 36035 35615
rect 36185 35581 36219 35615
rect 38117 35581 38151 35615
rect 38301 35581 38335 35615
rect 39865 35581 39899 35615
rect 41521 35581 41555 35615
rect 4537 35513 4571 35547
rect 11069 35513 11103 35547
rect 36093 35513 36127 35547
rect 4445 35445 4479 35479
rect 5917 35445 5951 35479
rect 10609 35445 10643 35479
rect 13461 35445 13495 35479
rect 17693 35445 17727 35479
rect 20545 35445 20579 35479
rect 21465 35445 21499 35479
rect 26985 35445 27019 35479
rect 29837 35445 29871 35479
rect 32873 35445 32907 35479
rect 34897 35445 34931 35479
rect 35357 35445 35391 35479
rect 37657 35445 37691 35479
rect 42165 35445 42199 35479
rect 3157 35241 3191 35275
rect 3985 35241 4019 35275
rect 4721 35241 4755 35275
rect 7113 35241 7147 35275
rect 8217 35241 8251 35275
rect 8677 35241 8711 35275
rect 12265 35241 12299 35275
rect 13737 35241 13771 35275
rect 15209 35241 15243 35275
rect 18521 35241 18555 35275
rect 24869 35241 24903 35275
rect 28641 35241 28675 35275
rect 31309 35241 31343 35275
rect 33885 35241 33919 35275
rect 36369 35241 36403 35275
rect 40141 35241 40175 35275
rect 41981 35241 42015 35275
rect 8033 35173 8067 35207
rect 5549 35105 5583 35139
rect 14105 35105 14139 35139
rect 15669 35105 15703 35139
rect 15853 35105 15887 35139
rect 17141 35105 17175 35139
rect 19993 35105 20027 35139
rect 22017 35105 22051 35139
rect 23397 35105 23431 35139
rect 25421 35105 25455 35139
rect 29285 35105 29319 35139
rect 29837 35105 29871 35139
rect 31953 35105 31987 35139
rect 32137 35105 32171 35139
rect 32413 35105 32447 35139
rect 36001 35105 36035 35139
rect 36093 35105 36127 35139
rect 39129 35105 39163 35139
rect 40693 35105 40727 35139
rect 3341 35037 3375 35071
rect 3525 35037 3559 35071
rect 3617 35037 3651 35071
rect 4169 35037 4203 35071
rect 4445 35037 4479 35071
rect 5273 35037 5307 35071
rect 7297 35037 7331 35071
rect 8493 35037 8527 35071
rect 8677 35037 8711 35071
rect 12449 35037 12483 35071
rect 12725 35037 12759 35071
rect 12909 35037 12943 35071
rect 13001 35037 13035 35071
rect 16037 35037 16071 35071
rect 17408 35037 17442 35071
rect 18705 35037 18739 35071
rect 19809 35037 19843 35071
rect 25237 35037 25271 35071
rect 26249 35037 26283 35071
rect 26893 35037 26927 35071
rect 29561 35037 29595 35071
rect 35265 35037 35299 35071
rect 37013 35037 37047 35071
rect 38301 35037 38335 35071
rect 40509 35037 40543 35071
rect 41521 35037 41555 35071
rect 41797 35037 41831 35071
rect 4705 34969 4739 35003
rect 4905 34969 4939 35003
rect 7481 34969 7515 35003
rect 8401 34969 8435 35003
rect 13185 34969 13219 35003
rect 13369 34969 13403 35003
rect 13829 34969 13863 35003
rect 20260 34969 20294 35003
rect 21833 34969 21867 35003
rect 23305 34969 23339 35003
rect 25697 34969 25731 35003
rect 27169 34969 27203 35003
rect 38945 34969 38979 35003
rect 4353 34901 4387 34935
rect 4537 34901 4571 34935
rect 7021 34901 7055 34935
rect 8191 34901 8225 34935
rect 14749 34901 14783 34935
rect 15577 34901 15611 34935
rect 16681 34901 16715 34935
rect 19257 34901 19291 34935
rect 21373 34901 21407 34935
rect 21465 34901 21499 34935
rect 21925 34901 21959 34935
rect 22845 34901 22879 34935
rect 23213 34901 23247 34935
rect 25329 34901 25363 34935
rect 28733 34901 28767 34935
rect 31401 34901 31435 34935
rect 34713 34901 34747 34935
rect 35541 34901 35575 34935
rect 35909 34901 35943 34935
rect 38577 34901 38611 34935
rect 39037 34901 39071 34935
rect 40601 34901 40635 34935
rect 40969 34901 41003 34935
rect 3985 34697 4019 34731
rect 11345 34697 11379 34731
rect 15117 34697 15151 34731
rect 17233 34697 17267 34731
rect 18705 34697 18739 34731
rect 19165 34697 19199 34731
rect 21281 34697 21315 34731
rect 22293 34697 22327 34731
rect 24869 34697 24903 34731
rect 25697 34697 25731 34731
rect 27537 34697 27571 34731
rect 27905 34697 27939 34731
rect 31493 34697 31527 34731
rect 31677 34697 31711 34731
rect 40141 34697 40175 34731
rect 40877 34697 40911 34731
rect 41245 34697 41279 34731
rect 41337 34697 41371 34731
rect 16681 34629 16715 34663
rect 18368 34629 18402 34663
rect 20168 34629 20202 34663
rect 23406 34629 23440 34663
rect 25237 34629 25271 34663
rect 26157 34629 26191 34663
rect 29101 34629 29135 34663
rect 33885 34629 33919 34663
rect 34345 34629 34379 34663
rect 35081 34629 35115 34663
rect 37013 34629 37047 34663
rect 37565 34629 37599 34663
rect 39865 34629 39899 34663
rect 41705 34629 41739 34663
rect 3893 34561 3927 34595
rect 4077 34561 4111 34595
rect 5181 34561 5215 34595
rect 5365 34561 5399 34595
rect 5457 34561 5491 34595
rect 8125 34561 8159 34595
rect 8493 34561 8527 34595
rect 8769 34561 8803 34595
rect 9137 34561 9171 34595
rect 9321 34561 9355 34595
rect 16241 34561 16275 34595
rect 17049 34561 17083 34595
rect 18613 34561 18647 34595
rect 19073 34561 19107 34595
rect 19901 34561 19935 34595
rect 24133 34561 24167 34595
rect 26065 34561 26099 34595
rect 31861 34561 31895 34595
rect 32137 34561 32171 34595
rect 39129 34561 39163 34595
rect 40693 34561 40727 34595
rect 41889 34561 41923 34595
rect 8953 34493 8987 34527
rect 9597 34493 9631 34527
rect 12081 34493 12115 34527
rect 12909 34493 12943 34527
rect 14657 34493 14691 34527
rect 16497 34493 16531 34527
rect 19257 34493 19291 34527
rect 23673 34493 23707 34527
rect 24225 34493 24259 34527
rect 24409 34493 24443 34527
rect 25329 34493 25363 34527
rect 25513 34493 25547 34527
rect 26249 34493 26283 34527
rect 27997 34493 28031 34527
rect 28181 34493 28215 34527
rect 28825 34493 28859 34527
rect 29745 34493 29779 34527
rect 30021 34493 30055 34527
rect 34437 34493 34471 34527
rect 34529 34493 34563 34527
rect 34805 34493 34839 34527
rect 37289 34493 37323 34527
rect 39037 34493 39071 34527
rect 41521 34493 41555 34527
rect 8585 34425 8619 34459
rect 8677 34425 8711 34459
rect 36553 34425 36587 34459
rect 5181 34357 5215 34391
rect 5641 34357 5675 34391
rect 8309 34357 8343 34391
rect 9854 34357 9888 34391
rect 11529 34357 11563 34391
rect 13172 34357 13206 34391
rect 23765 34357 23799 34391
rect 33977 34357 34011 34391
rect 36737 34357 36771 34391
rect 6101 34153 6135 34187
rect 8493 34153 8527 34187
rect 9689 34153 9723 34187
rect 11529 34153 11563 34187
rect 13737 34153 13771 34187
rect 14105 34153 14139 34187
rect 16405 34153 16439 34187
rect 21005 34153 21039 34187
rect 25881 34153 25915 34187
rect 27905 34153 27939 34187
rect 30205 34153 30239 34187
rect 33793 34153 33827 34187
rect 39037 34153 39071 34187
rect 40969 34153 41003 34187
rect 11345 34085 11379 34119
rect 15761 34085 15795 34119
rect 6745 34017 6779 34051
rect 9505 34017 9539 34051
rect 11161 34017 11195 34051
rect 11989 34017 12023 34051
rect 14657 34017 14691 34051
rect 16865 34017 16899 34051
rect 17049 34017 17083 34051
rect 19257 34017 19291 34051
rect 21649 34017 21683 34051
rect 26433 34017 26467 34051
rect 28457 34017 28491 34051
rect 30849 34017 30883 34051
rect 32045 34017 32079 34051
rect 32321 34017 32355 34051
rect 34989 34017 35023 34051
rect 37289 34017 37323 34051
rect 40693 34017 40727 34051
rect 41613 34017 41647 34051
rect 5917 33949 5951 33983
rect 6193 33949 6227 33983
rect 9873 33949 9907 33983
rect 9965 33949 9999 33983
rect 10241 33949 10275 33983
rect 10333 33949 10367 33983
rect 10517 33949 10551 33983
rect 14473 33949 14507 33983
rect 15485 33949 15519 33983
rect 15669 33949 15703 33983
rect 15853 33949 15887 33983
rect 22109 33949 22143 33983
rect 23581 33949 23615 33983
rect 24409 33949 24443 33983
rect 31033 33949 31067 33983
rect 40601 33949 40635 33983
rect 41337 33949 41371 33983
rect 7021 33881 7055 33915
rect 10057 33881 10091 33915
rect 10425 33881 10459 33915
rect 11713 33881 11747 33915
rect 12265 33881 12299 33915
rect 19533 33881 19567 33915
rect 23336 33881 23370 33915
rect 24676 33881 24710 33915
rect 26709 33881 26743 33915
rect 27445 33881 27479 33915
rect 28273 33881 28307 33915
rect 30573 33881 30607 33915
rect 35265 33881 35299 33915
rect 37565 33881 37599 33915
rect 5733 33813 5767 33847
rect 8953 33813 8987 33847
rect 10609 33813 10643 33847
rect 11503 33813 11537 33847
rect 14565 33813 14599 33847
rect 14933 33813 14967 33847
rect 16773 33813 16807 33847
rect 21097 33813 21131 33847
rect 21925 33813 21959 33847
rect 22201 33813 22235 33847
rect 25789 33813 25823 33847
rect 26249 33813 26283 33847
rect 26341 33813 26375 33847
rect 28365 33813 28399 33847
rect 30665 33813 30699 33847
rect 36737 33813 36771 33847
rect 40141 33813 40175 33847
rect 40509 33813 40543 33847
rect 41429 33813 41463 33847
rect 11253 33609 11287 33643
rect 12909 33609 12943 33643
rect 16681 33609 16715 33643
rect 19809 33609 19843 33643
rect 20269 33609 20303 33643
rect 21833 33609 21867 33643
rect 23857 33609 23891 33643
rect 23949 33609 23983 33643
rect 24777 33609 24811 33643
rect 26985 33609 27019 33643
rect 27905 33609 27939 33643
rect 30297 33609 30331 33643
rect 30757 33609 30791 33643
rect 31125 33609 31159 33643
rect 31493 33609 31527 33643
rect 31585 33609 31619 33643
rect 33517 33609 33551 33643
rect 33885 33609 33919 33643
rect 34345 33609 34379 33643
rect 36369 33609 36403 33643
rect 37933 33609 37967 33643
rect 38761 33609 38795 33643
rect 41337 33609 41371 33643
rect 41889 33609 41923 33643
rect 2329 33541 2363 33575
rect 2789 33541 2823 33575
rect 5825 33541 5859 33575
rect 7665 33541 7699 33575
rect 8401 33541 8435 33575
rect 12173 33541 12207 33575
rect 27445 33541 27479 33575
rect 30665 33541 30699 33575
rect 32229 33541 32263 33575
rect 39221 33541 39255 33575
rect 2053 33473 2087 33507
rect 2145 33473 2179 33507
rect 2605 33473 2639 33507
rect 2881 33473 2915 33507
rect 4905 33473 4939 33507
rect 5365 33473 5399 33507
rect 5457 33473 5491 33507
rect 5641 33473 5675 33507
rect 8953 33473 8987 33507
rect 9229 33473 9263 33507
rect 11069 33473 11103 33507
rect 11345 33473 11379 33507
rect 11713 33473 11747 33507
rect 15945 33473 15979 33507
rect 17794 33473 17828 33507
rect 18061 33473 18095 33507
rect 18475 33473 18509 33507
rect 18613 33473 18647 33507
rect 18705 33473 18739 33507
rect 18833 33473 18867 33507
rect 18981 33473 19015 33507
rect 20177 33473 20211 33507
rect 22385 33473 22419 33507
rect 23213 33473 23247 33507
rect 24501 33473 24535 33507
rect 25145 33473 25179 33507
rect 26709 33473 26743 33507
rect 27353 33473 27387 33507
rect 28273 33473 28307 33507
rect 28365 33473 28399 33507
rect 33057 33473 33091 33507
rect 33977 33473 34011 33507
rect 34713 33473 34747 33507
rect 38301 33473 38335 33507
rect 38393 33473 38427 33507
rect 39129 33473 39163 33507
rect 39957 33473 39991 33507
rect 40224 33473 40258 33507
rect 41797 33473 41831 33507
rect 4629 33405 4663 33439
rect 5181 33405 5215 33439
rect 5273 33405 5307 33439
rect 8677 33405 8711 33439
rect 8861 33405 8895 33439
rect 9505 33405 9539 33439
rect 11805 33405 11839 33439
rect 12357 33405 12391 33439
rect 13093 33405 13127 33439
rect 20453 33405 20487 33439
rect 25237 33405 25271 33439
rect 25329 33405 25363 33439
rect 27537 33405 27571 33439
rect 28457 33405 28491 33439
rect 30849 33405 30883 33439
rect 31677 33405 31711 33439
rect 32505 33405 32539 33439
rect 34069 33405 34103 33439
rect 34805 33405 34839 33439
rect 34989 33405 35023 33439
rect 36921 33405 36955 33439
rect 38577 33405 38611 33439
rect 39313 33405 39347 33439
rect 41981 33405 42015 33439
rect 11069 33337 11103 33371
rect 16497 33337 16531 33371
rect 41429 33337 41463 33371
rect 2329 33269 2363 33303
rect 2421 33269 2455 33303
rect 3157 33269 3191 33303
rect 4997 33269 5031 33303
rect 6009 33269 6043 33303
rect 8769 33269 8803 33303
rect 10977 33269 11011 33303
rect 11529 33269 11563 33303
rect 13645 33269 13679 33303
rect 18337 33269 18371 33303
rect 26157 33269 26191 33303
rect 33333 33269 33367 33303
rect 4721 33065 4755 33099
rect 4997 33065 5031 33099
rect 5549 33065 5583 33099
rect 7573 33065 7607 33099
rect 9505 33065 9539 33099
rect 12357 33065 12391 33099
rect 12449 33065 12483 33099
rect 17233 33065 17267 33099
rect 18429 33065 18463 33099
rect 21097 33065 21131 33099
rect 22937 33065 22971 33099
rect 24593 33065 24627 33099
rect 26709 33065 26743 33099
rect 38485 33065 38519 33099
rect 41705 33065 41739 33099
rect 3433 32997 3467 33031
rect 5733 32997 5767 33031
rect 10793 32997 10827 33031
rect 14657 32997 14691 33031
rect 15301 32997 15335 33031
rect 28549 32997 28583 33031
rect 32505 32997 32539 33031
rect 3157 32929 3191 32963
rect 3617 32929 3651 32963
rect 7481 32929 7515 32963
rect 10977 32929 11011 32963
rect 14197 32929 14231 32963
rect 14841 32929 14875 32963
rect 15485 32929 15519 32963
rect 16681 32929 16715 32963
rect 16773 32929 16807 32963
rect 19349 32929 19383 32963
rect 21189 32929 21223 32963
rect 29193 32929 29227 32963
rect 31125 32929 31159 32963
rect 33241 32929 33275 32963
rect 34253 32929 34287 32963
rect 35541 32929 35575 32963
rect 39129 32929 39163 32963
rect 3341 32861 3375 32895
rect 4445 32861 4479 32895
rect 4537 32861 4571 32895
rect 5178 32861 5212 32895
rect 5641 32861 5675 32895
rect 7757 32861 7791 32895
rect 7849 32861 7883 32895
rect 9689 32861 9723 32895
rect 9781 32861 9815 32895
rect 9873 32861 9907 32895
rect 9991 32861 10025 32895
rect 10149 32861 10183 32895
rect 10425 32861 10459 32895
rect 10701 32861 10735 32895
rect 10885 32861 10919 32895
rect 11244 32861 11278 32895
rect 13829 32861 13863 32895
rect 14289 32861 14323 32895
rect 14933 32861 14967 32895
rect 17785 32861 17819 32895
rect 19073 32861 19107 32895
rect 23029 32861 23063 32895
rect 25145 32861 25179 32895
rect 25329 32861 25363 32895
rect 27169 32861 27203 32895
rect 30665 32861 30699 32895
rect 36369 32861 36403 32895
rect 37105 32861 37139 32895
rect 40325 32861 40359 32895
rect 40592 32861 40626 32895
rect 2881 32793 2915 32827
rect 3617 32793 3651 32827
rect 4077 32793 4111 32827
rect 4169 32793 4203 32827
rect 7205 32793 7239 32827
rect 8125 32793 8159 32827
rect 8217 32793 8251 32827
rect 10609 32793 10643 32827
rect 13584 32793 13618 32827
rect 19625 32793 19659 32827
rect 21465 32793 21499 32827
rect 25596 32793 25630 32827
rect 27436 32793 27470 32827
rect 28641 32793 28675 32827
rect 31392 32793 31426 32827
rect 34069 32793 34103 32827
rect 35357 32793 35391 32827
rect 37372 32793 37406 32827
rect 1409 32725 1443 32759
rect 5181 32725 5215 32759
rect 10241 32725 10275 32759
rect 16037 32725 16071 32759
rect 16865 32725 16899 32759
rect 23213 32725 23247 32759
rect 30113 32725 30147 32759
rect 32597 32725 32631 32759
rect 33701 32725 33735 32759
rect 34161 32725 34195 32759
rect 34989 32725 35023 32759
rect 35449 32725 35483 32759
rect 35817 32725 35851 32759
rect 38577 32725 38611 32759
rect 2789 32521 2823 32555
rect 3249 32521 3283 32555
rect 4429 32521 4463 32555
rect 6009 32521 6043 32555
rect 8033 32521 8067 32555
rect 34161 32521 34195 32555
rect 36001 32521 36035 32555
rect 38669 32521 38703 32555
rect 41061 32521 41095 32555
rect 2421 32453 2455 32487
rect 4629 32453 4663 32487
rect 5641 32453 5675 32487
rect 12081 32453 12115 32487
rect 13737 32453 13771 32487
rect 16865 32453 16899 32487
rect 18153 32453 18187 32487
rect 20637 32453 20671 32487
rect 21189 32453 21223 32487
rect 21373 32453 21407 32487
rect 22201 32453 22235 32487
rect 24409 32453 24443 32487
rect 26249 32453 26283 32487
rect 30389 32453 30423 32487
rect 2237 32385 2271 32419
rect 2513 32385 2547 32419
rect 2605 32385 2639 32419
rect 3157 32385 3191 32419
rect 3525 32385 3559 32419
rect 4905 32385 4939 32419
rect 4997 32385 5031 32419
rect 5457 32385 5491 32419
rect 5733 32385 5767 32419
rect 5825 32385 5859 32419
rect 6377 32385 6411 32419
rect 7941 32385 7975 32419
rect 10149 32385 10183 32419
rect 13921 32385 13955 32419
rect 15862 32385 15896 32419
rect 16129 32385 16163 32419
rect 17693 32385 17727 32419
rect 17877 32385 17911 32419
rect 20545 32385 20579 32419
rect 20729 32385 20763 32419
rect 20913 32385 20947 32419
rect 21005 32385 21039 32419
rect 22063 32385 22097 32419
rect 22293 32385 22327 32419
rect 22477 32385 22511 32419
rect 24317 32385 24351 32419
rect 24593 32385 24627 32419
rect 25605 32385 25639 32419
rect 26157 32385 26191 32419
rect 27997 32385 28031 32419
rect 28089 32385 28123 32419
rect 28457 32385 28491 32419
rect 28724 32385 28758 32419
rect 30297 32385 30331 32419
rect 31585 32385 31619 32419
rect 33048 32385 33082 32419
rect 34529 32385 34563 32419
rect 34796 32385 34830 32419
rect 37545 32385 37579 32419
rect 39313 32385 39347 32419
rect 39681 32385 39715 32419
rect 39948 32385 39982 32419
rect 41705 32385 41739 32419
rect 41889 32385 41923 32419
rect 3709 32317 3743 32351
rect 5089 32317 5123 32351
rect 5181 32317 5215 32351
rect 14473 32317 14507 32351
rect 19625 32317 19659 32351
rect 24041 32317 24075 32351
rect 24777 32317 24811 32351
rect 26341 32317 26375 32351
rect 28273 32317 28307 32351
rect 30481 32317 30515 32351
rect 32781 32317 32815 32351
rect 36553 32317 36587 32351
rect 37289 32317 37323 32351
rect 6561 32249 6595 32283
rect 20361 32249 20395 32283
rect 25789 32249 25823 32283
rect 27629 32249 27663 32283
rect 29929 32249 29963 32283
rect 4261 32181 4295 32215
rect 4445 32181 4479 32215
rect 4721 32181 4755 32215
rect 10057 32181 10091 32215
rect 14749 32181 14783 32215
rect 21925 32181 21959 32215
rect 22569 32181 22603 32215
rect 25053 32181 25087 32215
rect 29837 32181 29871 32215
rect 31033 32181 31067 32215
rect 35909 32181 35943 32215
rect 38761 32181 38795 32215
rect 41153 32181 41187 32215
rect 42073 32181 42107 32215
rect 4629 31977 4663 32011
rect 5457 31977 5491 32011
rect 5641 31977 5675 32011
rect 13829 31977 13863 32011
rect 15485 31977 15519 32011
rect 15577 31977 15611 32011
rect 18153 31977 18187 32011
rect 19993 31977 20027 32011
rect 22293 31977 22327 32011
rect 24041 31977 24075 32011
rect 25789 31977 25823 32011
rect 27261 31977 27295 32011
rect 31125 31977 31159 32011
rect 34437 31977 34471 32011
rect 37289 31977 37323 32011
rect 38117 31977 38151 32011
rect 39865 31977 39899 32011
rect 28733 31909 28767 31943
rect 31217 31909 31251 31943
rect 9137 31841 9171 31875
rect 13185 31841 13219 31875
rect 13369 31841 13403 31875
rect 16221 31841 16255 31875
rect 16405 31841 16439 31875
rect 19441 31841 19475 31875
rect 35081 31841 35115 31875
rect 37749 31841 37783 31875
rect 37841 31841 37875 31875
rect 38577 31841 38611 31875
rect 38669 31841 38703 31875
rect 39129 31841 39163 31875
rect 40325 31841 40359 31875
rect 40417 31841 40451 31875
rect 41521 31841 41555 31875
rect 3249 31773 3283 31807
rect 4813 31773 4847 31807
rect 4997 31773 5031 31807
rect 6745 31773 6779 31807
rect 11529 31773 11563 31807
rect 12081 31773 12115 31807
rect 14105 31773 14139 31807
rect 16037 31773 16071 31807
rect 21925 31773 21959 31807
rect 23489 31773 23523 31807
rect 23673 31773 23707 31807
rect 23773 31773 23807 31807
rect 23881 31773 23915 31807
rect 24409 31773 24443 31807
rect 25881 31773 25915 31807
rect 27353 31773 27387 31807
rect 29745 31773 29779 31807
rect 30012 31773 30046 31807
rect 32597 31773 32631 31807
rect 33057 31773 33091 31807
rect 33324 31773 33358 31807
rect 39681 31773 39715 31807
rect 40785 31773 40819 31807
rect 41429 31773 41463 31807
rect 42165 31773 42199 31807
rect 5273 31705 5307 31739
rect 7021 31705 7055 31739
rect 9413 31705 9447 31739
rect 14372 31705 14406 31739
rect 16681 31705 16715 31739
rect 19625 31705 19659 31739
rect 22109 31705 22143 31739
rect 24676 31705 24710 31739
rect 26148 31705 26182 31739
rect 27620 31705 27654 31739
rect 28917 31705 28951 31739
rect 29285 31705 29319 31739
rect 32330 31705 32364 31739
rect 35357 31705 35391 31739
rect 3341 31637 3375 31671
rect 5473 31637 5507 31671
rect 8493 31637 8527 31671
rect 10885 31637 10919 31671
rect 10977 31637 11011 31671
rect 13461 31637 13495 31671
rect 15945 31637 15979 31671
rect 19533 31637 19567 31671
rect 36829 31637 36863 31671
rect 37657 31637 37691 31671
rect 38485 31637 38519 31671
rect 40233 31637 40267 31671
rect 7389 31433 7423 31467
rect 9321 31433 9355 31467
rect 14473 31433 14507 31467
rect 16957 31433 16991 31467
rect 17785 31433 17819 31467
rect 22109 31433 22143 31467
rect 23949 31433 23983 31467
rect 24869 31433 24903 31467
rect 25329 31433 25363 31467
rect 26065 31433 26099 31467
rect 30389 31433 30423 31467
rect 30849 31433 30883 31467
rect 31217 31433 31251 31467
rect 32137 31433 32171 31467
rect 32597 31433 32631 31467
rect 33333 31433 33367 31467
rect 33701 31433 33735 31467
rect 41061 31433 41095 31467
rect 7757 31365 7791 31399
rect 7895 31365 7929 31399
rect 8493 31365 8527 31399
rect 9045 31365 9079 31399
rect 9597 31365 9631 31399
rect 9689 31365 9723 31399
rect 9827 31365 9861 31399
rect 16129 31365 16163 31399
rect 19257 31365 19291 31399
rect 26433 31365 26467 31399
rect 28089 31365 28123 31399
rect 31585 31365 31619 31399
rect 7573 31297 7607 31331
rect 7665 31297 7699 31331
rect 8309 31297 8343 31331
rect 8861 31297 8895 31331
rect 8953 31297 8987 31331
rect 9505 31297 9539 31331
rect 14841 31297 14875 31331
rect 14933 31297 14967 31331
rect 15301 31297 15335 31331
rect 15853 31297 15887 31331
rect 17049 31297 17083 31331
rect 19533 31297 19567 31331
rect 22201 31297 22235 31331
rect 23857 31297 23891 31331
rect 25237 31297 25271 31331
rect 26525 31297 26559 31331
rect 26985 31297 27019 31331
rect 27537 31297 27571 31331
rect 28825 31297 28859 31331
rect 29092 31297 29126 31331
rect 30757 31297 30791 31331
rect 32505 31297 32539 31331
rect 33793 31297 33827 31331
rect 34161 31297 34195 31331
rect 34713 31297 34747 31331
rect 39057 31297 39091 31331
rect 39313 31297 39347 31331
rect 39688 31297 39722 31331
rect 39948 31297 39982 31331
rect 41797 31297 41831 31331
rect 1409 31229 1443 31263
rect 1685 31229 1719 31263
rect 3157 31229 3191 31263
rect 3801 31229 3835 31263
rect 3985 31229 4019 31263
rect 4261 31229 4295 31263
rect 8033 31229 8067 31263
rect 9965 31229 9999 31263
rect 10241 31229 10275 31263
rect 10333 31229 10367 31263
rect 10425 31229 10459 31263
rect 10517 31229 10551 31263
rect 11621 31229 11655 31263
rect 11897 31229 11931 31263
rect 13369 31229 13403 31263
rect 14013 31229 14047 31263
rect 15117 31229 15151 31263
rect 16405 31229 16439 31263
rect 16865 31229 16899 31263
rect 21925 31229 21959 31263
rect 24041 31229 24075 31263
rect 25421 31229 25455 31263
rect 26617 31229 26651 31263
rect 28181 31229 28215 31263
rect 28365 31229 28399 31263
rect 31033 31229 31067 31263
rect 31677 31229 31711 31263
rect 31861 31229 31895 31263
rect 32781 31229 32815 31263
rect 33977 31229 34011 31263
rect 8125 31161 8159 31195
rect 8677 31161 8711 31195
rect 9229 31161 9263 31195
rect 10057 31161 10091 31195
rect 13461 31161 13495 31195
rect 3249 31093 3283 31127
rect 5733 31093 5767 31127
rect 17417 31093 17451 31127
rect 22569 31093 22603 31127
rect 23489 31093 23523 31127
rect 27721 31093 27755 31127
rect 30205 31093 30239 31127
rect 37933 31093 37967 31127
rect 41245 31093 41279 31127
rect 1777 30889 1811 30923
rect 1961 30889 1995 30923
rect 4353 30889 4387 30923
rect 7849 30889 7883 30923
rect 10701 30889 10735 30923
rect 12633 30889 12667 30923
rect 17049 30889 17083 30923
rect 22109 30889 22143 30923
rect 23857 30889 23891 30923
rect 27721 30889 27755 30923
rect 28457 30889 28491 30923
rect 29561 30889 29595 30923
rect 31953 30889 31987 30923
rect 35265 30889 35299 30923
rect 39221 30889 39255 30923
rect 42165 30889 42199 30923
rect 5641 30821 5675 30855
rect 18337 30821 18371 30855
rect 2053 30753 2087 30787
rect 2881 30753 2915 30787
rect 3065 30753 3099 30787
rect 3157 30753 3191 30787
rect 3893 30753 3927 30787
rect 3985 30753 4019 30787
rect 8953 30753 8987 30787
rect 13277 30753 13311 30787
rect 17509 30753 17543 30787
rect 19901 30753 19935 30787
rect 22293 30753 22327 30787
rect 25789 30753 25823 30787
rect 28273 30753 28307 30787
rect 29009 30753 29043 30787
rect 30205 30753 30239 30787
rect 30941 30753 30975 30787
rect 31309 30753 31343 30787
rect 32045 30753 32079 30787
rect 35725 30753 35759 30787
rect 2237 30685 2271 30719
rect 2697 30685 2731 30719
rect 3249 30685 3283 30719
rect 3341 30685 3375 30719
rect 4077 30685 4111 30719
rect 4169 30685 4203 30719
rect 4905 30685 4939 30719
rect 5089 30685 5123 30719
rect 5549 30685 5583 30719
rect 5825 30685 5859 30719
rect 6193 30685 6227 30719
rect 7757 30685 7791 30719
rect 7941 30685 7975 30719
rect 8493 30685 8527 30719
rect 8769 30685 8803 30719
rect 13001 30685 13035 30719
rect 13461 30685 13495 30719
rect 13645 30685 13679 30719
rect 17233 30685 17267 30719
rect 17325 30685 17359 30719
rect 17601 30685 17635 30719
rect 18521 30685 18555 30719
rect 18613 30685 18647 30719
rect 18705 30685 18739 30719
rect 18889 30685 18923 30719
rect 20085 30685 20119 30719
rect 20178 30685 20212 30719
rect 20361 30685 20395 30719
rect 20453 30685 20487 30719
rect 20550 30685 20584 30719
rect 21557 30685 21591 30719
rect 21925 30685 21959 30719
rect 23305 30685 23339 30719
rect 23489 30685 23523 30719
rect 23581 30685 23615 30719
rect 23673 30685 23707 30719
rect 35449 30685 35483 30719
rect 35541 30685 35575 30719
rect 35817 30685 35851 30719
rect 37841 30685 37875 30719
rect 39865 30685 39899 30719
rect 39957 30685 39991 30719
rect 40141 30685 40175 30719
rect 40417 30685 40451 30719
rect 1823 30651 1857 30685
rect 1593 30617 1627 30651
rect 2329 30617 2363 30651
rect 2421 30617 2455 30651
rect 2559 30617 2593 30651
rect 6285 30617 6319 30651
rect 8585 30617 8619 30651
rect 9229 30617 9263 30651
rect 18153 30617 18187 30651
rect 21741 30617 21775 30651
rect 21833 30617 21867 30651
rect 22569 30617 22603 30651
rect 26065 30617 26099 30651
rect 29929 30617 29963 30651
rect 32321 30617 32355 30651
rect 38108 30617 38142 30651
rect 40693 30617 40727 30651
rect 5181 30549 5215 30583
rect 6009 30549 6043 30583
rect 8677 30549 8711 30583
rect 13093 30549 13127 30583
rect 13553 30549 13587 30583
rect 17877 30549 17911 30583
rect 19257 30549 19291 30583
rect 19625 30549 19659 30583
rect 19717 30549 19751 30583
rect 20729 30549 20763 30583
rect 27537 30549 27571 30583
rect 30021 30549 30055 30583
rect 30389 30549 30423 30583
rect 33793 30549 33827 30583
rect 40325 30549 40359 30583
rect 2421 30345 2455 30379
rect 5825 30345 5859 30379
rect 8861 30345 8895 30379
rect 16497 30345 16531 30379
rect 17417 30345 17451 30379
rect 32505 30345 32539 30379
rect 35081 30345 35115 30379
rect 35541 30345 35575 30379
rect 38209 30345 38243 30379
rect 40141 30345 40175 30379
rect 40509 30345 40543 30379
rect 40969 30345 41003 30379
rect 41429 30345 41463 30379
rect 3249 30277 3283 30311
rect 3341 30277 3375 30311
rect 4629 30277 4663 30311
rect 5457 30277 5491 30311
rect 9137 30277 9171 30311
rect 19533 30277 19567 30311
rect 20177 30277 20211 30311
rect 22109 30277 22143 30311
rect 26249 30277 26283 30311
rect 34697 30277 34731 30311
rect 34897 30277 34931 30311
rect 35817 30277 35851 30311
rect 39129 30277 39163 30311
rect 40601 30277 40635 30311
rect 2605 30209 2639 30243
rect 2789 30209 2823 30243
rect 2881 30209 2915 30243
rect 3157 30209 3191 30243
rect 4077 30209 4111 30243
rect 5365 30209 5399 30243
rect 6561 30209 6595 30243
rect 6837 30209 6871 30243
rect 9045 30209 9079 30243
rect 9229 30209 9263 30243
rect 9347 30209 9381 30243
rect 10425 30209 10459 30243
rect 11621 30209 11655 30243
rect 13553 30209 13587 30243
rect 13645 30209 13679 30243
rect 14013 30209 14047 30243
rect 14749 30209 14783 30243
rect 17233 30209 17267 30243
rect 17601 30209 17635 30243
rect 17693 30209 17727 30243
rect 17969 30209 18003 30243
rect 18521 30209 18555 30243
rect 18797 30209 18831 30243
rect 19165 30209 19199 30243
rect 19258 30209 19292 30243
rect 19441 30209 19475 30243
rect 19630 30209 19664 30243
rect 19901 30209 19935 30243
rect 20085 30209 20119 30243
rect 20269 30209 20303 30243
rect 21281 30209 21315 30243
rect 21373 30209 21407 30243
rect 21649 30209 21683 30243
rect 22012 30209 22046 30243
rect 22201 30209 22235 30243
rect 22329 30209 22363 30243
rect 22477 30209 22511 30243
rect 26433 30209 26467 30243
rect 26525 30209 26559 30243
rect 26801 30209 26835 30243
rect 31677 30209 31711 30243
rect 32689 30209 32723 30243
rect 32781 30209 32815 30243
rect 33057 30209 33091 30243
rect 34989 30209 35023 30243
rect 35173 30209 35207 30243
rect 35720 30209 35754 30243
rect 35909 30209 35943 30243
rect 36037 30209 36071 30243
rect 36185 30209 36219 30243
rect 36277 30209 36311 30243
rect 36461 30209 36495 30243
rect 36553 30209 36587 30243
rect 36645 30209 36679 30243
rect 37289 30209 37323 30243
rect 37437 30209 37471 30243
rect 37565 30209 37599 30243
rect 37657 30209 37691 30243
rect 37795 30209 37829 30243
rect 38577 30209 38611 30243
rect 41337 30209 41371 30243
rect 41797 30209 41831 30243
rect 2973 30141 3007 30175
rect 5641 30141 5675 30175
rect 5733 30141 5767 30175
rect 6009 30141 6043 30175
rect 6101 30141 6135 30175
rect 9505 30141 9539 30175
rect 9873 30141 9907 30175
rect 11897 30141 11931 30175
rect 15025 30141 15059 30175
rect 21557 30141 21591 30175
rect 23213 30141 23247 30175
rect 24685 30141 24719 30175
rect 24961 30141 24995 30175
rect 38669 30141 38703 30175
rect 38853 30141 38887 30175
rect 39957 30141 39991 30175
rect 40693 30141 40727 30175
rect 41521 30141 41555 30175
rect 3525 30073 3559 30107
rect 6653 30073 6687 30107
rect 6745 30073 6779 30107
rect 18705 30073 18739 30107
rect 19809 30073 19843 30107
rect 20453 30073 20487 30107
rect 21833 30073 21867 30107
rect 36829 30073 36863 30107
rect 3893 30005 3927 30039
rect 6377 30005 6411 30039
rect 13369 30005 13403 30039
rect 14013 30005 14047 30039
rect 14197 30005 14231 30039
rect 16681 30005 16715 30039
rect 17877 30005 17911 30039
rect 18337 30005 18371 30039
rect 21097 30005 21131 30039
rect 26709 30005 26743 30039
rect 32965 30005 32999 30039
rect 34529 30005 34563 30039
rect 34713 30005 34747 30039
rect 37933 30005 37967 30039
rect 41981 30005 42015 30039
rect 5365 29801 5399 29835
rect 9597 29801 9631 29835
rect 13093 29801 13127 29835
rect 16313 29801 16347 29835
rect 19257 29801 19291 29835
rect 19717 29801 19751 29835
rect 19901 29801 19935 29835
rect 21176 29801 21210 29835
rect 22661 29801 22695 29835
rect 24961 29801 24995 29835
rect 26157 29801 26191 29835
rect 26801 29801 26835 29835
rect 29285 29801 29319 29835
rect 30021 29801 30055 29835
rect 32965 29801 32999 29835
rect 33701 29801 33735 29835
rect 33885 29801 33919 29835
rect 34897 29801 34931 29835
rect 38945 29801 38979 29835
rect 40325 29801 40359 29835
rect 42165 29801 42199 29835
rect 13001 29733 13035 29767
rect 16589 29733 16623 29767
rect 19073 29733 19107 29767
rect 23949 29733 23983 29767
rect 34253 29733 34287 29767
rect 35633 29733 35667 29767
rect 36369 29733 36403 29767
rect 37289 29733 37323 29767
rect 4077 29665 4111 29699
rect 4169 29665 4203 29699
rect 5917 29665 5951 29699
rect 6377 29665 6411 29699
rect 6653 29665 6687 29699
rect 11253 29665 11287 29699
rect 14657 29665 14691 29699
rect 14841 29665 14875 29699
rect 16773 29665 16807 29699
rect 17141 29665 17175 29699
rect 18061 29665 18095 29699
rect 20913 29665 20947 29699
rect 24501 29665 24535 29699
rect 25697 29665 25731 29699
rect 25881 29665 25915 29699
rect 26617 29665 26651 29699
rect 30481 29665 30515 29699
rect 31861 29665 31895 29699
rect 32597 29665 32631 29699
rect 32781 29665 32815 29699
rect 34805 29665 34839 29699
rect 34989 29665 35023 29699
rect 39497 29665 39531 29699
rect 40693 29665 40727 29699
rect 2789 29597 2823 29631
rect 3065 29597 3099 29631
rect 3433 29597 3467 29631
rect 3985 29597 4019 29631
rect 4261 29597 4295 29631
rect 4721 29597 4755 29631
rect 4905 29597 4939 29631
rect 4997 29597 5031 29631
rect 5089 29597 5123 29631
rect 5641 29597 5675 29631
rect 5733 29597 5767 29631
rect 6285 29597 6319 29631
rect 9781 29597 9815 29631
rect 10057 29597 10091 29631
rect 13277 29597 13311 29631
rect 13369 29597 13403 29631
rect 14105 29597 14139 29631
rect 15209 29597 15243 29631
rect 16497 29597 16531 29631
rect 16681 29597 16715 29631
rect 16957 29597 16991 29631
rect 17325 29597 17359 29631
rect 18337 29597 18371 29631
rect 18521 29597 18555 29631
rect 18889 29597 18923 29631
rect 19441 29597 19475 29631
rect 19625 29597 19659 29631
rect 20269 29597 20303 29631
rect 20637 29597 20671 29631
rect 23305 29597 23339 29631
rect 23453 29597 23487 29631
rect 23673 29597 23707 29631
rect 23770 29597 23804 29631
rect 24409 29597 24443 29631
rect 24685 29597 24719 29631
rect 24777 29597 24811 29631
rect 25605 29597 25639 29631
rect 26341 29597 26375 29631
rect 26433 29597 26467 29631
rect 26709 29597 26743 29631
rect 26985 29597 27019 29631
rect 27077 29597 27111 29631
rect 27353 29597 27387 29631
rect 27445 29597 27479 29631
rect 27629 29597 27663 29631
rect 29561 29597 29595 29631
rect 29745 29597 29779 29631
rect 29837 29597 29871 29631
rect 30113 29597 30147 29631
rect 30205 29597 30239 29631
rect 30297 29597 30331 29631
rect 31125 29597 31159 29631
rect 33144 29597 33178 29631
rect 33241 29597 33275 29631
rect 33333 29597 33367 29631
rect 33461 29597 33495 29631
rect 33609 29597 33643 29631
rect 34713 29597 34747 29631
rect 35081 29597 35115 29631
rect 35265 29597 35299 29631
rect 35357 29597 35391 29631
rect 35449 29597 35483 29631
rect 35725 29597 35759 29631
rect 35818 29597 35852 29631
rect 36231 29597 36265 29631
rect 36645 29597 36679 29631
rect 36738 29597 36772 29631
rect 36921 29597 36955 29631
rect 37013 29597 37047 29631
rect 37151 29597 37185 29631
rect 39865 29597 39899 29631
rect 40141 29597 40175 29631
rect 40417 29597 40451 29631
rect 2605 29529 2639 29563
rect 3157 29529 3191 29563
rect 3249 29529 3283 29563
rect 6561 29529 6595 29563
rect 6929 29529 6963 29563
rect 9965 29529 9999 29563
rect 11529 29529 11563 29563
rect 15117 29529 15151 29563
rect 18705 29529 18739 29563
rect 18797 29529 18831 29563
rect 23581 29529 23615 29563
rect 27169 29529 27203 29563
rect 29193 29529 29227 29563
rect 33885 29529 33919 29563
rect 36001 29529 36035 29563
rect 36093 29529 36127 29563
rect 39957 29529 39991 29563
rect 2421 29461 2455 29495
rect 2881 29461 2915 29495
rect 3801 29461 3835 29495
rect 5549 29461 5583 29495
rect 8401 29461 8435 29495
rect 13737 29461 13771 29495
rect 15025 29461 15059 29495
rect 15393 29461 15427 29495
rect 17417 29461 17451 29495
rect 17785 29461 17819 29495
rect 19901 29461 19935 29495
rect 20453 29461 20487 29495
rect 25881 29461 25915 29495
rect 27537 29461 27571 29495
rect 30481 29461 30515 29495
rect 32137 29461 32171 29495
rect 32505 29461 32539 29495
rect 4813 29257 4847 29291
rect 5549 29257 5583 29291
rect 6377 29257 6411 29291
rect 12081 29257 12115 29291
rect 13645 29257 13679 29291
rect 17049 29257 17083 29291
rect 17417 29257 17451 29291
rect 18337 29257 18371 29291
rect 19993 29257 20027 29291
rect 24041 29257 24075 29291
rect 25973 29257 26007 29291
rect 26151 29257 26185 29291
rect 27077 29257 27111 29291
rect 31217 29257 31251 29291
rect 31401 29257 31435 29291
rect 33057 29257 33091 29291
rect 41337 29257 41371 29291
rect 2421 29189 2455 29223
rect 2559 29189 2593 29223
rect 3525 29189 3559 29223
rect 4445 29189 4479 29223
rect 5917 29189 5951 29223
rect 17233 29189 17267 29223
rect 18521 29189 18555 29223
rect 19901 29189 19935 29223
rect 20821 29189 20855 29223
rect 23857 29189 23891 29223
rect 26617 29189 26651 29223
rect 27261 29189 27295 29223
rect 27813 29189 27847 29223
rect 27905 29189 27939 29223
rect 28549 29189 28583 29223
rect 30481 29189 30515 29223
rect 32505 29189 32539 29223
rect 34405 29189 34439 29223
rect 34621 29189 34655 29223
rect 35357 29189 35391 29223
rect 37565 29189 37599 29223
rect 1777 29121 1811 29155
rect 1961 29121 1995 29155
rect 2237 29121 2271 29155
rect 2329 29121 2363 29155
rect 3433 29121 3467 29155
rect 4169 29121 4203 29155
rect 4261 29121 4295 29155
rect 4629 29121 4663 29155
rect 4997 29121 5031 29155
rect 5089 29121 5123 29155
rect 5181 29121 5215 29155
rect 5299 29121 5333 29155
rect 5733 29121 5767 29155
rect 5825 29121 5859 29155
rect 6101 29121 6135 29155
rect 6745 29121 6779 29155
rect 7389 29121 7423 29155
rect 7481 29121 7515 29155
rect 12357 29121 12391 29155
rect 12817 29121 12851 29155
rect 13461 29121 13495 29155
rect 13553 29121 13587 29155
rect 13737 29121 13771 29155
rect 16957 29121 16991 29155
rect 17325 29121 17359 29155
rect 17601 29121 17635 29155
rect 18153 29121 18187 29155
rect 18429 29121 18463 29155
rect 18613 29121 18647 29155
rect 19625 29121 19659 29155
rect 19809 29121 19843 29155
rect 20729 29121 20763 29155
rect 21097 29121 21131 29155
rect 21189 29121 21223 29155
rect 21373 29121 21407 29155
rect 21465 29121 21499 29155
rect 21833 29121 21867 29155
rect 21996 29121 22030 29155
rect 22109 29121 22143 29155
rect 22201 29121 22235 29155
rect 22845 29121 22879 29155
rect 22937 29121 22971 29155
rect 23121 29121 23155 29155
rect 23213 29121 23247 29155
rect 24133 29121 24167 29155
rect 24317 29121 24351 29155
rect 25237 29121 25271 29155
rect 25513 29121 25547 29155
rect 26065 29121 26099 29155
rect 26525 29121 26559 29155
rect 26985 29121 27019 29155
rect 27629 29121 27663 29155
rect 27997 29121 28031 29155
rect 28273 29121 28307 29155
rect 30113 29121 30147 29155
rect 30297 29121 30331 29155
rect 30573 29121 30607 29155
rect 30757 29121 30791 29155
rect 31033 29121 31067 29155
rect 31125 29121 31159 29155
rect 31677 29121 31711 29155
rect 31861 29121 31895 29155
rect 32137 29121 32171 29155
rect 32230 29121 32264 29155
rect 32413 29121 32447 29155
rect 32643 29121 32677 29155
rect 32873 29121 32907 29155
rect 33701 29121 33735 29155
rect 33793 29121 33827 29155
rect 33885 29121 33919 29155
rect 35173 29121 35207 29155
rect 35449 29121 35483 29155
rect 35817 29121 35851 29155
rect 36093 29121 36127 29155
rect 36185 29121 36219 29155
rect 39681 29121 39715 29155
rect 40325 29121 40359 29155
rect 41889 29121 41923 29155
rect 1869 29053 1903 29087
rect 2697 29053 2731 29087
rect 2789 29053 2823 29087
rect 5457 29053 5491 29087
rect 6653 29053 6687 29087
rect 9505 29053 9539 29087
rect 9781 29053 9815 29087
rect 12265 29053 12299 29087
rect 12725 29053 12759 29087
rect 17877 29053 17911 29087
rect 19211 29053 19245 29087
rect 19533 29053 19567 29087
rect 20177 29053 20211 29087
rect 24501 29053 24535 29087
rect 25329 29053 25363 29087
rect 25697 29053 25731 29087
rect 30021 29053 30055 29087
rect 30849 29053 30883 29087
rect 31493 29053 31527 29087
rect 33977 29053 34011 29087
rect 36369 29053 36403 29087
rect 37289 29053 37323 29087
rect 40877 29053 40911 29087
rect 41429 29053 41463 29087
rect 41521 29053 41555 29087
rect 11253 28985 11287 29019
rect 17233 28985 17267 29019
rect 17601 28985 17635 29019
rect 23489 28985 23523 29019
rect 25421 28985 25455 29019
rect 25789 28985 25823 29019
rect 28181 28985 28215 29019
rect 30573 28985 30607 29019
rect 34161 28985 34195 29019
rect 34253 28985 34287 29019
rect 35909 28985 35943 29019
rect 39037 28985 39071 29019
rect 40969 28985 41003 29019
rect 42073 28985 42107 29019
rect 2053 28917 2087 28951
rect 17969 28917 18003 28951
rect 21649 28917 21683 28951
rect 22477 28917 22511 28951
rect 23397 28917 23431 28951
rect 23857 28917 23891 28951
rect 25053 28917 25087 28951
rect 26433 28917 26467 28951
rect 27261 28917 27295 28951
rect 32781 28917 32815 28951
rect 34437 28917 34471 28951
rect 34989 28917 35023 28951
rect 3157 28713 3191 28747
rect 4721 28713 4755 28747
rect 4905 28713 4939 28747
rect 6101 28713 6135 28747
rect 6469 28713 6503 28747
rect 8217 28713 8251 28747
rect 13185 28713 13219 28747
rect 13921 28713 13955 28747
rect 18061 28713 18095 28747
rect 19257 28713 19291 28747
rect 21281 28713 21315 28747
rect 21465 28713 21499 28747
rect 22293 28713 22327 28747
rect 22569 28713 22603 28747
rect 22845 28713 22879 28747
rect 23673 28713 23707 28747
rect 25697 28713 25731 28747
rect 30205 28713 30239 28747
rect 30665 28713 30699 28747
rect 31033 28713 31067 28747
rect 34437 28713 34471 28747
rect 35173 28713 35207 28747
rect 36093 28713 36127 28747
rect 42165 28713 42199 28747
rect 3341 28645 3375 28679
rect 3801 28645 3835 28679
rect 10977 28645 11011 28679
rect 12725 28645 12759 28679
rect 14289 28645 14323 28679
rect 18889 28645 18923 28679
rect 21097 28645 21131 28679
rect 27169 28645 27203 28679
rect 31217 28645 31251 28679
rect 31401 28645 31435 28679
rect 35633 28645 35667 28679
rect 1409 28577 1443 28611
rect 1685 28577 1719 28611
rect 4077 28577 4111 28611
rect 9229 28577 9263 28611
rect 14933 28577 14967 28611
rect 18705 28577 18739 28611
rect 26341 28577 26375 28611
rect 30763 28577 30797 28611
rect 31309 28577 31343 28611
rect 34069 28577 34103 28611
rect 34805 28577 34839 28611
rect 35449 28577 35483 28611
rect 37933 28577 37967 28611
rect 40693 28577 40727 28611
rect 3525 28509 3559 28543
rect 4169 28509 4203 28543
rect 4537 28509 4571 28543
rect 4721 28509 4755 28543
rect 5089 28509 5123 28543
rect 5181 28509 5215 28543
rect 5457 28509 5491 28543
rect 6101 28509 6135 28543
rect 6285 28509 6319 28543
rect 7665 28509 7699 28543
rect 11529 28509 11563 28543
rect 13093 28509 13127 28543
rect 13277 28509 13311 28543
rect 13737 28509 13771 28543
rect 13921 28509 13955 28543
rect 14289 28509 14323 28543
rect 14565 28509 14599 28543
rect 14657 28509 14691 28543
rect 18245 28509 18279 28543
rect 18429 28509 18463 28543
rect 19073 28509 19107 28543
rect 19441 28509 19475 28543
rect 21005 28509 21039 28543
rect 21189 28509 21223 28543
rect 21833 28509 21867 28543
rect 22477 28509 22511 28543
rect 22753 28509 22787 28543
rect 22937 28509 22971 28543
rect 23029 28509 23063 28543
rect 23213 28509 23247 28543
rect 23305 28509 23339 28543
rect 23397 28509 23431 28543
rect 23949 28509 23983 28543
rect 25881 28509 25915 28543
rect 26157 28509 26191 28543
rect 26525 28509 26559 28543
rect 27077 28509 27111 28543
rect 29561 28509 29595 28543
rect 29654 28509 29688 28543
rect 29929 28509 29963 28543
rect 30026 28509 30060 28543
rect 30297 28509 30331 28543
rect 30481 28509 30515 28543
rect 31585 28509 31619 28543
rect 31861 28509 31895 28543
rect 32045 28509 32079 28543
rect 34253 28509 34287 28543
rect 35725 28509 35759 28543
rect 35817 28509 35851 28543
rect 35909 28509 35943 28543
rect 37657 28509 37691 28543
rect 40417 28509 40451 28543
rect 5273 28441 5307 28475
rect 9505 28441 9539 28475
rect 12357 28441 12391 28475
rect 12909 28441 12943 28475
rect 15209 28441 15243 28475
rect 16957 28441 16991 28475
rect 18337 28441 18371 28475
rect 18567 28441 18601 28475
rect 19625 28441 19659 28475
rect 21465 28441 21499 28475
rect 21925 28441 21959 28475
rect 22109 28441 22143 28475
rect 23765 28441 23799 28475
rect 24133 28441 24167 28475
rect 26617 28441 26651 28475
rect 27353 28441 27387 28475
rect 29193 28441 29227 28475
rect 29377 28441 29411 28475
rect 29837 28441 29871 28475
rect 30849 28441 30883 28475
rect 31049 28441 31083 28475
rect 31953 28441 31987 28475
rect 35173 28441 35207 28475
rect 35449 28441 35483 28475
rect 36093 28441 36127 28475
rect 37841 28441 37875 28475
rect 38209 28441 38243 28475
rect 14473 28373 14507 28407
rect 14749 28373 14783 28407
rect 26065 28373 26099 28407
rect 26985 28373 27019 28407
rect 27077 28373 27111 28407
rect 31769 28373 31803 28407
rect 35357 28373 35391 28407
rect 37473 28373 37507 28407
rect 39681 28373 39715 28407
rect 3709 28169 3743 28203
rect 5273 28169 5307 28203
rect 10517 28169 10551 28203
rect 10885 28169 10919 28203
rect 10977 28169 11011 28203
rect 11529 28169 11563 28203
rect 11989 28169 12023 28203
rect 15025 28169 15059 28203
rect 18521 28169 18555 28203
rect 19993 28169 20027 28203
rect 28641 28169 28675 28203
rect 29009 28169 29043 28203
rect 29653 28169 29687 28203
rect 30941 28169 30975 28203
rect 37749 28169 37783 28203
rect 38301 28169 38335 28203
rect 39681 28169 39715 28203
rect 39773 28169 39807 28203
rect 12541 28101 12575 28135
rect 14657 28101 14691 28135
rect 14857 28101 14891 28135
rect 18889 28101 18923 28135
rect 25513 28101 25547 28135
rect 34253 28101 34287 28135
rect 34437 28101 34471 28135
rect 38577 28101 38611 28135
rect 1685 28033 1719 28067
rect 5181 28033 5215 28067
rect 5549 28033 5583 28067
rect 5641 28033 5675 28067
rect 8686 28033 8720 28067
rect 8953 28033 8987 28067
rect 10158 28033 10192 28067
rect 11897 28033 11931 28067
rect 12449 28033 12483 28067
rect 12633 28033 12667 28067
rect 15393 28033 15427 28067
rect 18337 28033 18371 28067
rect 18797 28033 18831 28067
rect 18981 28033 19015 28067
rect 19901 28033 19935 28067
rect 20085 28033 20119 28067
rect 23581 28033 23615 28067
rect 23765 28033 23799 28067
rect 24777 28033 24811 28067
rect 24869 28033 24903 28067
rect 25145 28033 25179 28067
rect 25421 28033 25455 28067
rect 25605 28033 25639 28067
rect 25789 28033 25823 28067
rect 27721 28033 27755 28067
rect 27814 28033 27848 28067
rect 27997 28033 28031 28067
rect 28089 28033 28123 28067
rect 28186 28033 28220 28067
rect 28457 28033 28491 28067
rect 28825 28033 28859 28067
rect 29745 28033 29779 28067
rect 30205 28033 30239 28067
rect 30389 28033 30423 28067
rect 30481 28033 30515 28067
rect 30573 28033 30607 28067
rect 30849 28033 30883 28067
rect 31033 28033 31067 28067
rect 32321 28033 32355 28067
rect 32413 28033 32447 28067
rect 32689 28033 32723 28067
rect 33701 28033 33735 28067
rect 33977 28033 34011 28067
rect 37841 28033 37875 28067
rect 38485 28033 38519 28067
rect 38669 28033 38703 28067
rect 38853 28033 38887 28067
rect 39037 28033 39071 28067
rect 40233 28033 40267 28067
rect 40417 28033 40451 28067
rect 41521 28033 41555 28067
rect 41889 28033 41923 28067
rect 1961 27965 1995 27999
rect 2237 27965 2271 27999
rect 5273 27965 5307 27999
rect 10425 27965 10459 27999
rect 11069 27965 11103 27999
rect 12081 27965 12115 27999
rect 12725 27965 12759 27999
rect 13001 27965 13035 27999
rect 18153 27965 18187 27999
rect 29561 27965 29595 27999
rect 37565 27965 37599 27999
rect 39497 27965 39531 27999
rect 23765 27897 23799 27931
rect 25237 27897 25271 27931
rect 28365 27897 28399 27931
rect 30757 27897 30791 27931
rect 41705 27897 41739 27931
rect 1501 27829 1535 27863
rect 4997 27829 5031 27863
rect 5457 27829 5491 27863
rect 5733 27829 5767 27863
rect 7573 27829 7607 27863
rect 9045 27829 9079 27863
rect 14473 27829 14507 27863
rect 14841 27829 14875 27863
rect 15209 27829 15243 27863
rect 24593 27829 24627 27863
rect 25053 27829 25087 27863
rect 30113 27829 30147 27863
rect 32137 27829 32171 27863
rect 32597 27829 32631 27863
rect 33793 27829 33827 27863
rect 34161 27829 34195 27863
rect 34621 27829 34655 27863
rect 38209 27829 38243 27863
rect 39129 27829 39163 27863
rect 40141 27829 40175 27863
rect 40601 27829 40635 27863
rect 42073 27829 42107 27863
rect 14933 27625 14967 27659
rect 17141 27625 17175 27659
rect 19533 27625 19567 27659
rect 21741 27625 21775 27659
rect 24666 27625 24700 27659
rect 26157 27625 26191 27659
rect 31940 27625 31974 27659
rect 37749 27625 37783 27659
rect 40404 27625 40438 27659
rect 41889 27625 41923 27659
rect 4629 27557 4663 27591
rect 7665 27557 7699 27591
rect 8401 27557 8435 27591
rect 12909 27557 12943 27591
rect 14473 27557 14507 27591
rect 15301 27557 15335 27591
rect 17785 27557 17819 27591
rect 19901 27557 19935 27591
rect 19993 27557 20027 27591
rect 22017 27557 22051 27591
rect 26341 27557 26375 27591
rect 26801 27557 26835 27591
rect 33425 27557 33459 27591
rect 33517 27557 33551 27591
rect 39129 27557 39163 27591
rect 4997 27489 5031 27523
rect 7757 27489 7791 27523
rect 9045 27489 9079 27523
rect 10885 27489 10919 27523
rect 15393 27489 15427 27523
rect 19809 27489 19843 27523
rect 23029 27489 23063 27523
rect 24409 27489 24443 27523
rect 28549 27489 28583 27523
rect 29101 27489 29135 27523
rect 31677 27489 31711 27523
rect 34897 27489 34931 27523
rect 35081 27489 35115 27523
rect 35449 27489 35483 27523
rect 4629 27421 4663 27455
rect 4905 27421 4939 27455
rect 7113 27421 7147 27455
rect 7389 27421 7423 27455
rect 7481 27421 7515 27455
rect 7915 27421 7949 27455
rect 8217 27421 8251 27455
rect 9781 27421 9815 27455
rect 12725 27421 12759 27455
rect 14657 27421 14691 27455
rect 14749 27421 14783 27455
rect 15025 27421 15059 27455
rect 17509 27421 17543 27455
rect 18061 27421 18095 27455
rect 18153 27421 18187 27455
rect 18337 27421 18371 27455
rect 18429 27421 18463 27455
rect 18613 27421 18647 27455
rect 20361 27421 20395 27455
rect 20545 27421 20579 27455
rect 20637 27421 20671 27455
rect 21557 27421 21591 27455
rect 21741 27421 21775 27455
rect 21833 27421 21867 27455
rect 22017 27421 22051 27455
rect 22109 27421 22143 27455
rect 22477 27421 22511 27455
rect 24041 27421 24075 27455
rect 26525 27421 26559 27455
rect 28825 27421 28859 27455
rect 28917 27421 28951 27455
rect 29193 27421 29227 27455
rect 30665 27421 30699 27455
rect 30757 27421 30791 27455
rect 30941 27421 30975 27455
rect 31043 27399 31077 27433
rect 33655 27421 33689 27455
rect 33793 27421 33827 27455
rect 33885 27421 33919 27455
rect 34013 27421 34047 27455
rect 34161 27421 34195 27455
rect 34253 27421 34287 27455
rect 34437 27421 34471 27455
rect 34989 27421 35023 27455
rect 35173 27421 35207 27455
rect 35357 27421 35391 27455
rect 35633 27421 35667 27455
rect 35725 27421 35759 27455
rect 36001 27421 36035 27455
rect 39313 27421 39347 27455
rect 39681 27421 39715 27455
rect 40141 27421 40175 27455
rect 5273 27353 5307 27387
rect 7297 27353 7331 27387
rect 8033 27353 8067 27387
rect 8125 27353 8159 27387
rect 9689 27353 9723 27387
rect 11161 27353 11195 27387
rect 14933 27353 14967 27387
rect 15301 27353 15335 27387
rect 15669 27353 15703 27387
rect 17325 27353 17359 27387
rect 17693 27353 17727 27387
rect 17785 27353 17819 27387
rect 22661 27353 22695 27387
rect 22845 27353 22879 27387
rect 28273 27353 28307 27387
rect 28641 27353 28675 27387
rect 31493 27353 31527 27387
rect 34345 27353 34379 27387
rect 35909 27353 35943 27387
rect 36277 27353 36311 27387
rect 39405 27353 39439 27387
rect 39497 27353 39531 27387
rect 6745 27285 6779 27319
rect 10425 27285 10459 27319
rect 12633 27285 12667 27319
rect 15117 27285 15151 27319
rect 17969 27285 18003 27319
rect 18153 27285 18187 27319
rect 18521 27285 18555 27319
rect 30481 27285 30515 27319
rect 31217 27285 31251 27319
rect 34713 27285 34747 27319
rect 5457 27081 5491 27115
rect 6469 27081 6503 27115
rect 9321 27081 9355 27115
rect 11529 27081 11563 27115
rect 11989 27081 12023 27115
rect 15025 27081 15059 27115
rect 15485 27081 15519 27115
rect 16313 27081 16347 27115
rect 16865 27081 16899 27115
rect 17325 27081 17359 27115
rect 19809 27081 19843 27115
rect 20821 27081 20855 27115
rect 22861 27081 22895 27115
rect 23029 27081 23063 27115
rect 25513 27081 25547 27115
rect 28181 27081 28215 27115
rect 33149 27081 33183 27115
rect 36645 27081 36679 27115
rect 40049 27081 40083 27115
rect 40141 27081 40175 27115
rect 5089 27013 5123 27047
rect 5273 27013 5307 27047
rect 6745 27013 6779 27047
rect 9137 27013 9171 27047
rect 14657 27013 14691 27047
rect 14841 27013 14875 27047
rect 16405 27013 16439 27047
rect 18061 27013 18095 27047
rect 19993 27013 20027 27047
rect 20729 27013 20763 27047
rect 22661 27013 22695 27047
rect 24133 27013 24167 27047
rect 34621 27013 34655 27047
rect 35541 27013 35575 27047
rect 38393 27013 38427 27047
rect 38485 27013 38519 27047
rect 4169 26945 4203 26979
rect 4353 26945 4387 26979
rect 4629 26945 4663 26979
rect 4721 26945 4755 26979
rect 4905 26945 4939 26979
rect 4997 26945 5031 26979
rect 8953 26945 8987 26979
rect 10526 26945 10560 26979
rect 10793 26945 10827 26979
rect 11897 26945 11931 26979
rect 15117 26945 15151 26979
rect 17785 26945 17819 26979
rect 17969 26945 18003 26979
rect 18245 26945 18279 26979
rect 18429 26945 18463 26979
rect 18981 26945 19015 26979
rect 19349 26945 19383 26979
rect 19901 26945 19935 26979
rect 20453 26945 20487 26979
rect 20637 26945 20671 26979
rect 23397 26945 23431 26979
rect 25605 26945 25639 26979
rect 26157 26945 26191 26979
rect 26341 26945 26375 26979
rect 26433 26945 26467 26979
rect 26525 26945 26559 26979
rect 28273 26945 28307 26979
rect 28733 26945 28767 26979
rect 28917 26945 28951 26979
rect 29009 26945 29043 26979
rect 29101 26945 29135 26979
rect 29929 26945 29963 26979
rect 34897 26945 34931 26979
rect 35403 26945 35437 26979
rect 35633 26945 35667 26979
rect 35816 26945 35850 26979
rect 35909 26945 35943 26979
rect 36001 26945 36035 26979
rect 36149 26945 36183 26979
rect 36277 26945 36311 26979
rect 36369 26945 36403 26979
rect 36466 26945 36500 26979
rect 40601 26945 40635 26979
rect 40785 26945 40819 26979
rect 41889 26945 41923 26979
rect 2421 26877 2455 26911
rect 4261 26877 4295 26911
rect 12081 26877 12115 26911
rect 15209 26877 15243 26911
rect 16681 26877 16715 26911
rect 16773 26877 16807 26911
rect 17049 26877 17083 26911
rect 17141 26877 17175 26911
rect 19441 26877 19475 26911
rect 19625 26877 19659 26911
rect 20361 26877 20395 26911
rect 21005 26877 21039 26911
rect 25329 26877 25363 26911
rect 28089 26877 28123 26911
rect 32137 26877 32171 26911
rect 32413 26877 32447 26911
rect 38209 26877 38243 26911
rect 39865 26877 39899 26911
rect 4445 26809 4479 26843
rect 18245 26809 18279 26843
rect 35265 26809 35299 26843
rect 40509 26809 40543 26843
rect 2973 26741 3007 26775
rect 9413 26741 9447 26775
rect 15117 26741 15151 26775
rect 17601 26741 17635 26775
rect 18797 26741 18831 26775
rect 18981 26741 19015 26775
rect 22845 26741 22879 26775
rect 25973 26741 26007 26775
rect 26709 26741 26743 26775
rect 28641 26741 28675 26775
rect 29285 26741 29319 26775
rect 30192 26741 30226 26775
rect 31677 26741 31711 26775
rect 38853 26741 38887 26775
rect 40969 26741 41003 26775
rect 42073 26741 42107 26775
rect 3267 26537 3301 26571
rect 4445 26537 4479 26571
rect 4629 26537 4663 26571
rect 4905 26537 4939 26571
rect 9505 26537 9539 26571
rect 12081 26537 12115 26571
rect 15025 26537 15059 26571
rect 16497 26537 16531 26571
rect 18429 26537 18463 26571
rect 20821 26537 20855 26571
rect 30113 26537 30147 26571
rect 34161 26537 34195 26571
rect 35817 26537 35851 26571
rect 7941 26469 7975 26503
rect 8769 26469 8803 26503
rect 16957 26469 16991 26503
rect 23765 26469 23799 26503
rect 23949 26469 23983 26503
rect 31953 26469 31987 26503
rect 35449 26469 35483 26503
rect 36001 26469 36035 26503
rect 36645 26469 36679 26503
rect 37289 26469 37323 26503
rect 1501 26401 1535 26435
rect 10333 26401 10367 26435
rect 13645 26401 13679 26435
rect 13921 26401 13955 26435
rect 15393 26401 15427 26435
rect 15485 26401 15519 26435
rect 16681 26401 16715 26435
rect 17141 26401 17175 26435
rect 18245 26401 18279 26435
rect 19257 26401 19291 26435
rect 19717 26401 19751 26435
rect 19809 26401 19843 26435
rect 20913 26401 20947 26435
rect 23121 26401 23155 26435
rect 23581 26401 23615 26435
rect 24501 26401 24535 26435
rect 30573 26401 30607 26435
rect 34805 26401 34839 26435
rect 38393 26401 38427 26435
rect 40417 26401 40451 26435
rect 40693 26401 40727 26435
rect 42165 26401 42199 26435
rect 3525 26333 3559 26367
rect 4077 26333 4111 26367
rect 5084 26333 5118 26367
rect 5273 26333 5307 26367
rect 5456 26333 5490 26367
rect 5549 26333 5583 26367
rect 5733 26333 5767 26367
rect 5825 26333 5859 26367
rect 6193 26333 6227 26367
rect 6653 26333 6687 26367
rect 6929 26333 6963 26367
rect 7297 26333 7331 26367
rect 8033 26333 8067 26367
rect 8217 26333 8251 26367
rect 8401 26333 8435 26367
rect 8493 26333 8527 26367
rect 8585 26333 8619 26367
rect 8953 26333 8987 26367
rect 9137 26333 9171 26367
rect 9229 26333 9263 26367
rect 9321 26333 9355 26367
rect 9597 26333 9631 26367
rect 15301 26333 15335 26367
rect 15761 26333 15795 26367
rect 15853 26333 15887 26367
rect 15946 26333 15980 26367
rect 16221 26333 16255 26367
rect 16318 26333 16352 26367
rect 16589 26333 16623 26367
rect 16773 26333 16807 26367
rect 17233 26333 17267 26367
rect 17325 26333 17359 26367
rect 17417 26333 17451 26367
rect 17877 26333 17911 26367
rect 17969 26333 18003 26367
rect 18337 26333 18371 26367
rect 18521 26333 18555 26367
rect 20085 26333 20119 26367
rect 20821 26333 20855 26367
rect 21097 26333 21131 26367
rect 21465 26333 21499 26367
rect 21649 26333 21683 26367
rect 21741 26333 21775 26367
rect 21925 26333 21959 26367
rect 22477 26333 22511 26367
rect 23305 26333 23339 26367
rect 23489 26333 23523 26367
rect 23857 26333 23891 26367
rect 23949 26333 23983 26367
rect 24133 26333 24167 26367
rect 30297 26333 30331 26367
rect 30389 26333 30423 26367
rect 30665 26333 30699 26367
rect 31309 26333 31343 26367
rect 31457 26333 31491 26367
rect 31677 26333 31711 26367
rect 31774 26333 31808 26367
rect 33609 26333 33643 26367
rect 33885 26333 33919 26367
rect 33977 26333 34011 26367
rect 34989 26333 35023 26367
rect 36093 26333 36127 26367
rect 36369 26333 36403 26367
rect 36461 26333 36495 26367
rect 36737 26333 36771 26367
rect 36921 26333 36955 26367
rect 37013 26333 37047 26367
rect 37105 26333 37139 26367
rect 37381 26333 37415 26367
rect 37473 26333 37507 26367
rect 37657 26333 37691 26367
rect 37749 26333 37783 26367
rect 38301 26333 38335 26367
rect 39037 26333 39071 26367
rect 5181 26265 5215 26299
rect 10241 26265 10275 26299
rect 10609 26265 10643 26299
rect 16129 26265 16163 26299
rect 17760 26265 17794 26299
rect 20453 26265 20487 26299
rect 20570 26265 20604 26299
rect 24777 26265 24811 26299
rect 31585 26265 31619 26299
rect 33793 26265 33827 26299
rect 35081 26265 35115 26299
rect 35633 26265 35667 26299
rect 35833 26265 35867 26299
rect 36277 26265 36311 26299
rect 4445 26197 4479 26231
rect 6009 26197 6043 26231
rect 12173 26197 12207 26231
rect 15669 26197 15703 26231
rect 17601 26197 17635 26231
rect 19441 26197 19475 26231
rect 20361 26197 20395 26231
rect 20729 26197 20763 26231
rect 21281 26197 21315 26231
rect 21465 26197 21499 26231
rect 22109 26197 22143 26231
rect 22293 26197 22327 26231
rect 23581 26197 23615 26231
rect 26249 26197 26283 26231
rect 37933 26197 37967 26231
rect 38117 26197 38151 26231
rect 1501 25993 1535 26027
rect 4445 25993 4479 26027
rect 4629 25993 4663 26027
rect 7113 25993 7147 26027
rect 8309 25993 8343 26027
rect 8953 25993 8987 26027
rect 9413 25993 9447 26027
rect 11529 25993 11563 26027
rect 11989 25993 12023 26027
rect 14749 25993 14783 26027
rect 14933 25993 14967 26027
rect 16037 25993 16071 26027
rect 22293 25993 22327 26027
rect 23581 25993 23615 26027
rect 24961 25993 24995 26027
rect 29377 25993 29411 26027
rect 32413 25993 32447 26027
rect 32505 25993 32539 26027
rect 39037 25993 39071 26027
rect 39865 25993 39899 26027
rect 40509 25993 40543 26027
rect 42073 25993 42107 26027
rect 8033 25925 8067 25959
rect 8677 25925 8711 25959
rect 10526 25925 10560 25959
rect 11897 25925 11931 25959
rect 21465 25925 21499 25959
rect 21649 25925 21683 25959
rect 22385 25925 22419 25959
rect 22661 25925 22695 25959
rect 37565 25925 37599 25959
rect 39313 25925 39347 25959
rect 39497 25925 39531 25959
rect 40789 25925 40823 25959
rect 1685 25857 1719 25891
rect 2697 25857 2731 25891
rect 3157 25857 3191 25891
rect 3709 25857 3743 25891
rect 3893 25857 3927 25891
rect 3986 25857 4020 25891
rect 4353 25857 4387 25891
rect 4537 25857 4571 25891
rect 5089 25857 5123 25891
rect 5825 25857 5859 25891
rect 5917 25857 5951 25891
rect 6101 25857 6135 25891
rect 7297 25857 7331 25891
rect 7389 25857 7423 25891
rect 7665 25857 7699 25891
rect 7757 25857 7791 25891
rect 7941 25857 7975 25891
rect 8125 25857 8159 25891
rect 8401 25857 8435 25891
rect 8585 25857 8619 25891
rect 8769 25857 8803 25891
rect 10793 25857 10827 25891
rect 12541 25857 12575 25891
rect 12725 25857 12759 25891
rect 14381 25857 14415 25891
rect 14535 25857 14569 25891
rect 14841 25857 14875 25891
rect 15025 25857 15059 25891
rect 15117 25857 15151 25891
rect 15209 25857 15243 25891
rect 15393 25857 15427 25891
rect 15485 25857 15519 25891
rect 16129 25857 16163 25891
rect 16957 25857 16991 25891
rect 19993 25857 20027 25891
rect 20085 25857 20119 25891
rect 20361 25857 20395 25891
rect 21097 25857 21131 25891
rect 21281 25857 21315 25891
rect 21373 25857 21407 25891
rect 22017 25857 22051 25891
rect 22470 25857 22504 25891
rect 22559 25857 22593 25891
rect 22845 25857 22879 25891
rect 23305 25857 23339 25891
rect 23489 25857 23523 25891
rect 23857 25857 23891 25891
rect 25145 25857 25179 25891
rect 25421 25857 25455 25891
rect 40049 25857 40083 25891
rect 40141 25857 40175 25891
rect 40233 25857 40267 25891
rect 40417 25857 40451 25891
rect 40693 25857 40727 25891
rect 40877 25857 40911 25891
rect 41061 25857 41095 25891
rect 41889 25857 41923 25891
rect 3525 25789 3559 25823
rect 4261 25789 4295 25823
rect 4997 25789 5031 25823
rect 5273 25789 5307 25823
rect 5457 25789 5491 25823
rect 5549 25789 5583 25823
rect 12173 25789 12207 25823
rect 16681 25789 16715 25823
rect 20269 25789 20303 25823
rect 23949 25789 23983 25823
rect 27629 25789 27663 25823
rect 27905 25789 27939 25823
rect 32229 25789 32263 25823
rect 37289 25789 37323 25823
rect 5641 25721 5675 25755
rect 7573 25721 7607 25755
rect 16773 25721 16807 25755
rect 16865 25721 16899 25755
rect 21281 25721 21315 25755
rect 24225 25721 24259 25755
rect 5733 25653 5767 25687
rect 6009 25653 6043 25687
rect 12541 25653 12575 25687
rect 15669 25653 15703 25687
rect 21557 25653 21591 25687
rect 23029 25653 23063 25687
rect 23765 25653 23799 25687
rect 23857 25653 23891 25687
rect 25329 25653 25363 25687
rect 32873 25653 32907 25687
rect 39129 25653 39163 25687
rect 14749 25449 14783 25483
rect 15393 25449 15427 25483
rect 17325 25449 17359 25483
rect 18153 25449 18187 25483
rect 24961 25449 24995 25483
rect 28181 25449 28215 25483
rect 40325 25449 40359 25483
rect 41889 25449 41923 25483
rect 30205 25381 30239 25415
rect 30573 25381 30607 25415
rect 2881 25313 2915 25347
rect 3157 25313 3191 25347
rect 15117 25313 15151 25347
rect 15853 25313 15887 25347
rect 28825 25313 28859 25347
rect 34529 25313 34563 25347
rect 4997 25245 5031 25279
rect 7665 25245 7699 25279
rect 7849 25245 7883 25279
rect 13461 25245 13495 25279
rect 15025 25245 15059 25279
rect 15485 25245 15519 25279
rect 15577 25245 15611 25279
rect 18061 25245 18095 25279
rect 18245 25245 18279 25279
rect 21281 25245 21315 25279
rect 21649 25245 21683 25279
rect 21741 25245 21775 25279
rect 22293 25245 22327 25279
rect 23213 25245 23247 25279
rect 23305 25245 23339 25279
rect 23673 25245 23707 25279
rect 25145 25245 25179 25279
rect 25237 25245 25271 25279
rect 25513 25245 25547 25279
rect 25605 25245 25639 25279
rect 25789 25245 25823 25279
rect 26985 25245 27019 25279
rect 27169 25245 27203 25279
rect 29653 25245 29687 25279
rect 30297 25245 30331 25279
rect 30389 25245 30423 25279
rect 30849 25245 30883 25279
rect 31125 25245 31159 25279
rect 35449 25245 35483 25279
rect 35725 25245 35759 25279
rect 36001 25245 36035 25279
rect 36369 25245 36403 25279
rect 36645 25245 36679 25279
rect 37013 25245 37047 25279
rect 41337 25245 41371 25279
rect 14381 25177 14415 25211
rect 14565 25177 14599 25211
rect 17509 25177 17543 25211
rect 17877 25177 17911 25211
rect 21419 25177 21453 25211
rect 21557 25177 21591 25211
rect 21925 25177 21959 25211
rect 23397 25177 23431 25211
rect 23535 25177 23569 25211
rect 25329 25177 25363 25211
rect 25973 25177 26007 25211
rect 30021 25177 30055 25211
rect 30573 25177 30607 25211
rect 32505 25177 32539 25211
rect 34253 25177 34287 25211
rect 35541 25177 35575 25211
rect 35909 25177 35943 25211
rect 36185 25177 36219 25211
rect 40509 25177 40543 25211
rect 40693 25177 40727 25211
rect 41797 25177 41831 25211
rect 1409 25109 1443 25143
rect 5181 25109 5215 25143
rect 7849 25109 7883 25143
rect 13369 25109 13403 25143
rect 14841 25109 14875 25143
rect 18429 25109 18463 25143
rect 22109 25109 22143 25143
rect 23029 25109 23063 25143
rect 27077 25109 27111 25143
rect 28549 25109 28583 25143
rect 28641 25109 28675 25143
rect 29745 25109 29779 25143
rect 30665 25109 30699 25143
rect 31033 25109 31067 25143
rect 35449 25109 35483 25143
rect 36553 25109 36587 25143
rect 40877 25109 40911 25143
rect 41521 25109 41555 25143
rect 7205 24905 7239 24939
rect 7573 24905 7607 24939
rect 8217 24905 8251 24939
rect 8861 24905 8895 24939
rect 12817 24905 12851 24939
rect 20177 24905 20211 24939
rect 22201 24905 22235 24939
rect 25053 24905 25087 24939
rect 28733 24905 28767 24939
rect 31861 24905 31895 24939
rect 33885 24905 33919 24939
rect 40693 24905 40727 24939
rect 7113 24837 7147 24871
rect 13461 24837 13495 24871
rect 19809 24837 19843 24871
rect 25697 24837 25731 24871
rect 25897 24837 25931 24871
rect 26525 24837 26559 24871
rect 27445 24837 27479 24871
rect 29653 24837 29687 24871
rect 35817 24837 35851 24871
rect 36737 24837 36771 24871
rect 37381 24837 37415 24871
rect 39129 24837 39163 24871
rect 41061 24837 41095 24871
rect 42073 24837 42107 24871
rect 1409 24769 1443 24803
rect 3709 24769 3743 24803
rect 3801 24769 3835 24803
rect 3893 24769 3927 24803
rect 4445 24769 4479 24803
rect 4537 24769 4571 24803
rect 4629 24769 4663 24803
rect 4813 24769 4847 24803
rect 4905 24769 4939 24803
rect 5089 24769 5123 24803
rect 5273 24769 5307 24803
rect 6561 24769 6595 24803
rect 6745 24769 6779 24803
rect 6837 24769 6871 24803
rect 7205 24769 7239 24803
rect 7757 24769 7791 24803
rect 7849 24769 7883 24803
rect 7941 24769 7975 24803
rect 8493 24769 8527 24803
rect 8585 24769 8619 24803
rect 9045 24769 9079 24803
rect 9229 24769 9263 24803
rect 9321 24769 9355 24803
rect 9689 24769 9723 24803
rect 9873 24769 9907 24803
rect 9965 24769 9999 24803
rect 10057 24769 10091 24803
rect 12725 24769 12759 24803
rect 13737 24769 13771 24803
rect 14381 24769 14415 24803
rect 14657 24769 14691 24803
rect 14749 24769 14783 24803
rect 14933 24769 14967 24803
rect 15669 24769 15703 24803
rect 15853 24769 15887 24803
rect 15945 24769 15979 24803
rect 17141 24769 17175 24803
rect 19165 24769 19199 24803
rect 19349 24769 19383 24803
rect 19625 24769 19659 24803
rect 19901 24769 19935 24803
rect 20085 24769 20119 24803
rect 20361 24769 20395 24803
rect 22293 24769 22327 24803
rect 22937 24769 22971 24803
rect 24777 24769 24811 24803
rect 25329 24769 25363 24803
rect 26341 24769 26375 24803
rect 26433 24769 26467 24803
rect 27169 24769 27203 24803
rect 27262 24769 27296 24803
rect 27537 24769 27571 24803
rect 27675 24769 27709 24803
rect 27997 24769 28031 24803
rect 28457 24769 28491 24803
rect 28641 24769 28675 24803
rect 28917 24769 28951 24803
rect 29009 24769 29043 24803
rect 29101 24769 29135 24803
rect 29239 24769 29273 24803
rect 29469 24769 29503 24803
rect 29837 24769 29871 24803
rect 32321 24769 32355 24803
rect 32689 24769 32723 24803
rect 32782 24769 32816 24803
rect 32965 24769 32999 24803
rect 33057 24769 33091 24803
rect 33154 24769 33188 24803
rect 33701 24769 33735 24803
rect 35081 24769 35115 24803
rect 35265 24769 35299 24803
rect 35357 24769 35391 24803
rect 35449 24769 35483 24803
rect 35607 24769 35641 24803
rect 35725 24769 35759 24803
rect 35909 24769 35943 24803
rect 36093 24769 36127 24803
rect 36645 24769 36679 24803
rect 38209 24769 38243 24803
rect 40877 24769 40911 24803
rect 40969 24769 41003 24803
rect 41245 24769 41279 24803
rect 41337 24769 41371 24803
rect 4077 24701 4111 24735
rect 4997 24701 5031 24735
rect 6101 24701 6135 24735
rect 6653 24701 6687 24735
rect 7113 24701 7147 24735
rect 7481 24701 7515 24735
rect 8033 24701 8067 24735
rect 8401 24701 8435 24735
rect 8677 24701 8711 24735
rect 11161 24701 11195 24735
rect 12081 24701 12115 24735
rect 14565 24701 14599 24735
rect 18153 24701 18187 24735
rect 19441 24701 19475 24735
rect 22477 24701 22511 24735
rect 25053 24701 25087 24735
rect 25513 24701 25547 24735
rect 26709 24701 26743 24735
rect 28549 24701 28583 24735
rect 29377 24701 29411 24735
rect 30113 24701 30147 24735
rect 30389 24701 30423 24735
rect 32137 24701 32171 24735
rect 33425 24701 33459 24735
rect 36461 24701 36495 24735
rect 38853 24701 38887 24735
rect 40601 24701 40635 24735
rect 1593 24633 1627 24667
rect 4169 24633 4203 24667
rect 7297 24633 7331 24667
rect 10517 24633 10551 24667
rect 12357 24633 12391 24667
rect 18429 24633 18463 24667
rect 19349 24633 19383 24667
rect 22753 24633 22787 24667
rect 24869 24633 24903 24667
rect 25145 24633 25179 24667
rect 26157 24633 26191 24667
rect 28181 24633 28215 24667
rect 33333 24633 33367 24667
rect 41797 24633 41831 24667
rect 6929 24565 6963 24599
rect 10241 24565 10275 24599
rect 12541 24565 12575 24599
rect 13001 24565 13035 24599
rect 13093 24565 13127 24599
rect 13185 24565 13219 24599
rect 14013 24565 14047 24599
rect 14197 24565 14231 24599
rect 17049 24565 17083 24599
rect 18613 24565 18647 24599
rect 21833 24565 21867 24599
rect 25881 24565 25915 24599
rect 26065 24565 26099 24599
rect 27813 24565 27847 24599
rect 33517 24565 33551 24599
rect 34897 24565 34931 24599
rect 37105 24565 37139 24599
rect 41521 24565 41555 24599
rect 4905 24361 4939 24395
rect 5089 24361 5123 24395
rect 6745 24361 6779 24395
rect 7849 24361 7883 24395
rect 8033 24361 8067 24395
rect 9229 24361 9263 24395
rect 11345 24361 11379 24395
rect 13185 24361 13219 24395
rect 15025 24361 15059 24395
rect 20361 24361 20395 24395
rect 25421 24361 25455 24395
rect 26341 24361 26375 24395
rect 26617 24361 26651 24395
rect 29929 24361 29963 24395
rect 30297 24361 30331 24395
rect 30757 24361 30791 24395
rect 30941 24361 30975 24395
rect 32965 24361 32999 24395
rect 42165 24361 42199 24395
rect 6285 24293 6319 24327
rect 7021 24293 7055 24327
rect 23949 24293 23983 24327
rect 25605 24293 25639 24327
rect 30113 24293 30147 24327
rect 1593 24225 1627 24259
rect 7573 24225 7607 24259
rect 13277 24225 13311 24259
rect 14657 24225 14691 24259
rect 16773 24225 16807 24259
rect 20177 24225 20211 24259
rect 21833 24225 21867 24259
rect 22109 24225 22143 24259
rect 22201 24225 22235 24259
rect 25789 24225 25823 24259
rect 26893 24225 26927 24259
rect 32505 24225 32539 24259
rect 35909 24225 35943 24259
rect 36277 24225 36311 24259
rect 37013 24225 37047 24259
rect 37289 24225 37323 24259
rect 39037 24225 39071 24259
rect 40693 24225 40727 24259
rect 3617 24157 3651 24191
rect 4353 24157 4387 24191
rect 4537 24157 4571 24191
rect 5181 24157 5215 24191
rect 5365 24157 5399 24191
rect 6101 24157 6135 24191
rect 6561 24157 6595 24191
rect 6653 24157 6687 24191
rect 6837 24157 6871 24191
rect 6929 24157 6963 24191
rect 7113 24157 7147 24191
rect 7205 24157 7239 24191
rect 8401 24157 8435 24191
rect 8493 24157 8527 24191
rect 9045 24157 9079 24191
rect 9229 24157 9263 24191
rect 9321 24157 9355 24191
rect 9505 24157 9539 24191
rect 9597 24157 9631 24191
rect 9689 24157 9723 24191
rect 9965 24157 9999 24191
rect 11805 24157 11839 24191
rect 14565 24157 14599 24191
rect 14933 24157 14967 24191
rect 15209 24157 15243 24191
rect 15393 24157 15427 24191
rect 16865 24157 16899 24191
rect 17233 24157 17267 24191
rect 18061 24157 18095 24191
rect 18705 24157 18739 24191
rect 18981 24157 19015 24191
rect 19257 24157 19291 24191
rect 19441 24157 19475 24191
rect 19717 24157 19751 24191
rect 24593 24157 24627 24191
rect 24869 24157 24903 24191
rect 24961 24157 24995 24191
rect 25145 24157 25179 24191
rect 25237 24157 25271 24191
rect 25513 24157 25547 24191
rect 25881 24157 25915 24191
rect 26249 24157 26283 24191
rect 26341 24157 26375 24191
rect 26525 24157 26559 24191
rect 26617 24157 26651 24191
rect 26801 24157 26835 24191
rect 30481 24157 30515 24191
rect 30573 24157 30607 24191
rect 30849 24157 30883 24191
rect 32597 24157 32631 24191
rect 34713 24157 34747 24191
rect 35541 24157 35575 24191
rect 35633 24157 35667 24191
rect 40049 24157 40083 24191
rect 40417 24157 40451 24191
rect 1869 24089 1903 24123
rect 5273 24089 5307 24123
rect 6285 24089 6319 24123
rect 7389 24089 7423 24123
rect 7665 24089 7699 24123
rect 7865 24089 7899 24123
rect 8677 24089 8711 24123
rect 10210 24089 10244 24123
rect 12072 24089 12106 24123
rect 13921 24089 13955 24123
rect 14473 24089 14507 24123
rect 17141 24089 17175 24123
rect 18245 24089 18279 24123
rect 19809 24089 19843 24123
rect 19901 24089 19935 24123
rect 20039 24089 20073 24123
rect 22477 24089 22511 24123
rect 24685 24089 24719 24123
rect 26157 24089 26191 24123
rect 27169 24089 27203 24123
rect 29745 24089 29779 24123
rect 29945 24089 29979 24123
rect 31125 24089 31159 24123
rect 31309 24089 31343 24123
rect 34897 24089 34931 24123
rect 35081 24089 35115 24123
rect 35265 24089 35299 24123
rect 36001 24089 36035 24123
rect 39313 24089 39347 24123
rect 39497 24089 39531 24123
rect 3801 24021 3835 24055
rect 4905 24021 4939 24055
rect 6469 24021 6503 24055
rect 8401 24021 8435 24055
rect 9873 24021 9907 24055
rect 14105 24021 14139 24055
rect 15301 24021 15335 24055
rect 16589 24021 16623 24055
rect 16957 24021 16991 24055
rect 18429 24021 18463 24055
rect 18521 24021 18555 24055
rect 18889 24021 18923 24055
rect 19349 24021 19383 24055
rect 19533 24021 19567 24055
rect 24770 24021 24804 24055
rect 28641 24021 28675 24055
rect 34989 24021 35023 24055
rect 35357 24021 35391 24055
rect 36461 24021 36495 24055
rect 36553 24021 36587 24055
rect 36921 24021 36955 24055
rect 39681 24021 39715 24055
rect 40233 24021 40267 24055
rect 2329 23817 2363 23851
rect 3985 23817 4019 23851
rect 8953 23817 8987 23851
rect 13369 23817 13403 23851
rect 19901 23817 19935 23851
rect 20361 23817 20395 23851
rect 21925 23817 21959 23851
rect 22661 23817 22695 23851
rect 23121 23817 23155 23851
rect 26985 23817 27019 23851
rect 27537 23817 27571 23851
rect 30297 23817 30331 23851
rect 35005 23817 35039 23851
rect 2145 23749 2179 23783
rect 4629 23749 4663 23783
rect 9505 23749 9539 23783
rect 10232 23749 10266 23783
rect 17785 23749 17819 23783
rect 18613 23749 18647 23783
rect 24593 23749 24627 23783
rect 27905 23749 27939 23783
rect 28365 23749 28399 23783
rect 31309 23749 31343 23783
rect 34805 23749 34839 23783
rect 37565 23749 37599 23783
rect 39773 23749 39807 23783
rect 41705 23749 41739 23783
rect 1409 23681 1443 23715
rect 2421 23681 2455 23715
rect 3709 23681 3743 23715
rect 3801 23681 3835 23715
rect 4077 23681 4111 23715
rect 6653 23681 6687 23715
rect 7205 23681 7239 23715
rect 7389 23681 7423 23715
rect 7481 23681 7515 23715
rect 7573 23681 7607 23715
rect 8861 23681 8895 23715
rect 9321 23681 9355 23715
rect 9597 23681 9631 23715
rect 9689 23681 9723 23715
rect 9965 23681 9999 23715
rect 11989 23681 12023 23715
rect 12256 23681 12290 23715
rect 13829 23681 13863 23715
rect 14841 23681 14875 23715
rect 16221 23681 16255 23715
rect 16405 23681 16439 23715
rect 16497 23681 16531 23715
rect 17049 23681 17083 23715
rect 17647 23681 17681 23715
rect 17877 23681 17911 23715
rect 18005 23681 18039 23715
rect 18153 23681 18187 23715
rect 18429 23681 18463 23715
rect 18521 23681 18555 23715
rect 18797 23681 18831 23715
rect 20269 23681 20303 23715
rect 20545 23681 20579 23715
rect 20637 23681 20671 23715
rect 22109 23681 22143 23715
rect 23029 23681 23063 23715
rect 24317 23681 24351 23715
rect 27169 23681 27203 23715
rect 30205 23681 30239 23715
rect 31125 23681 31159 23715
rect 31677 23681 31711 23715
rect 35357 23681 35391 23715
rect 35449 23681 35483 23715
rect 37289 23681 37323 23715
rect 39497 23681 39531 23715
rect 41521 23681 41555 23715
rect 41613 23681 41647 23715
rect 41889 23681 41923 23715
rect 3617 23613 3651 23647
rect 4353 23613 4387 23647
rect 6101 23613 6135 23647
rect 13921 23613 13955 23647
rect 14013 23613 14047 23647
rect 14289 23613 14323 23647
rect 17141 23613 17175 23647
rect 17417 23613 17451 23647
rect 20177 23613 20211 23647
rect 20361 23613 20395 23647
rect 23305 23613 23339 23647
rect 27445 23613 27479 23647
rect 27997 23613 28031 23647
rect 28089 23613 28123 23647
rect 28917 23613 28951 23647
rect 30941 23613 30975 23647
rect 31401 23613 31435 23647
rect 35633 23613 35667 23647
rect 39037 23613 39071 23647
rect 41245 23613 41279 23647
rect 2145 23545 2179 23579
rect 13461 23545 13495 23579
rect 17509 23545 17543 23579
rect 26065 23545 26099 23579
rect 27353 23545 27387 23579
rect 31585 23545 31619 23579
rect 35173 23545 35207 23579
rect 1593 23477 1627 23511
rect 4261 23477 4295 23511
rect 6469 23477 6503 23511
rect 7849 23477 7883 23511
rect 9873 23477 9907 23511
rect 11345 23477 11379 23511
rect 16037 23477 16071 23511
rect 18245 23477 18279 23511
rect 20177 23477 20211 23511
rect 31493 23477 31527 23511
rect 34989 23477 35023 23511
rect 35541 23477 35575 23511
rect 41337 23477 41371 23511
rect 1409 23273 1443 23307
rect 5457 23273 5491 23307
rect 5641 23273 5675 23307
rect 21925 23273 21959 23307
rect 39129 23273 39163 23307
rect 7389 23205 7423 23239
rect 11529 23205 11563 23239
rect 14381 23205 14415 23239
rect 14841 23205 14875 23239
rect 17417 23205 17451 23239
rect 13737 23137 13771 23171
rect 14197 23137 14231 23171
rect 15209 23137 15243 23171
rect 19717 23137 19751 23171
rect 19901 23137 19935 23171
rect 30941 23137 30975 23171
rect 31401 23137 31435 23171
rect 31769 23137 31803 23171
rect 31861 23137 31895 23171
rect 34529 23137 34563 23171
rect 35357 23137 35391 23171
rect 35725 23137 35759 23171
rect 36093 23137 36127 23171
rect 36829 23137 36863 23171
rect 39957 23137 39991 23171
rect 40693 23137 40727 23171
rect 3157 23069 3191 23103
rect 7113 23069 7147 23103
rect 7297 23069 7331 23103
rect 7481 23069 7515 23103
rect 7573 23069 7607 23103
rect 10149 23069 10183 23103
rect 10405 23069 10439 23103
rect 13461 23069 13495 23103
rect 13645 23069 13679 23103
rect 13829 23069 13863 23103
rect 14473 23069 14507 23103
rect 14657 23069 14691 23103
rect 14841 23069 14875 23103
rect 15117 23069 15151 23103
rect 15301 23069 15335 23103
rect 15393 23069 15427 23103
rect 15669 23069 15703 23103
rect 17693 23069 17727 23103
rect 20637 23069 20671 23103
rect 22661 23069 22695 23103
rect 25605 23069 25639 23103
rect 25881 23069 25915 23103
rect 25973 23069 26007 23103
rect 29009 23069 29043 23103
rect 31493 23069 31527 23103
rect 33517 23069 33551 23103
rect 34253 23069 34287 23103
rect 34345 23069 34379 23103
rect 35817 23069 35851 23103
rect 36461 23069 36495 23103
rect 36553 23069 36587 23103
rect 38669 23069 38703 23103
rect 39313 23069 39347 23103
rect 39405 23069 39439 23103
rect 39497 23069 39531 23103
rect 39681 23069 39715 23103
rect 40417 23069 40451 23103
rect 2881 23001 2915 23035
rect 5273 23001 5307 23035
rect 15945 23001 15979 23035
rect 19625 23001 19659 23035
rect 25789 23001 25823 23035
rect 28764 23001 28798 23035
rect 30757 23001 30791 23035
rect 33272 23001 33306 23035
rect 34529 23001 34563 23035
rect 36185 23001 36219 23035
rect 36921 23001 36955 23035
rect 40141 23001 40175 23035
rect 40325 23001 40359 23035
rect 5483 22933 5517 22967
rect 7757 22933 7791 22967
rect 12909 22933 12943 22967
rect 14197 22933 14231 22967
rect 15577 22933 15611 22967
rect 19257 22933 19291 22967
rect 23213 22933 23247 22967
rect 26157 22933 26191 22967
rect 27629 22933 27663 22967
rect 30389 22933 30423 22967
rect 30849 22933 30883 22967
rect 31217 22933 31251 22967
rect 32137 22933 32171 22967
rect 34713 22933 34747 22967
rect 35081 22933 35115 22967
rect 35173 22933 35207 22967
rect 35541 22933 35575 22967
rect 36277 22933 36311 22967
rect 38025 22933 38059 22967
rect 42165 22933 42199 22967
rect 7941 22729 7975 22763
rect 10609 22729 10643 22763
rect 12633 22729 12667 22763
rect 13829 22729 13863 22763
rect 16037 22729 16071 22763
rect 20269 22729 20303 22763
rect 24225 22729 24259 22763
rect 26157 22729 26191 22763
rect 31769 22729 31803 22763
rect 33425 22729 33459 22763
rect 35265 22729 35299 22763
rect 36461 22729 36495 22763
rect 36553 22729 36587 22763
rect 38669 22729 38703 22763
rect 40325 22729 40359 22763
rect 41153 22729 41187 22763
rect 8033 22661 8067 22695
rect 11713 22661 11747 22695
rect 13921 22661 13955 22695
rect 14565 22661 14599 22695
rect 17601 22661 17635 22695
rect 18797 22661 18831 22695
rect 20729 22661 20763 22695
rect 24685 22661 24719 22695
rect 30297 22661 30331 22695
rect 34897 22661 34931 22695
rect 7757 22593 7791 22627
rect 8125 22593 8159 22627
rect 8381 22593 8415 22627
rect 10241 22593 10275 22627
rect 14289 22593 14323 22627
rect 16221 22593 16255 22627
rect 17969 22593 18003 22627
rect 18153 22593 18187 22627
rect 18245 22593 18279 22627
rect 20637 22593 20671 22627
rect 20821 22593 20855 22627
rect 21005 22593 21039 22627
rect 21097 22593 21131 22627
rect 21373 22593 21407 22627
rect 21465 22593 21499 22627
rect 22836 22593 22870 22627
rect 24593 22593 24627 22627
rect 25053 22593 25087 22627
rect 25789 22593 25823 22627
rect 27169 22593 27203 22627
rect 27813 22593 27847 22627
rect 30021 22593 30055 22627
rect 32689 22593 32723 22627
rect 35173 22593 35207 22627
rect 35449 22593 35483 22627
rect 35633 22593 35667 22627
rect 38577 22593 38611 22627
rect 39773 22593 39807 22627
rect 40233 22593 40267 22627
rect 41061 22593 41095 22627
rect 2881 22525 2915 22559
rect 3157 22525 3191 22559
rect 3433 22525 3467 22559
rect 3801 22525 3835 22559
rect 7665 22525 7699 22559
rect 11253 22525 11287 22559
rect 12173 22525 12207 22559
rect 12725 22525 12759 22559
rect 12909 22525 12943 22559
rect 14013 22525 14047 22559
rect 16773 22525 16807 22559
rect 18521 22525 18555 22559
rect 21833 22525 21867 22559
rect 22569 22525 22603 22559
rect 24777 22525 24811 22559
rect 25605 22525 25639 22559
rect 26801 22525 26835 22559
rect 33333 22525 33367 22559
rect 36277 22525 36311 22559
rect 38761 22525 38795 22559
rect 40417 22525 40451 22559
rect 41245 22525 41279 22559
rect 42073 22525 42107 22559
rect 7573 22457 7607 22491
rect 9597 22457 9631 22491
rect 11989 22457 12023 22491
rect 22477 22457 22511 22491
rect 23949 22457 23983 22491
rect 39589 22457 39623 22491
rect 1409 22389 1443 22423
rect 5181 22389 5215 22423
rect 9505 22389 9539 22423
rect 12265 22389 12299 22423
rect 13461 22389 13495 22423
rect 16405 22389 16439 22423
rect 17785 22389 17819 22423
rect 20453 22389 20487 22423
rect 21189 22389 21223 22423
rect 21649 22389 21683 22423
rect 25973 22389 26007 22423
rect 27721 22389 27755 22423
rect 36921 22389 36955 22423
rect 38209 22389 38243 22423
rect 39865 22389 39899 22423
rect 40693 22389 40727 22423
rect 41521 22389 41555 22423
rect 7757 22185 7791 22219
rect 14749 22185 14783 22219
rect 17496 22185 17530 22219
rect 18981 22185 19015 22219
rect 23121 22185 23155 22219
rect 34713 22185 34747 22219
rect 36540 22185 36574 22219
rect 41245 22185 41279 22219
rect 16129 22117 16163 22151
rect 3893 22049 3927 22083
rect 7389 22049 7423 22083
rect 7849 22049 7883 22083
rect 9137 22049 9171 22083
rect 15761 22049 15795 22083
rect 17233 22049 17267 22083
rect 23581 22049 23615 22083
rect 23765 22049 23799 22083
rect 24961 22049 24995 22083
rect 30205 22049 30239 22083
rect 36277 22049 36311 22083
rect 38025 22049 38059 22083
rect 41981 22049 42015 22083
rect 1409 21981 1443 22015
rect 4261 21981 4295 22015
rect 6837 21981 6871 22015
rect 7113 21981 7147 22015
rect 7297 21981 7331 22015
rect 7481 21981 7515 22015
rect 7757 21981 7791 22015
rect 8493 21981 8527 22015
rect 12541 21981 12575 22015
rect 12808 21981 12842 22015
rect 14105 21981 14139 22015
rect 15209 21981 15243 22015
rect 15301 21981 15335 22015
rect 15577 21981 15611 22015
rect 15669 21981 15703 22015
rect 15945 21981 15979 22015
rect 16221 21981 16255 22015
rect 19993 21981 20027 22015
rect 21465 21981 21499 22015
rect 21732 21981 21766 22015
rect 23949 21981 23983 22015
rect 25145 21981 25179 22015
rect 26617 21981 26651 22015
rect 30941 21981 30975 22015
rect 31309 21981 31343 22015
rect 31401 21981 31435 22015
rect 31677 21981 31711 22015
rect 32137 21981 32171 22015
rect 34161 21981 34195 22015
rect 34897 21981 34931 22015
rect 35265 21981 35299 22015
rect 39037 21981 39071 22015
rect 39865 21981 39899 22015
rect 41337 21981 41371 22015
rect 6745 21913 6779 21947
rect 9413 21913 9447 21947
rect 11161 21913 11195 21947
rect 15393 21913 15427 21947
rect 20260 21913 20294 21947
rect 24409 21913 24443 21947
rect 25412 21913 25446 21947
rect 26862 21913 26896 21947
rect 28273 21913 28307 21947
rect 29009 21913 29043 21947
rect 30021 21913 30055 21947
rect 31493 21913 31527 21947
rect 32404 21913 32438 21947
rect 33609 21913 33643 21947
rect 34989 21913 35023 21947
rect 35081 21913 35115 21947
rect 38209 21913 38243 21947
rect 40132 21913 40166 21947
rect 1593 21845 1627 21879
rect 5687 21845 5721 21879
rect 6929 21845 6963 21879
rect 7573 21845 7607 21879
rect 13921 21845 13955 21879
rect 15025 21845 15059 21879
rect 16313 21845 16347 21879
rect 21373 21845 21407 21879
rect 22845 21845 22879 21879
rect 23489 21845 23523 21879
rect 24133 21845 24167 21879
rect 26525 21845 26559 21879
rect 27997 21845 28031 21879
rect 29561 21845 29595 21879
rect 29929 21845 29963 21879
rect 30389 21845 30423 21879
rect 31125 21845 31159 21879
rect 33517 21845 33551 21879
rect 4445 21641 4479 21675
rect 8309 21641 8343 21675
rect 9597 21641 9631 21675
rect 13001 21641 13035 21675
rect 15577 21641 15611 21675
rect 17049 21641 17083 21675
rect 22293 21641 22327 21675
rect 24869 21641 24903 21675
rect 25605 21641 25639 21675
rect 28365 21641 28399 21675
rect 29837 21641 29871 21675
rect 32413 21641 32447 21675
rect 41337 21641 41371 21675
rect 5089 21573 5123 21607
rect 9229 21573 9263 21607
rect 9321 21573 9355 21607
rect 11888 21573 11922 21607
rect 16773 21573 16807 21607
rect 17325 21573 17359 21607
rect 23756 21573 23790 21607
rect 25329 21573 25363 21607
rect 28724 21573 28758 21607
rect 32781 21573 32815 21607
rect 34161 21573 34195 21607
rect 34253 21573 34287 21607
rect 34713 21573 34747 21607
rect 34805 21573 34839 21607
rect 4629 21505 4663 21539
rect 4721 21505 4755 21539
rect 4905 21505 4939 21539
rect 4997 21505 5031 21539
rect 5273 21505 5307 21539
rect 5365 21505 5399 21539
rect 5549 21505 5583 21539
rect 5641 21505 5675 21539
rect 5917 21505 5951 21539
rect 9045 21505 9079 21539
rect 9413 21505 9447 21539
rect 11621 21505 11655 21539
rect 15301 21505 15335 21539
rect 18889 21505 18923 21539
rect 19156 21505 19190 21539
rect 22201 21505 22235 21539
rect 25053 21505 25087 21539
rect 25237 21505 25271 21539
rect 25421 21505 25455 21539
rect 26985 21505 27019 21539
rect 27252 21505 27286 21539
rect 32597 21505 32631 21539
rect 32689 21505 32723 21539
rect 32965 21505 32999 21539
rect 34069 21505 34103 21539
rect 34437 21505 34471 21539
rect 34529 21505 34563 21539
rect 34897 21505 34931 21539
rect 37933 21505 37967 21539
rect 39957 21505 39991 21539
rect 40224 21505 40258 21539
rect 3157 21437 3191 21471
rect 6193 21437 6227 21471
rect 6377 21437 6411 21471
rect 6745 21437 6779 21471
rect 8861 21437 8895 21471
rect 16129 21437 16163 21471
rect 17509 21437 17543 21471
rect 21005 21437 21039 21471
rect 22385 21437 22419 21471
rect 22661 21437 22695 21471
rect 23213 21437 23247 21471
rect 23489 21437 23523 21471
rect 25881 21437 25915 21471
rect 26525 21437 26559 21471
rect 28457 21437 28491 21471
rect 30665 21437 30699 21471
rect 31861 21437 31895 21471
rect 33241 21437 33275 21471
rect 35633 21437 35667 21471
rect 41981 21437 42015 21471
rect 20269 21369 20303 21403
rect 2605 21301 2639 21335
rect 6009 21301 6043 21335
rect 6101 21301 6135 21335
rect 8171 21301 8205 21335
rect 14749 21301 14783 21335
rect 20361 21301 20395 21335
rect 21833 21301 21867 21335
rect 30113 21301 30147 21335
rect 31217 21301 31251 21335
rect 33793 21301 33827 21335
rect 33885 21301 33919 21335
rect 35081 21301 35115 21335
rect 36277 21301 36311 21335
rect 41429 21301 41463 21335
rect 5181 21097 5215 21131
rect 6101 21097 6135 21131
rect 8125 21097 8159 21131
rect 15485 21097 15519 21131
rect 17509 21097 17543 21131
rect 19257 21097 19291 21131
rect 22293 21097 22327 21131
rect 29009 21097 29043 21131
rect 38669 21097 38703 21131
rect 3157 21029 3191 21063
rect 4537 21029 4571 21063
rect 10885 21029 10919 21063
rect 18337 21029 18371 21063
rect 27629 21029 27663 21063
rect 6377 20961 6411 20995
rect 11529 20961 11563 20995
rect 11805 20961 11839 20995
rect 16037 20961 16071 20995
rect 16221 20961 16255 20995
rect 18429 20961 18463 20995
rect 24869 20961 24903 20995
rect 24961 20961 24995 20995
rect 28273 20961 28307 20995
rect 30021 20961 30055 20995
rect 30205 20961 30239 20995
rect 30481 20961 30515 20995
rect 39221 20961 39255 20995
rect 39405 20961 39439 20995
rect 40417 20961 40451 20995
rect 1777 20893 1811 20927
rect 2044 20893 2078 20927
rect 3249 20893 3283 20927
rect 3433 20893 3467 20927
rect 4353 20893 4387 20927
rect 4813 20893 4847 20927
rect 4997 20893 5031 20927
rect 5181 20893 5215 20927
rect 6009 20893 6043 20927
rect 6193 20893 6227 20927
rect 8677 20893 8711 20927
rect 9505 20893 9539 20927
rect 11897 20893 11931 20927
rect 12541 20893 12575 20927
rect 13185 20893 13219 20927
rect 14105 20893 14139 20927
rect 16957 20893 16991 20927
rect 17233 20893 17267 20927
rect 17785 20893 17819 20927
rect 17969 20893 18003 20927
rect 18153 20893 18187 20927
rect 19809 20893 19843 20927
rect 20545 20893 20579 20927
rect 20913 20893 20947 20927
rect 25789 20893 25823 20927
rect 26249 20893 26283 20927
rect 28457 20893 28491 20927
rect 28733 20893 28767 20927
rect 28825 20893 28859 20927
rect 29929 20893 29963 20927
rect 30748 20893 30782 20927
rect 32229 20893 32263 20927
rect 32496 20893 32530 20927
rect 36286 20893 36320 20927
rect 36553 20893 36587 20927
rect 37289 20893 37323 20927
rect 37556 20893 37590 20927
rect 4537 20825 4571 20859
rect 6653 20825 6687 20859
rect 9772 20825 9806 20859
rect 14372 20825 14406 20859
rect 15945 20825 15979 20859
rect 16405 20825 16439 20859
rect 18061 20825 18095 20859
rect 19993 20825 20027 20859
rect 21180 20825 21214 20859
rect 24777 20825 24811 20859
rect 25237 20825 25271 20859
rect 26494 20825 26528 20859
rect 28641 20825 28675 20859
rect 40693 20825 40727 20859
rect 3341 20757 3375 20791
rect 3801 20757 3835 20791
rect 4721 20757 4755 20791
rect 10977 20757 11011 20791
rect 12265 20757 12299 20791
rect 15577 20757 15611 20791
rect 19073 20757 19107 20791
rect 24409 20757 24443 20791
rect 27721 20757 27755 20791
rect 29561 20757 29595 20791
rect 31861 20757 31895 20791
rect 33609 20757 33643 20791
rect 35173 20757 35207 20791
rect 38761 20757 38795 20791
rect 39129 20757 39163 20791
rect 42165 20757 42199 20791
rect 3065 20553 3099 20587
rect 4537 20553 4571 20587
rect 6377 20553 6411 20587
rect 9781 20553 9815 20587
rect 13277 20553 13311 20587
rect 18429 20553 18463 20587
rect 22293 20553 22327 20587
rect 24869 20553 24903 20587
rect 26157 20553 26191 20587
rect 27813 20553 27847 20587
rect 40233 20553 40267 20587
rect 41153 20553 41187 20587
rect 41613 20553 41647 20587
rect 8401 20485 8435 20519
rect 12164 20485 12198 20519
rect 14740 20485 14774 20519
rect 18972 20485 19006 20519
rect 23397 20485 23431 20519
rect 25881 20485 25915 20519
rect 32873 20485 32907 20519
rect 32965 20485 32999 20519
rect 36277 20485 36311 20519
rect 40785 20485 40819 20519
rect 1593 20417 1627 20451
rect 1860 20417 1894 20451
rect 3433 20417 3467 20451
rect 4629 20417 4663 20451
rect 6745 20417 6779 20451
rect 9137 20417 9171 20451
rect 9413 20417 9447 20451
rect 11897 20417 11931 20451
rect 16129 20417 16163 20451
rect 16681 20417 16715 20451
rect 21649 20417 21683 20451
rect 22201 20417 22235 20451
rect 25605 20417 25639 20451
rect 25789 20417 25823 20451
rect 25973 20417 26007 20451
rect 28365 20417 28399 20451
rect 32689 20417 32723 20451
rect 33057 20417 33091 20451
rect 35193 20417 35227 20451
rect 35449 20417 35483 20451
rect 37289 20417 37323 20451
rect 37556 20417 37590 20451
rect 38853 20417 38887 20451
rect 39120 20417 39154 20451
rect 40693 20417 40727 20451
rect 41521 20417 41555 20451
rect 3341 20349 3375 20383
rect 3893 20349 3927 20383
rect 6653 20349 6687 20383
rect 9321 20349 9355 20383
rect 14473 20349 14507 20383
rect 16221 20349 16255 20383
rect 16957 20349 16991 20383
rect 18705 20349 18739 20383
rect 21097 20349 21131 20383
rect 22385 20349 22419 20383
rect 23121 20349 23155 20383
rect 27905 20349 27939 20383
rect 28089 20349 28123 20383
rect 28641 20349 28675 20383
rect 30113 20349 30147 20383
rect 33333 20349 33367 20383
rect 35541 20349 35575 20383
rect 36921 20349 36955 20383
rect 40877 20349 40911 20383
rect 41705 20349 41739 20383
rect 15853 20281 15887 20315
rect 40325 20281 40359 20315
rect 2973 20213 3007 20247
rect 5273 20213 5307 20247
rect 6745 20213 6779 20247
rect 16497 20213 16531 20247
rect 20085 20213 20119 20247
rect 21833 20213 21867 20247
rect 27445 20213 27479 20247
rect 33241 20213 33275 20247
rect 33977 20213 34011 20247
rect 34069 20213 34103 20247
rect 36185 20213 36219 20247
rect 38669 20213 38703 20247
rect 3617 20009 3651 20043
rect 4261 20009 4295 20043
rect 5825 20009 5859 20043
rect 11437 20009 11471 20043
rect 17325 20009 17359 20043
rect 19257 20009 19291 20043
rect 19717 20009 19751 20043
rect 36185 20009 36219 20043
rect 10517 19941 10551 19975
rect 32413 19941 32447 19975
rect 5641 19873 5675 19907
rect 8217 19873 8251 19907
rect 8953 19873 8987 19907
rect 11989 19873 12023 19907
rect 17877 19873 17911 19907
rect 18705 19873 18739 19907
rect 22017 19873 22051 19907
rect 26617 19873 26651 19907
rect 32965 19873 32999 19907
rect 33057 19873 33091 19907
rect 33333 19873 33367 19907
rect 38853 19873 38887 19907
rect 39957 19873 39991 19907
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 3985 19805 4019 19839
rect 4169 19805 4203 19839
rect 5733 19805 5767 19839
rect 5917 19805 5951 19839
rect 6745 19805 6779 19839
rect 8125 19805 8159 19839
rect 8309 19805 8343 19839
rect 8493 19805 8527 19839
rect 8585 19805 8619 19839
rect 10885 19805 10919 19839
rect 11345 19805 11379 19839
rect 11529 19805 11563 19839
rect 11621 19805 11655 19839
rect 14841 19805 14875 19839
rect 15485 19805 15519 19839
rect 19441 19805 19475 19839
rect 19533 19805 19567 19839
rect 19809 19805 19843 19839
rect 22293 19805 22327 19839
rect 23305 19805 23339 19839
rect 24041 19805 24075 19839
rect 31033 19805 31067 19839
rect 34713 19805 34747 19839
rect 34969 19805 35003 19839
rect 36369 19805 36403 19839
rect 36461 19805 36495 19839
rect 36737 19805 36771 19839
rect 39037 19805 39071 19839
rect 2504 19737 2538 19771
rect 3801 19737 3835 19771
rect 5374 19737 5408 19771
rect 6377 19737 6411 19771
rect 6653 19737 6687 19771
rect 7113 19737 7147 19771
rect 8769 19737 8803 19771
rect 9198 19737 9232 19771
rect 12256 19737 12290 19771
rect 14105 19737 14139 19771
rect 15761 19737 15795 19771
rect 17693 19737 17727 19771
rect 18153 19737 18187 19771
rect 22477 19737 22511 19771
rect 26893 19737 26927 19771
rect 31300 19737 31334 19771
rect 36553 19737 36587 19771
rect 38577 19737 38611 19771
rect 40233 19737 40267 19771
rect 6561 19669 6595 19703
rect 6929 19669 6963 19703
rect 7205 19669 7239 19703
rect 10333 19669 10367 19703
rect 10425 19669 10459 19703
rect 11805 19669 11839 19703
rect 13369 19669 13403 19703
rect 17233 19669 17267 19703
rect 17785 19669 17819 19703
rect 20545 19669 20579 19703
rect 23489 19669 23523 19703
rect 28365 19669 28399 19703
rect 32505 19669 32539 19703
rect 32873 19669 32907 19703
rect 33977 19669 34011 19703
rect 36093 19669 36127 19703
rect 37105 19669 37139 19703
rect 39589 19669 39623 19703
rect 41705 19669 41739 19703
rect 1777 19465 1811 19499
rect 9689 19465 9723 19499
rect 11161 19465 11195 19499
rect 12449 19465 12483 19499
rect 16681 19465 16715 19499
rect 17141 19465 17175 19499
rect 25605 19465 25639 19499
rect 26433 19465 26467 19499
rect 31585 19465 31619 19499
rect 32137 19465 32171 19499
rect 36829 19465 36863 19499
rect 38485 19465 38519 19499
rect 40233 19465 40267 19499
rect 40693 19465 40727 19499
rect 41521 19465 41555 19499
rect 2513 19397 2547 19431
rect 3249 19397 3283 19431
rect 8677 19397 8711 19431
rect 8861 19397 8895 19431
rect 10048 19397 10082 19431
rect 17049 19397 17083 19431
rect 34345 19397 34379 19431
rect 34437 19397 34471 19431
rect 38025 19397 38059 19431
rect 1961 19329 1995 19363
rect 3801 19329 3835 19363
rect 4261 19329 4295 19363
rect 4813 19329 4847 19363
rect 4997 19329 5031 19363
rect 5181 19329 5215 19363
rect 6009 19329 6043 19363
rect 6653 19329 6687 19363
rect 6920 19329 6954 19363
rect 9045 19329 9079 19363
rect 9321 19329 9355 19363
rect 9781 19329 9815 19363
rect 11713 19329 11747 19363
rect 11897 19329 11931 19363
rect 12265 19329 12299 19363
rect 13737 19329 13771 19363
rect 17693 19329 17727 19363
rect 19901 19329 19935 19363
rect 22017 19329 22051 19363
rect 23857 19329 23891 19363
rect 26341 19329 26375 19363
rect 26985 19329 27019 19363
rect 27997 19329 28031 19363
rect 29837 19329 29871 19363
rect 33885 19329 33919 19363
rect 38117 19329 38151 19363
rect 40601 19329 40635 19363
rect 41061 19329 41095 19363
rect 41245 19329 41279 19363
rect 2145 19261 2179 19295
rect 3893 19261 3927 19295
rect 4169 19261 4203 19295
rect 5089 19261 5123 19295
rect 5733 19261 5767 19295
rect 5825 19261 5859 19295
rect 5917 19261 5951 19295
rect 9229 19261 9263 19295
rect 9413 19261 9447 19295
rect 9505 19261 9539 19295
rect 11989 19261 12023 19295
rect 12081 19261 12115 19295
rect 17325 19261 17359 19295
rect 17969 19261 18003 19295
rect 19441 19261 19475 19295
rect 20177 19261 20211 19295
rect 21649 19261 21683 19295
rect 22293 19261 22327 19295
rect 24133 19261 24167 19295
rect 26525 19261 26559 19295
rect 27537 19261 27571 19295
rect 28273 19261 28307 19295
rect 29745 19261 29779 19295
rect 30113 19261 30147 19295
rect 33609 19261 33643 19295
rect 34621 19261 34655 19295
rect 35081 19261 35115 19295
rect 35357 19261 35391 19295
rect 37933 19261 37967 19295
rect 40785 19261 40819 19295
rect 42165 19261 42199 19295
rect 23765 19193 23799 19227
rect 33977 19193 34011 19227
rect 6193 19125 6227 19159
rect 8033 19125 8067 19159
rect 25973 19125 26007 19159
rect 41153 19125 41187 19159
rect 4077 18921 4111 18955
rect 4537 18921 4571 18955
rect 6837 18921 6871 18955
rect 10149 18921 10183 18955
rect 10885 18921 10919 18955
rect 17877 18921 17911 18955
rect 18337 18921 18371 18955
rect 19441 18921 19475 18955
rect 20729 18921 20763 18955
rect 22753 18921 22787 18955
rect 24409 18921 24443 18955
rect 26709 18921 26743 18955
rect 28457 18921 28491 18955
rect 30481 18921 30515 18955
rect 34345 18921 34379 18955
rect 38301 18921 38335 18955
rect 41245 18921 41279 18955
rect 6653 18853 6687 18887
rect 7205 18853 7239 18887
rect 9597 18853 9631 18887
rect 12173 18853 12207 18887
rect 40233 18853 40267 18887
rect 3893 18785 3927 18819
rect 8125 18785 8159 18819
rect 8309 18785 8343 18819
rect 12357 18785 12391 18819
rect 12541 18785 12575 18819
rect 17233 18785 17267 18819
rect 18981 18785 19015 18819
rect 21281 18785 21315 18819
rect 23213 18785 23247 18819
rect 23305 18785 23339 18819
rect 24961 18785 24995 18819
rect 29009 18785 29043 18819
rect 31033 18785 31067 18819
rect 34989 18785 35023 18819
rect 37657 18785 37691 18819
rect 41797 18785 41831 18819
rect 3801 18717 3835 18751
rect 4077 18717 4111 18751
rect 7573 18717 7607 18751
rect 8401 18717 8435 18751
rect 9781 18717 9815 18751
rect 10885 18717 10919 18751
rect 11069 18717 11103 18751
rect 12081 18717 12115 18751
rect 12265 18717 12299 18751
rect 12633 18717 12667 18751
rect 12726 18717 12760 18751
rect 12817 18717 12851 18751
rect 13277 18717 13311 18751
rect 13369 18717 13403 18751
rect 13553 18717 13587 18751
rect 13645 18717 13679 18751
rect 13829 18717 13863 18751
rect 18705 18717 18739 18751
rect 21097 18717 21131 18751
rect 23121 18717 23155 18751
rect 25329 18717 25363 18751
rect 25596 18717 25630 18751
rect 28825 18717 28859 18751
rect 30849 18717 30883 18751
rect 32137 18717 32171 18751
rect 32597 18717 32631 18751
rect 39313 18717 39347 18751
rect 40049 18717 40083 18751
rect 40233 18717 40267 18751
rect 40969 18717 41003 18751
rect 4353 18649 4387 18683
rect 4553 18649 4587 18683
rect 7757 18649 7791 18683
rect 9965 18649 9999 18683
rect 11345 18649 11379 18683
rect 13001 18649 13035 18683
rect 13185 18649 13219 18683
rect 19717 18649 19751 18683
rect 24869 18649 24903 18683
rect 32873 18649 32907 18683
rect 35265 18649 35299 18683
rect 4261 18581 4295 18615
rect 4721 18581 4755 18615
rect 6837 18581 6871 18615
rect 7389 18581 7423 18615
rect 8125 18581 8159 18615
rect 9873 18581 9907 18615
rect 10701 18581 10735 18615
rect 13737 18581 13771 18615
rect 18797 18581 18831 18615
rect 21189 18581 21223 18615
rect 24777 18581 24811 18615
rect 28917 18581 28951 18615
rect 30941 18581 30975 18615
rect 36737 18581 36771 18615
rect 38669 18581 38703 18615
rect 40325 18581 40359 18615
rect 8309 18377 8343 18411
rect 11069 18377 11103 18411
rect 17141 18377 17175 18411
rect 19901 18377 19935 18411
rect 21465 18377 21499 18411
rect 26341 18377 26375 18411
rect 33425 18377 33459 18411
rect 33793 18377 33827 18411
rect 35817 18377 35851 18411
rect 36185 18377 36219 18411
rect 41613 18377 41647 18411
rect 9873 18309 9907 18343
rect 14206 18309 14240 18343
rect 27721 18309 27755 18343
rect 28089 18309 28123 18343
rect 32873 18309 32907 18343
rect 36277 18309 36311 18343
rect 40141 18309 40175 18343
rect 42165 18309 42199 18343
rect 1409 18241 1443 18275
rect 7849 18241 7883 18275
rect 9229 18241 9263 18275
rect 9597 18241 9631 18275
rect 10057 18241 10091 18275
rect 10149 18241 10183 18275
rect 10609 18241 10643 18275
rect 10885 18241 10919 18275
rect 12081 18241 12115 18275
rect 12449 18241 12483 18275
rect 14473 18241 14507 18275
rect 17049 18241 17083 18275
rect 18153 18241 18187 18275
rect 21373 18241 21407 18275
rect 26249 18241 26283 18275
rect 26985 18241 27019 18275
rect 28733 18241 28767 18275
rect 31677 18241 31711 18275
rect 32137 18241 32171 18275
rect 33885 18241 33919 18275
rect 8033 18173 8067 18207
rect 8861 18173 8895 18207
rect 9137 18173 9171 18207
rect 10701 18173 10735 18207
rect 12541 18173 12575 18207
rect 17325 18173 17359 18207
rect 18429 18173 18463 18207
rect 22385 18173 22419 18207
rect 26433 18173 26467 18207
rect 27537 18173 27571 18207
rect 29009 18173 29043 18207
rect 34069 18173 34103 18207
rect 36461 18173 36495 18207
rect 37565 18173 37599 18207
rect 37841 18173 37875 18207
rect 39865 18173 39899 18207
rect 10333 18105 10367 18139
rect 11897 18105 11931 18139
rect 13093 18105 13127 18139
rect 21833 18105 21867 18139
rect 41797 18105 41831 18139
rect 1593 18037 1627 18071
rect 7665 18037 7699 18071
rect 9597 18037 9631 18071
rect 9781 18037 9815 18071
rect 9873 18037 9907 18071
rect 10885 18037 10919 18071
rect 12173 18037 12207 18071
rect 16681 18037 16715 18071
rect 25881 18037 25915 18071
rect 30481 18037 30515 18071
rect 31401 18037 31435 18071
rect 39313 18037 39347 18071
rect 41705 18037 41739 18071
rect 5733 17833 5767 17867
rect 10333 17833 10367 17867
rect 10425 17833 10459 17867
rect 10885 17833 10919 17867
rect 19257 17833 19291 17867
rect 24409 17833 24443 17867
rect 26985 17833 27019 17867
rect 35725 17833 35759 17867
rect 41613 17833 41647 17867
rect 14105 17765 14139 17799
rect 16957 17765 16991 17799
rect 22385 17765 22419 17799
rect 1777 17697 1811 17731
rect 4905 17697 4939 17731
rect 6101 17697 6135 17731
rect 10241 17697 10275 17731
rect 12541 17697 12575 17731
rect 12817 17697 12851 17731
rect 13921 17697 13955 17731
rect 17509 17697 17543 17731
rect 17693 17697 17727 17731
rect 18429 17697 18463 17731
rect 19809 17697 19843 17731
rect 20637 17697 20671 17731
rect 24225 17697 24259 17731
rect 24961 17697 24995 17731
rect 25237 17697 25271 17731
rect 25513 17697 25547 17731
rect 30849 17697 30883 17731
rect 32597 17697 32631 17731
rect 33241 17697 33275 17731
rect 36369 17697 36403 17731
rect 39405 17697 39439 17731
rect 40417 17697 40451 17731
rect 40969 17697 41003 17731
rect 41521 17697 41555 17731
rect 1409 17629 1443 17663
rect 3203 17629 3237 17663
rect 4353 17629 4387 17663
rect 5089 17629 5123 17663
rect 5181 17629 5215 17663
rect 5917 17629 5951 17663
rect 6009 17629 6043 17663
rect 6193 17629 6227 17663
rect 6377 17629 6411 17663
rect 7113 17629 7147 17663
rect 10057 17629 10091 17663
rect 10609 17629 10643 17663
rect 10977 17629 11011 17663
rect 15485 17629 15519 17663
rect 15577 17629 15611 17663
rect 15844 17629 15878 17663
rect 17877 17629 17911 17663
rect 19625 17629 19659 17663
rect 22477 17629 22511 17663
rect 27077 17629 27111 17663
rect 29193 17629 29227 17663
rect 29377 17629 29411 17663
rect 30297 17629 30331 17663
rect 30573 17629 30607 17663
rect 30757 17629 30791 17663
rect 33425 17629 33459 17663
rect 33609 17629 33643 17663
rect 36553 17629 36587 17663
rect 37105 17629 37139 17663
rect 37657 17629 37691 17663
rect 41797 17629 41831 17663
rect 41981 17629 42015 17663
rect 42165 17629 42199 17663
rect 5273 17561 5307 17595
rect 5641 17561 5675 17595
rect 7380 17561 7414 17595
rect 10333 17561 10367 17595
rect 12332 17561 12366 17595
rect 15218 17561 15252 17595
rect 20913 17561 20947 17595
rect 22753 17561 22787 17595
rect 27353 17561 27387 17595
rect 31125 17561 31159 17595
rect 32689 17561 32723 17595
rect 35357 17561 35391 17595
rect 35541 17561 35575 17595
rect 36093 17561 36127 17595
rect 37933 17561 37967 17595
rect 41889 17561 41923 17595
rect 3801 17493 3835 17527
rect 8493 17493 8527 17527
rect 9873 17493 9907 17527
rect 12173 17493 12207 17527
rect 12449 17493 12483 17527
rect 13277 17493 13311 17527
rect 17049 17493 17083 17527
rect 17417 17493 17451 17527
rect 19717 17493 19751 17527
rect 28825 17493 28859 17527
rect 29285 17493 29319 17527
rect 29653 17493 29687 17527
rect 30389 17493 30423 17527
rect 33517 17493 33551 17527
rect 35173 17493 35207 17527
rect 36185 17493 36219 17527
rect 39865 17493 39899 17527
rect 4491 17289 4525 17323
rect 5181 17289 5215 17323
rect 6101 17289 6135 17323
rect 7481 17289 7515 17323
rect 10517 17289 10551 17323
rect 12541 17289 12575 17323
rect 13001 17289 13035 17323
rect 17509 17289 17543 17323
rect 27905 17289 27939 17323
rect 29377 17289 29411 17323
rect 30297 17289 30331 17323
rect 31125 17289 31159 17323
rect 34621 17289 34655 17323
rect 37933 17289 37967 17323
rect 38577 17289 38611 17323
rect 41981 17289 42015 17323
rect 6929 17221 6963 17255
rect 23765 17221 23799 17255
rect 24409 17221 24443 17255
rect 28273 17221 28307 17255
rect 28411 17221 28445 17255
rect 29285 17221 29319 17255
rect 29745 17221 29779 17255
rect 30665 17221 30699 17255
rect 33701 17221 33735 17255
rect 34437 17221 34471 17255
rect 35541 17221 35575 17255
rect 38853 17221 38887 17255
rect 38945 17221 38979 17255
rect 39773 17221 39807 17255
rect 41153 17221 41187 17255
rect 1409 17153 1443 17187
rect 3065 17153 3099 17187
rect 4905 17153 4939 17187
rect 5089 17153 5123 17187
rect 5549 17153 5583 17187
rect 6009 17153 6043 17187
rect 6193 17153 6227 17187
rect 6653 17153 6687 17187
rect 7205 17153 7239 17187
rect 7389 17153 7423 17187
rect 7573 17153 7607 17187
rect 8116 17153 8150 17187
rect 9413 17153 9447 17187
rect 9505 17153 9539 17187
rect 9873 17153 9907 17187
rect 10701 17153 10735 17187
rect 10977 17153 11011 17187
rect 12173 17153 12207 17187
rect 12449 17153 12483 17187
rect 12725 17153 12759 17187
rect 14114 17153 14148 17187
rect 19901 17153 19935 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 22385 17153 22419 17187
rect 23673 17153 23707 17187
rect 23857 17153 23891 17187
rect 24041 17153 24075 17187
rect 24133 17153 24167 17187
rect 27445 17153 27479 17187
rect 27629 17153 27663 17187
rect 28089 17153 28123 17187
rect 28181 17153 28215 17187
rect 28733 17153 28767 17187
rect 29561 17153 29595 17187
rect 29653 17153 29687 17187
rect 29929 17153 29963 17187
rect 30205 17153 30239 17187
rect 30481 17153 30515 17187
rect 30757 17153 30791 17187
rect 30849 17153 30883 17187
rect 32137 17153 32171 17187
rect 32689 17153 32723 17187
rect 32965 17153 32999 17187
rect 33149 17153 33183 17187
rect 33241 17153 33275 17187
rect 33609 17153 33643 17187
rect 33793 17153 33827 17187
rect 34253 17153 34287 17187
rect 34529 17153 34563 17187
rect 34805 17153 34839 17187
rect 34897 17153 34931 17187
rect 34989 17153 35023 17187
rect 35173 17153 35207 17187
rect 37473 17153 37507 17187
rect 38117 17153 38151 17187
rect 38209 17153 38243 17187
rect 38301 17153 38335 17187
rect 38485 17153 38519 17187
rect 38761 17153 38795 17187
rect 39129 17153 39163 17187
rect 39589 17153 39623 17187
rect 39865 17153 39899 17187
rect 39957 17153 39991 17187
rect 41797 17153 41831 17187
rect 41889 17153 41923 17187
rect 42073 17153 42107 17187
rect 2697 17085 2731 17119
rect 5641 17085 5675 17119
rect 5825 17085 5859 17119
rect 6377 17085 6411 17119
rect 6929 17085 6963 17119
rect 7849 17085 7883 17119
rect 10793 17085 10827 17119
rect 14381 17085 14415 17119
rect 18153 17085 18187 17119
rect 20177 17085 20211 17119
rect 25881 17085 25915 17119
rect 26525 17085 26559 17119
rect 28549 17085 28583 17119
rect 31677 17085 31711 17119
rect 32781 17085 32815 17119
rect 33517 17085 33551 17119
rect 35265 17085 35299 17119
rect 37565 17085 37599 17119
rect 40417 17085 40451 17119
rect 6837 17017 6871 17051
rect 10057 17017 10091 17051
rect 12265 17017 12299 17051
rect 21649 17017 21683 17051
rect 23489 17017 23523 17051
rect 25973 17017 26007 17051
rect 31033 17017 31067 17051
rect 32873 17017 32907 17051
rect 33425 17017 33459 17051
rect 37841 17017 37875 17051
rect 40141 17017 40175 17051
rect 1593 16949 1627 16983
rect 4629 16949 4663 16983
rect 4905 16949 4939 16983
rect 6469 16949 6503 16983
rect 7113 16949 7147 16983
rect 9229 16949 9263 16983
rect 9873 16949 9907 16983
rect 10701 16949 10735 16983
rect 12909 16949 12943 16983
rect 21925 16949 21959 16983
rect 23029 16949 23063 16983
rect 27813 16949 27847 16983
rect 32321 16949 32355 16983
rect 32505 16949 32539 16983
rect 33333 16949 33367 16983
rect 34345 16949 34379 16983
rect 37013 16949 37047 16983
rect 41061 16949 41095 16983
rect 5089 16745 5123 16779
rect 6285 16745 6319 16779
rect 8033 16745 8067 16779
rect 8217 16745 8251 16779
rect 8953 16745 8987 16779
rect 10793 16745 10827 16779
rect 10977 16745 11011 16779
rect 11437 16745 11471 16779
rect 12633 16745 12667 16779
rect 12817 16745 12851 16779
rect 13093 16745 13127 16779
rect 13277 16745 13311 16779
rect 13921 16745 13955 16779
rect 20821 16745 20855 16779
rect 23765 16745 23799 16779
rect 24409 16745 24443 16779
rect 25789 16745 25823 16779
rect 28917 16745 28951 16779
rect 34805 16745 34839 16779
rect 36001 16745 36035 16779
rect 5825 16677 5859 16711
rect 25145 16677 25179 16711
rect 29653 16677 29687 16711
rect 33057 16677 33091 16711
rect 36093 16677 36127 16711
rect 1777 16609 1811 16643
rect 3203 16609 3237 16643
rect 4353 16609 4387 16643
rect 5273 16609 5307 16643
rect 5365 16609 5399 16643
rect 5457 16609 5491 16643
rect 5549 16609 5583 16643
rect 5733 16609 5767 16643
rect 9321 16609 9355 16643
rect 10609 16609 10643 16643
rect 13645 16609 13679 16643
rect 15945 16609 15979 16643
rect 20637 16609 20671 16643
rect 22109 16609 22143 16643
rect 24133 16609 24167 16643
rect 25053 16609 25087 16643
rect 27629 16609 27663 16643
rect 27721 16609 27755 16643
rect 31677 16609 31711 16643
rect 32137 16609 32171 16643
rect 32689 16609 32723 16643
rect 35357 16609 35391 16643
rect 38853 16609 38887 16643
rect 39865 16609 39899 16643
rect 40233 16609 40267 16643
rect 40509 16609 40543 16643
rect 1409 16541 1443 16575
rect 4813 16541 4847 16575
rect 6009 16541 6043 16575
rect 6377 16541 6411 16575
rect 8493 16541 8527 16575
rect 9137 16541 9171 16575
rect 9229 16541 9263 16575
rect 9413 16541 9447 16575
rect 10793 16541 10827 16575
rect 11621 16541 11655 16575
rect 11713 16541 11747 16575
rect 11805 16541 11839 16575
rect 13553 16541 13587 16575
rect 15669 16541 15703 16575
rect 17509 16541 17543 16575
rect 18337 16541 18371 16575
rect 18521 16541 18555 16575
rect 18705 16541 18739 16575
rect 18797 16541 18831 16575
rect 19441 16541 19475 16575
rect 19809 16541 19843 16575
rect 20085 16541 20119 16575
rect 21005 16541 21039 16575
rect 21097 16541 21131 16575
rect 21373 16541 21407 16575
rect 21465 16541 21499 16575
rect 22385 16541 22419 16575
rect 22569 16541 22603 16575
rect 22753 16541 22787 16575
rect 24041 16541 24075 16575
rect 25329 16541 25363 16575
rect 25513 16541 25547 16575
rect 25697 16541 25731 16575
rect 25789 16541 25823 16575
rect 25967 16541 26001 16575
rect 26065 16541 26099 16575
rect 26249 16541 26283 16575
rect 28733 16541 28767 16575
rect 29101 16541 29135 16575
rect 29285 16541 29319 16575
rect 29377 16541 29411 16575
rect 29745 16541 29779 16575
rect 29837 16541 29871 16575
rect 32597 16541 32631 16575
rect 33977 16541 34011 16575
rect 34069 16541 34103 16575
rect 34437 16541 34471 16575
rect 35541 16541 35575 16575
rect 35817 16541 35851 16575
rect 36369 16541 36403 16575
rect 36553 16541 36587 16575
rect 38117 16541 38151 16575
rect 40049 16541 40083 16575
rect 40141 16541 40175 16575
rect 4905 16473 4939 16507
rect 5089 16473 5123 16507
rect 8401 16473 8435 16507
rect 10517 16473 10551 16507
rect 12449 16473 12483 16507
rect 12665 16473 12699 16507
rect 12909 16473 12943 16507
rect 13109 16473 13143 16507
rect 19533 16473 19567 16507
rect 19625 16473 19659 16507
rect 21189 16473 21223 16507
rect 22477 16473 22511 16507
rect 25421 16473 25455 16507
rect 27537 16473 27571 16507
rect 28181 16473 28215 16507
rect 29561 16473 29595 16507
rect 31401 16473 31435 16507
rect 31769 16473 31803 16507
rect 31953 16473 31987 16507
rect 33333 16473 33367 16507
rect 34161 16473 34195 16507
rect 34299 16473 34333 16507
rect 35633 16473 35667 16507
rect 3801 16405 3835 16439
rect 8201 16405 8235 16439
rect 8585 16405 8619 16439
rect 17417 16405 17451 16439
rect 18153 16405 18187 16439
rect 18429 16405 18463 16439
rect 18981 16405 19015 16439
rect 19257 16405 19291 16439
rect 22201 16405 22235 16439
rect 26065 16405 26099 16439
rect 27169 16405 27203 16439
rect 29929 16405 29963 16439
rect 32229 16405 32263 16439
rect 32873 16405 32907 16439
rect 33793 16405 33827 16439
rect 36277 16405 36311 16439
rect 39865 16405 39899 16439
rect 41981 16405 42015 16439
rect 5457 16201 5491 16235
rect 8585 16201 8619 16235
rect 15669 16201 15703 16235
rect 17693 16201 17727 16235
rect 21097 16201 21131 16235
rect 24133 16201 24167 16235
rect 24225 16201 24259 16235
rect 29377 16201 29411 16235
rect 31125 16201 31159 16235
rect 31217 16201 31251 16235
rect 35265 16201 35299 16235
rect 37749 16201 37783 16235
rect 5733 16133 5767 16167
rect 8737 16133 8771 16167
rect 8953 16133 8987 16167
rect 12541 16133 12575 16167
rect 15117 16133 15151 16167
rect 20203 16133 20237 16167
rect 23765 16133 23799 16167
rect 27261 16133 27295 16167
rect 31493 16133 31527 16167
rect 31585 16133 31619 16167
rect 33793 16133 33827 16167
rect 39773 16133 39807 16167
rect 1409 16065 1443 16099
rect 2973 16065 3007 16099
rect 4399 16065 4433 16099
rect 5365 16065 5399 16099
rect 5917 16065 5951 16099
rect 6101 16065 6135 16099
rect 11713 16065 11747 16099
rect 12357 16065 12391 16099
rect 12449 16065 12483 16099
rect 12725 16065 12759 16099
rect 12817 16065 12851 16099
rect 13001 16065 13035 16099
rect 14206 16065 14240 16099
rect 15209 16065 15243 16099
rect 15485 16065 15519 16099
rect 15761 16065 15795 16099
rect 17049 16065 17083 16099
rect 17141 16065 17175 16099
rect 17509 16065 17543 16099
rect 19901 16065 19935 16099
rect 19993 16065 20027 16099
rect 20085 16065 20119 16099
rect 20729 16065 20763 16099
rect 21833 16065 21867 16099
rect 22017 16065 22051 16099
rect 23949 16065 23983 16099
rect 24869 16065 24903 16099
rect 25053 16065 25087 16099
rect 29653 16065 29687 16099
rect 30481 16065 30515 16099
rect 31401 16065 31435 16099
rect 31769 16065 31803 16099
rect 33517 16065 33551 16099
rect 35357 16065 35391 16099
rect 35541 16065 35575 16099
rect 37657 16065 37691 16099
rect 38209 16065 38243 16099
rect 40048 16065 40082 16099
rect 40141 16065 40175 16099
rect 40601 16065 40635 16099
rect 41245 16065 41279 16099
rect 41613 16065 41647 16099
rect 41797 16065 41831 16099
rect 2605 15997 2639 16031
rect 11805 15997 11839 16031
rect 11897 15997 11931 16031
rect 11989 15997 12023 16031
rect 14473 15997 14507 16031
rect 16497 15997 16531 16031
rect 17325 15997 17359 16031
rect 17877 15997 17911 16031
rect 18153 15997 18187 16031
rect 20361 15997 20395 16031
rect 20637 15997 20671 16031
rect 21189 15997 21223 16031
rect 21649 15997 21683 16031
rect 21925 15997 21959 16031
rect 24685 15997 24719 16031
rect 24777 15997 24811 16031
rect 26985 15997 27019 16031
rect 29285 15997 29319 16031
rect 29377 15997 29411 16031
rect 35449 15997 35483 16031
rect 37933 15997 37967 16031
rect 38945 15997 38979 16031
rect 39497 15997 39531 16031
rect 40233 15997 40267 16031
rect 40509 15997 40543 16031
rect 41061 15997 41095 16031
rect 41521 15997 41555 16031
rect 13093 15929 13127 15963
rect 19717 15929 19751 15963
rect 21373 15929 21407 15963
rect 24409 15929 24443 15963
rect 28917 15929 28951 15963
rect 29561 15929 29595 15963
rect 41705 15929 41739 15963
rect 1593 15861 1627 15895
rect 8769 15861 8803 15895
rect 11529 15861 11563 15895
rect 12173 15861 12207 15895
rect 12909 15861 12943 15895
rect 15301 15861 15335 15895
rect 15853 15861 15887 15895
rect 16681 15861 16715 15895
rect 19625 15861 19659 15895
rect 25237 15861 25271 15895
rect 28733 15861 28767 15895
rect 28825 15861 28859 15895
rect 37289 15861 37323 15895
rect 41429 15861 41463 15895
rect 3571 15657 3605 15691
rect 5733 15657 5767 15691
rect 7665 15657 7699 15691
rect 8401 15657 8435 15691
rect 12265 15657 12299 15691
rect 13829 15657 13863 15691
rect 16773 15657 16807 15691
rect 18889 15657 18923 15691
rect 18981 15657 19015 15691
rect 19901 15657 19935 15691
rect 19993 15657 20027 15691
rect 20821 15657 20855 15691
rect 22293 15657 22327 15691
rect 24409 15657 24443 15691
rect 37013 15657 37047 15691
rect 37454 15657 37488 15691
rect 41613 15657 41647 15691
rect 5641 15589 5675 15623
rect 8309 15589 8343 15623
rect 10701 15589 10735 15623
rect 21097 15589 21131 15623
rect 22661 15589 22695 15623
rect 24685 15589 24719 15623
rect 25881 15589 25915 15623
rect 28917 15589 28951 15623
rect 29009 15589 29043 15623
rect 29561 15589 29595 15623
rect 1777 15521 1811 15555
rect 5365 15521 5399 15555
rect 7205 15521 7239 15555
rect 9781 15521 9815 15555
rect 10333 15521 10367 15555
rect 17141 15521 17175 15555
rect 18613 15521 18647 15555
rect 19073 15521 19107 15555
rect 21189 15521 21223 15555
rect 22109 15521 22143 15555
rect 31493 15521 31527 15555
rect 31677 15521 31711 15555
rect 35265 15521 35299 15555
rect 37197 15521 37231 15555
rect 38945 15521 38979 15555
rect 1409 15453 1443 15487
rect 2145 15453 2179 15487
rect 5273 15453 5307 15487
rect 7481 15453 7515 15487
rect 8125 15453 8159 15487
rect 8309 15453 8343 15487
rect 8585 15453 8619 15487
rect 8769 15453 8803 15487
rect 9873 15453 9907 15487
rect 10057 15453 10091 15487
rect 10885 15453 10919 15487
rect 12909 15453 12943 15487
rect 13093 15453 13127 15487
rect 13277 15453 13311 15487
rect 13369 15453 13403 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 15393 15453 15427 15487
rect 16865 15453 16899 15487
rect 18797 15453 18831 15487
rect 19349 15453 19383 15487
rect 20177 15453 20211 15487
rect 20366 15453 20400 15487
rect 21005 15453 21039 15487
rect 21281 15453 21315 15487
rect 21465 15453 21499 15487
rect 21863 15453 21897 15487
rect 22017 15453 22051 15487
rect 22385 15453 22419 15487
rect 22569 15453 22603 15487
rect 22753 15453 22787 15487
rect 22937 15453 22971 15487
rect 23121 15453 23155 15487
rect 24593 15453 24627 15487
rect 24777 15453 24811 15487
rect 24869 15453 24903 15487
rect 25053 15453 25087 15487
rect 25513 15453 25547 15487
rect 25697 15453 25731 15487
rect 25789 15453 25823 15487
rect 25966 15453 26000 15487
rect 26157 15453 26191 15487
rect 26801 15453 26835 15487
rect 26893 15453 26927 15487
rect 27629 15453 27663 15487
rect 28641 15453 28675 15487
rect 28825 15453 28859 15487
rect 29101 15453 29135 15487
rect 29561 15453 29595 15487
rect 29745 15453 29779 15487
rect 31861 15453 31895 15487
rect 39129 15453 39163 15487
rect 39589 15453 39623 15487
rect 40049 15453 40083 15487
rect 40141 15453 40175 15487
rect 40417 15453 40451 15487
rect 41429 15453 41463 15487
rect 7941 15385 7975 15419
rect 9965 15385 9999 15419
rect 11130 15385 11164 15419
rect 15660 15385 15694 15419
rect 19993 15385 20027 15419
rect 20269 15385 20303 15419
rect 26341 15385 26375 15419
rect 26525 15385 26559 15419
rect 27261 15385 27295 15419
rect 29285 15385 29319 15419
rect 31401 15385 31435 15419
rect 32505 15385 32539 15419
rect 35541 15385 35575 15419
rect 40233 15385 40267 15419
rect 40785 15385 40819 15419
rect 41889 15385 41923 15419
rect 1593 15317 1627 15351
rect 9137 15317 9171 15351
rect 10793 15317 10827 15351
rect 12357 15317 12391 15351
rect 21649 15317 21683 15351
rect 22109 15317 22143 15351
rect 23029 15317 23063 15351
rect 25605 15317 25639 15351
rect 27169 15317 27203 15351
rect 31033 15317 31067 15351
rect 39221 15317 39255 15351
rect 39313 15317 39347 15351
rect 39865 15317 39899 15351
rect 4491 15113 4525 15147
rect 4721 15113 4755 15147
rect 5441 15113 5475 15147
rect 6653 15113 6687 15147
rect 10149 15113 10183 15147
rect 13001 15113 13035 15147
rect 13553 15113 13587 15147
rect 16497 15113 16531 15147
rect 18153 15113 18187 15147
rect 19073 15113 19107 15147
rect 19809 15113 19843 15147
rect 20269 15113 20303 15147
rect 20729 15113 20763 15147
rect 26525 15113 26559 15147
rect 31861 15113 31895 15147
rect 32781 15113 32815 15147
rect 36001 15113 36035 15147
rect 36369 15113 36403 15147
rect 41889 15113 41923 15147
rect 5641 15045 5675 15079
rect 14666 15045 14700 15079
rect 20361 15045 20395 15079
rect 20545 15045 20579 15079
rect 22385 15045 22419 15079
rect 24777 15045 24811 15079
rect 26065 15045 26099 15079
rect 26249 15045 26283 15079
rect 28181 15045 28215 15079
rect 30748 15045 30782 15079
rect 35265 15045 35299 15079
rect 4629 14977 4663 15011
rect 4905 14977 4939 15011
rect 6101 14977 6135 15011
rect 6561 14977 6595 15011
rect 6837 14977 6871 15011
rect 8217 14977 8251 15011
rect 8933 14977 8967 15011
rect 12633 14977 12667 15011
rect 14933 14977 14967 15011
rect 15117 14977 15151 15011
rect 15384 14977 15418 15011
rect 16681 14977 16715 15011
rect 18061 14977 18095 15011
rect 18889 14977 18923 15011
rect 19073 14977 19107 15011
rect 19901 14977 19935 15011
rect 19993 14977 20027 15011
rect 21005 14977 21039 15011
rect 22109 14977 22143 15011
rect 22293 14977 22327 15011
rect 22477 14977 22511 15011
rect 24685 14977 24719 15011
rect 24869 14977 24903 15011
rect 25007 14977 25041 15011
rect 26433 14977 26467 15011
rect 26525 14977 26559 15011
rect 26709 14977 26743 15011
rect 27261 14977 27295 15011
rect 27445 14977 27479 15011
rect 28641 14977 28675 15011
rect 29101 14977 29135 15011
rect 29285 14977 29319 15011
rect 29377 14977 29411 15011
rect 29469 14977 29503 15011
rect 30481 14977 30515 15011
rect 32689 14977 32723 15011
rect 33241 14977 33275 15011
rect 34069 14977 34103 15011
rect 34253 14977 34287 15011
rect 34989 14977 35023 15011
rect 35173 14977 35207 15011
rect 35357 14977 35391 15011
rect 37473 14977 37507 15011
rect 40141 14977 40175 15011
rect 2697 14909 2731 14943
rect 3065 14909 3099 14943
rect 7573 14909 7607 14943
rect 8125 14909 8159 14943
rect 8585 14909 8619 14943
rect 8677 14909 8711 14943
rect 10701 14909 10735 14943
rect 12725 14909 12759 14943
rect 17417 14909 17451 14943
rect 18337 14909 18371 14943
rect 19165 14909 19199 14943
rect 21097 14909 21131 14943
rect 25145 14909 25179 14943
rect 25421 14909 25455 14943
rect 28733 14909 28767 14943
rect 29745 14909 29779 14943
rect 30297 14909 30331 14943
rect 32965 14909 32999 14943
rect 33885 14909 33919 14943
rect 36461 14909 36495 14943
rect 36553 14909 36587 14943
rect 37749 14909 37783 14943
rect 39221 14909 39255 14943
rect 39865 14909 39899 14943
rect 40417 14909 40451 14943
rect 5917 14841 5951 14875
rect 29009 14841 29043 14875
rect 29653 14841 29687 14875
rect 4905 14773 4939 14807
rect 5273 14773 5307 14807
rect 5457 14773 5491 14807
rect 10057 14773 10091 14807
rect 17693 14773 17727 14807
rect 19901 14773 19935 14807
rect 21281 14773 21315 14807
rect 22661 14773 22695 14807
rect 24501 14773 24535 14807
rect 25973 14773 26007 14807
rect 27169 14773 27203 14807
rect 32321 14773 32355 14807
rect 35541 14773 35575 14807
rect 39313 14773 39347 14807
rect 3801 14569 3835 14603
rect 5070 14569 5104 14603
rect 10333 14569 10367 14603
rect 17969 14569 18003 14603
rect 21925 14569 21959 14603
rect 26893 14569 26927 14603
rect 38025 14569 38059 14603
rect 39589 14569 39623 14603
rect 40877 14569 40911 14603
rect 41797 14569 41831 14603
rect 34529 14501 34563 14535
rect 39865 14501 39899 14535
rect 1409 14433 1443 14467
rect 4813 14433 4847 14467
rect 8953 14433 8987 14467
rect 10517 14433 10551 14467
rect 15945 14433 15979 14467
rect 17693 14433 17727 14467
rect 20545 14433 20579 14467
rect 23673 14433 23707 14467
rect 24961 14433 24995 14467
rect 28917 14433 28951 14467
rect 29561 14433 29595 14467
rect 29837 14433 29871 14467
rect 31953 14433 31987 14467
rect 32229 14433 32263 14467
rect 34253 14433 34287 14467
rect 38945 14433 38979 14467
rect 40233 14433 40267 14467
rect 1777 14365 1811 14399
rect 3203 14365 3237 14399
rect 4353 14365 4387 14399
rect 6929 14365 6963 14399
rect 9209 14365 9243 14399
rect 10701 14365 10735 14399
rect 10793 14365 10827 14399
rect 18613 14365 18647 14399
rect 18705 14365 18739 14399
rect 18889 14365 18923 14399
rect 19073 14365 19107 14399
rect 19441 14365 19475 14399
rect 19743 14365 19777 14399
rect 19901 14365 19935 14399
rect 21281 14365 21315 14399
rect 21373 14365 21407 14399
rect 21649 14365 21683 14399
rect 26801 14365 26835 14399
rect 26985 14365 27019 14399
rect 31493 14365 31527 14399
rect 34161 14365 34195 14399
rect 35173 14365 35207 14399
rect 38209 14365 38243 14399
rect 38393 14365 38427 14399
rect 38511 14365 38545 14399
rect 38669 14365 38703 14399
rect 39129 14365 39163 14399
rect 39313 14365 39347 14399
rect 39405 14365 39439 14399
rect 39497 14365 39531 14399
rect 39681 14365 39715 14399
rect 39865 14365 39899 14399
rect 39957 14365 39991 14399
rect 41521 14365 41555 14399
rect 10517 14297 10551 14331
rect 16221 14297 16255 14331
rect 19533 14297 19567 14331
rect 19625 14297 19659 14331
rect 21465 14297 21499 14331
rect 23397 14297 23431 14331
rect 25237 14297 25271 14331
rect 28641 14297 28675 14331
rect 31861 14297 31895 14331
rect 35817 14297 35851 14331
rect 38301 14297 38335 14331
rect 40141 14297 40175 14331
rect 6561 14229 6595 14263
rect 19257 14229 19291 14263
rect 19993 14229 20027 14263
rect 21097 14229 21131 14263
rect 26709 14229 26743 14263
rect 27169 14229 27203 14263
rect 31309 14229 31343 14263
rect 33701 14229 33735 14263
rect 2329 14025 2363 14059
rect 5825 14025 5859 14059
rect 6745 14025 6779 14059
rect 11713 14025 11747 14059
rect 11989 14025 12023 14059
rect 12173 14025 12207 14059
rect 18429 14025 18463 14059
rect 20269 14025 20303 14059
rect 22109 14025 22143 14059
rect 23765 14025 23799 14059
rect 25605 14025 25639 14059
rect 25697 14025 25731 14059
rect 26065 14025 26099 14059
rect 32505 14025 32539 14059
rect 34989 14025 35023 14059
rect 38301 14025 38335 14059
rect 38945 14025 38979 14059
rect 41061 14025 41095 14059
rect 5273 13957 5307 13991
rect 5473 13957 5507 13991
rect 6009 13957 6043 13991
rect 6653 13957 6687 13991
rect 9873 13957 9907 13991
rect 12725 13957 12759 13991
rect 24133 13957 24167 13991
rect 29101 13957 29135 13991
rect 36461 13957 36495 13991
rect 40049 13957 40083 13991
rect 1685 13889 1719 13923
rect 5733 13889 5767 13923
rect 9597 13889 9631 13923
rect 11529 13889 11563 13923
rect 11897 13889 11931 13923
rect 12081 13889 12115 13923
rect 12173 13889 12207 13923
rect 12357 13889 12391 13923
rect 12909 13889 12943 13923
rect 21005 13889 21039 13923
rect 23121 13889 23155 13923
rect 23857 13889 23891 13923
rect 27537 13889 27571 13923
rect 30205 13889 30239 13923
rect 34713 13889 34747 13923
rect 38209 13889 38243 13923
rect 38669 13889 38703 13923
rect 39865 13889 39899 13923
rect 40969 13889 41003 13923
rect 41521 13889 41555 13923
rect 2973 13821 3007 13855
rect 3065 13821 3099 13855
rect 3341 13821 3375 13855
rect 5089 13821 5123 13855
rect 16681 13821 16715 13855
rect 18521 13821 18555 13855
rect 18797 13821 18831 13855
rect 21649 13821 21683 13855
rect 22661 13821 22695 13855
rect 26157 13821 26191 13855
rect 26341 13821 26375 13855
rect 28365 13821 28399 13855
rect 28457 13821 28491 13855
rect 30481 13821 30515 13855
rect 31953 13821 31987 13855
rect 33977 13821 34011 13855
rect 34253 13821 34287 13855
rect 34621 13821 34655 13855
rect 36737 13821 36771 13855
rect 38945 13821 38979 13855
rect 40233 13821 40267 13855
rect 41153 13821 41187 13855
rect 42165 13821 42199 13855
rect 6009 13753 6043 13787
rect 34345 13753 34379 13787
rect 1501 13685 1535 13719
rect 5457 13685 5491 13719
rect 5641 13685 5675 13719
rect 11345 13685 11379 13719
rect 12541 13685 12575 13719
rect 16944 13685 16978 13719
rect 26985 13685 27019 13719
rect 27721 13685 27755 13719
rect 38761 13685 38795 13719
rect 40601 13685 40635 13719
rect 3203 13481 3237 13515
rect 5273 13481 5307 13515
rect 6561 13481 6595 13515
rect 8493 13481 8527 13515
rect 10977 13481 11011 13515
rect 15301 13481 15335 13515
rect 32597 13481 32631 13515
rect 38485 13481 38519 13515
rect 39405 13481 39439 13515
rect 42165 13481 42199 13515
rect 4997 13413 5031 13447
rect 19257 13413 19291 13447
rect 22017 13413 22051 13447
rect 23857 13413 23891 13447
rect 25237 13413 25271 13447
rect 27077 13413 27111 13447
rect 28089 13413 28123 13447
rect 33701 13413 33735 13447
rect 34713 13413 34747 13447
rect 37289 13413 37323 13447
rect 1777 13345 1811 13379
rect 8309 13345 8343 13379
rect 17601 13345 17635 13379
rect 17785 13345 17819 13379
rect 20269 13345 20303 13379
rect 20545 13345 20579 13379
rect 22109 13345 22143 13379
rect 25605 13345 25639 13379
rect 33057 13345 33091 13379
rect 34345 13345 34379 13379
rect 35541 13345 35575 13379
rect 40417 13345 40451 13379
rect 40693 13345 40727 13379
rect 1409 13277 1443 13311
rect 4721 13277 4755 13311
rect 5089 13277 5123 13311
rect 5273 13277 5307 13311
rect 5825 13277 5859 13311
rect 6009 13277 6043 13311
rect 6285 13277 6319 13311
rect 8401 13277 8435 13311
rect 10885 13277 10919 13311
rect 11161 13277 11195 13311
rect 11253 13277 11287 13311
rect 11897 13277 11931 13311
rect 14657 13277 14691 13311
rect 17049 13277 17083 13311
rect 19441 13277 19475 13311
rect 19809 13277 19843 13311
rect 24685 13277 24719 13311
rect 24961 13277 24995 13311
rect 25053 13277 25087 13311
rect 25329 13277 25363 13311
rect 27537 13277 27571 13311
rect 27721 13277 27755 13311
rect 27905 13277 27939 13311
rect 28733 13277 28767 13311
rect 31125 13277 31159 13311
rect 34897 13277 34931 13311
rect 34989 13277 35023 13311
rect 35081 13277 35115 13311
rect 35265 13277 35299 13311
rect 37473 13277 37507 13311
rect 38669 13277 38703 13311
rect 38945 13277 38979 13311
rect 39129 13277 39163 13311
rect 39221 13277 39255 13311
rect 39405 13277 39439 13311
rect 4997 13209 5031 13243
rect 6101 13209 6135 13243
rect 8033 13209 8067 13243
rect 12173 13209 12207 13243
rect 16773 13209 16807 13243
rect 19533 13209 19567 13243
rect 19625 13209 19659 13243
rect 22385 13209 22419 13243
rect 24869 13209 24903 13243
rect 27813 13209 27847 13243
rect 28549 13209 28583 13243
rect 35817 13209 35851 13243
rect 4813 13141 4847 13175
rect 6009 13141 6043 13175
rect 6469 13141 6503 13175
rect 9597 13141 9631 13175
rect 11621 13141 11655 13175
rect 13645 13141 13679 13175
rect 14105 13141 14139 13175
rect 17141 13141 17175 13175
rect 17509 13141 17543 13175
rect 28273 13141 28307 13175
rect 28917 13141 28951 13175
rect 33609 13141 33643 13175
rect 39589 13141 39623 13175
rect 4813 12937 4847 12971
rect 6761 12937 6795 12971
rect 6929 12937 6963 12971
rect 18613 12937 18647 12971
rect 22477 12937 22511 12971
rect 22937 12937 22971 12971
rect 29009 12937 29043 12971
rect 29469 12937 29503 12971
rect 32137 12937 32171 12971
rect 32505 12937 32539 12971
rect 33425 12937 33459 12971
rect 35449 12937 35483 12971
rect 36185 12937 36219 12971
rect 36553 12937 36587 12971
rect 40877 12937 40911 12971
rect 6561 12869 6595 12903
rect 9137 12869 9171 12903
rect 13261 12869 13295 12903
rect 13461 12869 13495 12903
rect 19073 12869 19107 12903
rect 26065 12869 26099 12903
rect 32597 12869 32631 12903
rect 38853 12869 38887 12903
rect 4077 12801 4111 12835
rect 4261 12801 4295 12835
rect 5365 12801 5399 12835
rect 8861 12801 8895 12835
rect 9045 12801 9079 12835
rect 10057 12801 10091 12835
rect 10211 12801 10245 12835
rect 10885 12801 10919 12835
rect 12633 12801 12667 12835
rect 13001 12801 13035 12835
rect 15301 12801 15335 12835
rect 18613 12801 18647 12835
rect 18797 12801 18831 12835
rect 19533 12801 19567 12835
rect 19901 12801 19935 12835
rect 22845 12801 22879 12835
rect 25237 12801 25271 12835
rect 27445 12801 27479 12835
rect 27629 12801 27663 12835
rect 27721 12801 27755 12835
rect 27997 12801 28031 12835
rect 28181 12801 28215 12835
rect 28825 12801 28859 12835
rect 29101 12801 29135 12835
rect 29285 12801 29319 12835
rect 33333 12801 33367 12835
rect 33793 12801 33827 12835
rect 35633 12801 35667 12835
rect 35725 12801 35759 12835
rect 36645 12801 36679 12835
rect 39497 12801 39531 12835
rect 41061 12801 41095 12835
rect 1501 12733 1535 12767
rect 1777 12733 1811 12767
rect 3249 12733 3283 12767
rect 3893 12733 3927 12767
rect 5089 12733 5123 12767
rect 10425 12733 10459 12767
rect 10977 12733 11011 12767
rect 11161 12733 11195 12767
rect 11529 12733 11563 12767
rect 12081 12733 12115 12767
rect 12541 12733 12575 12767
rect 12909 12733 12943 12767
rect 15025 12733 15059 12767
rect 23121 12733 23155 12767
rect 28457 12733 28491 12767
rect 31125 12733 31159 12767
rect 31401 12733 31435 12767
rect 32781 12733 32815 12767
rect 33517 12733 33551 12767
rect 34345 12733 34379 12767
rect 35081 12733 35115 12767
rect 36737 12733 36771 12767
rect 37381 12733 37415 12767
rect 39129 12733 39163 12767
rect 39221 12733 39255 12767
rect 40693 12733 40727 12767
rect 41245 12733 41279 12767
rect 3341 12665 3375 12699
rect 8769 12665 8803 12699
rect 12357 12665 12391 12699
rect 27905 12665 27939 12699
rect 4077 12597 4111 12631
rect 5181 12597 5215 12631
rect 6745 12597 6779 12631
rect 10517 12597 10551 12631
rect 13093 12597 13127 12631
rect 13277 12597 13311 12631
rect 13553 12597 13587 12631
rect 18981 12597 19015 12631
rect 27813 12597 27847 12631
rect 28641 12597 28675 12631
rect 29653 12597 29687 12631
rect 32965 12597 32999 12631
rect 34529 12597 34563 12631
rect 35909 12597 35943 12631
rect 40141 12597 40175 12631
rect 1593 12393 1627 12427
rect 5181 12393 5215 12427
rect 5733 12393 5767 12427
rect 6653 12393 6687 12427
rect 11253 12393 11287 12427
rect 11437 12393 11471 12427
rect 12541 12393 12575 12427
rect 14105 12393 14139 12427
rect 17785 12393 17819 12427
rect 22201 12393 22235 12427
rect 24133 12393 24167 12427
rect 29285 12393 29319 12427
rect 30665 12393 30699 12427
rect 32965 12393 32999 12427
rect 34345 12393 34379 12427
rect 3801 12325 3835 12359
rect 6285 12325 6319 12359
rect 11161 12325 11195 12359
rect 12357 12325 12391 12359
rect 13921 12325 13955 12359
rect 20177 12325 20211 12359
rect 34529 12325 34563 12359
rect 39681 12325 39715 12359
rect 41521 12325 41555 12359
rect 2053 12257 2087 12291
rect 4997 12257 5031 12291
rect 5641 12257 5675 12291
rect 6193 12257 6227 12291
rect 6745 12257 6779 12291
rect 9413 12257 9447 12291
rect 9689 12257 9723 12291
rect 12265 12257 12299 12291
rect 13461 12257 13495 12291
rect 20361 12257 20395 12291
rect 22661 12257 22695 12291
rect 22845 12257 22879 12291
rect 24961 12257 24995 12291
rect 25145 12257 25179 12291
rect 27353 12257 27387 12291
rect 29101 12257 29135 12291
rect 30297 12257 30331 12291
rect 32873 12257 32907 12291
rect 33701 12257 33735 12291
rect 33885 12257 33919 12291
rect 34161 12257 34195 12291
rect 35357 12257 35391 12291
rect 35541 12257 35575 12291
rect 38117 12257 38151 12291
rect 38945 12257 38979 12291
rect 39865 12257 39899 12291
rect 40509 12257 40543 12291
rect 1961 12189 1995 12223
rect 3157 12189 3191 12223
rect 3525 12189 3559 12223
rect 3985 12189 4019 12223
rect 4169 12189 4203 12223
rect 5273 12189 5307 12223
rect 5917 12189 5951 12223
rect 6101 12189 6135 12223
rect 6377 12189 6411 12223
rect 6929 12189 6963 12223
rect 7389 12189 7423 12223
rect 7573 12189 7607 12223
rect 7665 12189 7699 12223
rect 7849 12189 7883 12223
rect 11897 12189 11931 12223
rect 11989 12189 12023 12223
rect 12081 12189 12115 12223
rect 12541 12189 12575 12223
rect 12633 12189 12667 12223
rect 13553 12189 13587 12223
rect 14289 12189 14323 12223
rect 14381 12189 14415 12223
rect 14749 12189 14783 12223
rect 16405 12189 16439 12223
rect 16681 12189 16715 12223
rect 16865 12189 16899 12223
rect 17601 12189 17635 12223
rect 17693 12189 17727 12223
rect 17877 12189 17911 12223
rect 19349 12189 19383 12223
rect 20269 12189 20303 12223
rect 22109 12189 22143 12223
rect 23581 12189 23615 12223
rect 26065 12189 26099 12223
rect 26617 12189 26651 12223
rect 29193 12189 29227 12223
rect 29745 12189 29779 12223
rect 30481 12189 30515 12223
rect 32597 12189 32631 12223
rect 32965 12189 32999 12223
rect 33609 12189 33643 12223
rect 34345 12189 34379 12223
rect 36369 12189 36403 12223
rect 37197 12189 37231 12223
rect 38393 12189 38427 12223
rect 39175 12189 39209 12223
rect 39401 12189 39435 12223
rect 39497 12189 39531 12223
rect 40141 12189 40175 12223
rect 40233 12189 40267 12223
rect 40325 12189 40359 12223
rect 41153 12189 41187 12223
rect 41337 12189 41371 12223
rect 41521 12189 41555 12223
rect 2421 12121 2455 12155
rect 5549 12121 5583 12155
rect 6653 12121 6687 12155
rect 7757 12121 7791 12155
rect 11405 12121 11439 12155
rect 11621 12121 11655 12155
rect 12817 12121 12851 12155
rect 14657 12121 14691 12155
rect 16957 12121 16991 12155
rect 21833 12121 21867 12155
rect 23857 12121 23891 12155
rect 27629 12121 27663 12155
rect 30113 12121 30147 12155
rect 32321 12121 32355 12155
rect 32689 12121 32723 12155
rect 34069 12121 34103 12155
rect 37381 12121 37415 12155
rect 39313 12121 39347 12155
rect 40003 12121 40037 12155
rect 3341 12053 3375 12087
rect 4721 12053 4755 12087
rect 5825 12053 5859 12087
rect 6561 12053 6595 12087
rect 7113 12053 7147 12087
rect 7481 12053 7515 12087
rect 11713 12053 11747 12087
rect 16221 12053 16255 12087
rect 19993 12053 20027 12087
rect 22569 12053 22603 12087
rect 23029 12053 23063 12087
rect 24501 12053 24535 12087
rect 24869 12053 24903 12087
rect 25513 12053 25547 12087
rect 30849 12053 30883 12087
rect 33149 12053 33183 12087
rect 33241 12053 33275 12087
rect 34897 12053 34931 12087
rect 35265 12053 35299 12087
rect 35817 12053 35851 12087
rect 36553 12053 36587 12087
rect 40601 12053 40635 12087
rect 3249 11849 3283 11883
rect 4369 11849 4403 11883
rect 4813 11849 4847 11883
rect 6929 11849 6963 11883
rect 7481 11849 7515 11883
rect 12173 11849 12207 11883
rect 12817 11849 12851 11883
rect 12909 11849 12943 11883
rect 19165 11849 19199 11883
rect 19625 11849 19659 11883
rect 26801 11849 26835 11883
rect 29653 11849 29687 11883
rect 30481 11849 30515 11883
rect 36277 11849 36311 11883
rect 36737 11849 36771 11883
rect 36829 11849 36863 11883
rect 40693 11849 40727 11883
rect 4169 11781 4203 11815
rect 4629 11781 4663 11815
rect 6653 11781 6687 11815
rect 7389 11781 7423 11815
rect 7941 11781 7975 11815
rect 8585 11781 8619 11815
rect 8677 11781 8711 11815
rect 9045 11781 9079 11815
rect 13829 11781 13863 11815
rect 16497 11781 16531 11815
rect 16957 11781 16991 11815
rect 21097 11781 21131 11815
rect 24501 11781 24535 11815
rect 27445 11781 27479 11815
rect 28181 11781 28215 11815
rect 31677 11781 31711 11815
rect 31861 11781 31895 11815
rect 32965 11781 32999 11815
rect 34805 11781 34839 11815
rect 39221 11781 39255 11815
rect 3525 11713 3559 11747
rect 4905 11713 4939 11747
rect 5917 11713 5951 11747
rect 6101 11713 6135 11747
rect 6469 11713 6503 11747
rect 7113 11713 7147 11747
rect 7665 11713 7699 11747
rect 8125 11713 8159 11747
rect 8309 11713 8343 11747
rect 8401 11713 8435 11747
rect 8769 11713 8803 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 10425 11713 10459 11747
rect 11989 11713 12023 11747
rect 12265 11713 12299 11747
rect 12357 11713 12391 11747
rect 12633 11713 12667 11747
rect 13093 11713 13127 11747
rect 13553 11713 13587 11747
rect 13645 11713 13679 11747
rect 14565 11713 14599 11747
rect 16129 11713 16163 11747
rect 16313 11713 16347 11747
rect 19533 11713 19567 11747
rect 20361 11713 20395 11747
rect 21373 11713 21407 11747
rect 22385 11713 22419 11747
rect 24225 11713 24259 11747
rect 26433 11713 26467 11747
rect 27169 11713 27203 11747
rect 27537 11713 27571 11747
rect 27721 11713 27755 11747
rect 27905 11713 27939 11747
rect 30389 11713 30423 11747
rect 30941 11713 30975 11747
rect 32689 11713 32723 11747
rect 34529 11713 34563 11747
rect 1501 11645 1535 11679
rect 1777 11645 1811 11679
rect 5733 11645 5767 11679
rect 7297 11645 7331 11679
rect 7757 11645 7791 11679
rect 9689 11645 9723 11679
rect 12449 11645 12483 11679
rect 13277 11645 13311 11679
rect 14105 11645 14139 11679
rect 14473 11645 14507 11679
rect 16681 11645 16715 11679
rect 19717 11645 19751 11679
rect 20913 11645 20947 11679
rect 21281 11645 21315 11679
rect 22661 11645 22695 11679
rect 26525 11645 26559 11679
rect 27261 11645 27295 11679
rect 30665 11645 30699 11679
rect 31585 11645 31619 11679
rect 37013 11645 37047 11679
rect 38945 11645 38979 11679
rect 4629 11577 4663 11611
rect 8309 11577 8343 11611
rect 10333 11577 10367 11611
rect 11989 11577 12023 11611
rect 18429 11577 18463 11611
rect 26985 11577 27019 11611
rect 34437 11577 34471 11611
rect 36369 11577 36403 11611
rect 4353 11509 4387 11543
rect 4537 11509 4571 11543
rect 6837 11509 6871 11543
rect 7389 11509 7423 11543
rect 7665 11509 7699 11543
rect 8953 11509 8987 11543
rect 10149 11509 10183 11543
rect 12633 11509 12667 11543
rect 13829 11509 13863 11543
rect 14749 11509 14783 11543
rect 21097 11509 21131 11543
rect 21557 11509 21591 11543
rect 24133 11509 24167 11543
rect 25973 11509 26007 11543
rect 26433 11509 26467 11543
rect 27169 11509 27203 11543
rect 30021 11509 30055 11543
rect 3341 11305 3375 11339
rect 9210 11305 9244 11339
rect 11713 11305 11747 11339
rect 12541 11305 12575 11339
rect 13277 11305 13311 11339
rect 13461 11305 13495 11339
rect 13737 11305 13771 11339
rect 13921 11305 13955 11339
rect 14933 11305 14967 11339
rect 17555 11305 17589 11339
rect 22569 11305 22603 11339
rect 31493 11305 31527 11339
rect 35541 11305 35575 11339
rect 37565 11305 37599 11339
rect 8217 11237 8251 11271
rect 10701 11237 10735 11271
rect 12909 11237 12943 11271
rect 31309 11237 31343 11271
rect 1593 11169 1627 11203
rect 3801 11169 3835 11203
rect 8953 11169 8987 11203
rect 11621 11169 11655 11203
rect 12357 11169 12391 11203
rect 13645 11169 13679 11203
rect 14289 11169 14323 11203
rect 15761 11169 15795 11203
rect 18797 11169 18831 11203
rect 18889 11169 18923 11203
rect 19533 11169 19567 11203
rect 21005 11169 21039 11203
rect 23213 11169 23247 11203
rect 24133 11169 24167 11203
rect 24961 11169 24995 11203
rect 26709 11169 26743 11203
rect 27353 11169 27387 11203
rect 29561 11169 29595 11203
rect 35633 11169 35667 11203
rect 35817 11169 35851 11203
rect 36093 11169 36127 11203
rect 3433 11101 3467 11135
rect 3617 11101 3651 11135
rect 6745 11101 6779 11135
rect 8401 11101 8435 11135
rect 8493 11101 8527 11135
rect 8585 11101 8619 11135
rect 8677 11101 8711 11135
rect 11989 11101 12023 11135
rect 12633 11101 12667 11135
rect 12731 11101 12765 11135
rect 12909 11101 12943 11135
rect 13553 11101 13587 11135
rect 16129 11101 16163 11135
rect 19257 11101 19291 11135
rect 22017 11101 22051 11135
rect 22109 11101 22143 11135
rect 22385 11101 22419 11135
rect 23029 11101 23063 11135
rect 28273 11101 28307 11135
rect 32505 11101 32539 11135
rect 34805 11101 34839 11135
rect 34897 11101 34931 11135
rect 35357 11101 35391 11135
rect 35449 11101 35483 11135
rect 37657 11101 37691 11135
rect 37841 11101 37875 11135
rect 38025 11101 38059 11135
rect 1869 11033 1903 11067
rect 3525 11033 3559 11067
rect 4077 11033 4111 11067
rect 13093 11033 13127 11067
rect 18705 11033 18739 11067
rect 22201 11033 22235 11067
rect 22937 11033 22971 11067
rect 23581 11033 23615 11067
rect 25237 11033 25271 11067
rect 29837 11033 29871 11067
rect 31769 11033 31803 11067
rect 37749 11033 37783 11067
rect 5549 10965 5583 10999
rect 6561 10965 6595 10999
rect 11805 10965 11839 10999
rect 11897 10965 11931 10999
rect 12081 10965 12115 10999
rect 13293 10965 13327 10999
rect 18337 10965 18371 10999
rect 21833 10965 21867 10999
rect 26801 10965 26835 10999
rect 27721 10965 27755 10999
rect 31953 10965 31987 10999
rect 38209 10965 38243 10999
rect 1501 10761 1535 10795
rect 2513 10761 2547 10795
rect 4537 10761 4571 10795
rect 4705 10761 4739 10795
rect 8309 10761 8343 10795
rect 8493 10761 8527 10795
rect 9137 10761 9171 10795
rect 14013 10761 14047 10795
rect 20177 10761 20211 10795
rect 22937 10761 22971 10795
rect 25513 10761 25547 10795
rect 25973 10761 26007 10795
rect 27353 10761 27387 10795
rect 28733 10761 28767 10795
rect 32137 10761 32171 10795
rect 32597 10761 32631 10795
rect 35357 10761 35391 10795
rect 40601 10761 40635 10795
rect 4905 10693 4939 10727
rect 13553 10693 13587 10727
rect 13645 10693 13679 10727
rect 15485 10693 15519 10727
rect 18613 10693 18647 10727
rect 23673 10693 23707 10727
rect 25881 10693 25915 10727
rect 27445 10693 27479 10727
rect 34529 10693 34563 10727
rect 35725 10693 35759 10727
rect 36185 10693 36219 10727
rect 1685 10625 1719 10659
rect 2421 10625 2455 10659
rect 2605 10625 2639 10659
rect 2789 10625 2823 10659
rect 2881 10625 2915 10659
rect 3065 10625 3099 10659
rect 3249 10625 3283 10659
rect 3985 10625 4019 10659
rect 4169 10625 4203 10659
rect 4261 10625 4295 10659
rect 5733 10625 5767 10659
rect 5825 10625 5859 10659
rect 6377 10625 6411 10659
rect 6561 10625 6595 10659
rect 7389 10625 7423 10659
rect 7941 10625 7975 10659
rect 8125 10625 8159 10659
rect 8677 10625 8711 10659
rect 9045 10625 9079 10659
rect 9689 10625 9723 10659
rect 11529 10625 11563 10659
rect 13369 10625 13403 10659
rect 13737 10625 13771 10659
rect 15761 10625 15795 10659
rect 23949 10625 23983 10659
rect 24041 10625 24075 10659
rect 24133 10625 24167 10659
rect 24317 10625 24351 10659
rect 26709 10625 26743 10659
rect 28825 10625 28859 10659
rect 29377 10625 29411 10659
rect 32505 10625 32539 10659
rect 32965 10625 32999 10659
rect 34253 10625 34287 10659
rect 35536 10625 35570 10659
rect 35633 10625 35667 10659
rect 35908 10625 35942 10659
rect 36001 10625 36035 10659
rect 36093 10625 36127 10659
rect 36277 10625 36311 10659
rect 37657 10625 37691 10659
rect 37933 10625 37967 10659
rect 40509 10625 40543 10659
rect 40785 10625 40819 10659
rect 3893 10557 3927 10591
rect 5917 10557 5951 10591
rect 6009 10557 6043 10591
rect 7481 10557 7515 10591
rect 7849 10557 7883 10591
rect 8585 10557 8619 10591
rect 9413 10557 9447 10591
rect 11805 10557 11839 10591
rect 18337 10557 18371 10591
rect 20729 10557 20763 10591
rect 22293 10557 22327 10591
rect 23029 10557 23063 10591
rect 26065 10557 26099 10591
rect 27537 10557 27571 10591
rect 28549 10557 28583 10591
rect 29929 10557 29963 10591
rect 32781 10557 32815 10591
rect 33517 10557 33551 10591
rect 34529 10557 34563 10591
rect 37749 10557 37783 10591
rect 38209 10557 38243 10591
rect 39681 10557 39715 10591
rect 40325 10557 40359 10591
rect 5549 10489 5583 10523
rect 3065 10421 3099 10455
rect 4169 10421 4203 10455
rect 4445 10421 4479 10455
rect 4721 10421 4755 10455
rect 6469 10421 6503 10455
rect 7389 10421 7423 10455
rect 7757 10421 7791 10455
rect 9597 10421 9631 10455
rect 13277 10421 13311 10455
rect 13921 10421 13955 10455
rect 20085 10421 20119 10455
rect 23765 10421 23799 10455
rect 26433 10421 26467 10455
rect 26985 10421 27019 10455
rect 29193 10421 29227 10455
rect 34345 10421 34379 10455
rect 37473 10421 37507 10455
rect 39773 10421 39807 10455
rect 3341 10217 3375 10251
rect 5549 10217 5583 10251
rect 7021 10217 7055 10251
rect 11621 10217 11655 10251
rect 13369 10217 13403 10251
rect 14105 10217 14139 10251
rect 22201 10217 22235 10251
rect 23305 10217 23339 10251
rect 25697 10217 25731 10251
rect 28917 10217 28951 10251
rect 33149 10217 33183 10251
rect 36829 10217 36863 10251
rect 38577 10217 38611 10251
rect 27997 10149 28031 10183
rect 28825 10149 28859 10183
rect 30849 10149 30883 10183
rect 31033 10149 31067 10183
rect 34713 10149 34747 10183
rect 37841 10149 37875 10183
rect 11805 10081 11839 10115
rect 12265 10081 12299 10115
rect 13277 10081 13311 10115
rect 13645 10081 13679 10115
rect 15577 10081 15611 10115
rect 20729 10081 20763 10115
rect 22753 10081 22787 10115
rect 25329 10081 25363 10115
rect 26249 10081 26283 10115
rect 26525 10081 26559 10115
rect 30113 10081 30147 10115
rect 31217 10081 31251 10115
rect 31401 10081 31435 10115
rect 33241 10081 33275 10115
rect 34529 10081 34563 10115
rect 35173 10081 35207 10115
rect 35357 10081 35391 10115
rect 36369 10081 36403 10115
rect 37933 10081 37967 10115
rect 3157 10013 3191 10047
rect 3341 10013 3375 10047
rect 5365 10013 5399 10047
rect 5549 10013 5583 10047
rect 5641 10013 5675 10047
rect 5825 10013 5859 10047
rect 6009 10013 6043 10047
rect 6101 10013 6135 10047
rect 6193 10013 6227 10047
rect 6285 10013 6319 10047
rect 6561 10013 6595 10047
rect 6837 10013 6871 10047
rect 7113 10013 7147 10047
rect 7297 10013 7331 10047
rect 11897 10013 11931 10047
rect 12633 10013 12667 10047
rect 13737 10013 13771 10047
rect 15853 10013 15887 10047
rect 20453 10013 20487 10047
rect 22477 10013 22511 10047
rect 22661 10013 22695 10047
rect 22845 10013 22879 10047
rect 23029 10013 23063 10047
rect 23305 10013 23339 10047
rect 23489 10013 23523 10047
rect 23581 10013 23615 10047
rect 23674 10013 23708 10047
rect 23857 10013 23891 10047
rect 23949 10013 23983 10047
rect 24046 10013 24080 10047
rect 24961 10013 24995 10047
rect 25145 10013 25179 10047
rect 25237 10013 25271 10047
rect 25513 10013 25547 10047
rect 28089 10015 28123 10049
rect 28273 10013 28307 10047
rect 28365 10013 28399 10047
rect 28457 10013 28491 10047
rect 28641 10013 28675 10047
rect 30297 10013 30331 10047
rect 30573 10013 30607 10047
rect 30665 10013 30699 10047
rect 30941 10013 30975 10047
rect 33425 10013 33459 10047
rect 33517 10013 33551 10047
rect 33614 10023 33648 10057
rect 36093 10013 36127 10047
rect 36277 10013 36311 10047
rect 36553 10013 36587 10047
rect 36645 10013 36679 10047
rect 37289 10013 37323 10047
rect 37565 10013 37599 10047
rect 37657 10013 37691 10047
rect 38853 10013 38887 10047
rect 38945 10013 38979 10047
rect 39221 10013 39255 10047
rect 39865 10013 39899 10047
rect 40417 10013 40451 10047
rect 5733 9945 5767 9979
rect 23213 9945 23247 9979
rect 29101 9945 29135 9979
rect 29285 9945 29319 9979
rect 30481 9945 30515 9979
rect 31677 9945 31711 9979
rect 33287 9945 33321 9979
rect 35081 9945 35115 9979
rect 35541 9945 35575 9979
rect 37473 9945 37507 9979
rect 39037 9945 39071 9979
rect 40693 9945 40727 9979
rect 6469 9877 6503 9911
rect 6653 9877 6687 9911
rect 7205 9877 7239 9911
rect 24225 9877 24259 9911
rect 29561 9877 29595 9911
rect 31217 9877 31251 9911
rect 33885 9877 33919 9911
rect 38669 9877 38703 9911
rect 40785 9877 40819 9911
rect 6653 9673 6687 9707
rect 8217 9673 8251 9707
rect 31217 9673 31251 9707
rect 38301 9673 38335 9707
rect 3065 9605 3099 9639
rect 8401 9605 8435 9639
rect 20545 9605 20579 9639
rect 23305 9605 23339 9639
rect 27261 9605 27295 9639
rect 27353 9605 27387 9639
rect 29469 9605 29503 9639
rect 32137 9605 32171 9639
rect 33885 9605 33919 9639
rect 35449 9605 35483 9639
rect 36185 9605 36219 9639
rect 36461 9605 36495 9639
rect 38945 9605 38979 9639
rect 2513 9537 2547 9571
rect 2697 9537 2731 9571
rect 2973 9537 3007 9571
rect 3157 9537 3191 9571
rect 5273 9537 5307 9571
rect 5457 9537 5491 9571
rect 5549 9537 5583 9571
rect 6009 9537 6043 9571
rect 6650 9537 6684 9571
rect 7297 9537 7331 9571
rect 8309 9537 8343 9571
rect 10057 9537 10091 9571
rect 10425 9537 10459 9571
rect 11253 9537 11287 9571
rect 11621 9537 11655 9571
rect 18429 9537 18463 9571
rect 19441 9537 19475 9571
rect 19579 9537 19613 9571
rect 19717 9537 19751 9571
rect 19809 9537 19843 9571
rect 19901 9537 19935 9571
rect 20177 9537 20211 9571
rect 20361 9537 20395 9571
rect 21465 9537 21499 9571
rect 21649 9537 21683 9571
rect 26709 9537 26743 9571
rect 27169 9537 27203 9571
rect 27537 9537 27571 9571
rect 29745 9537 29779 9571
rect 30665 9537 30699 9571
rect 30941 9537 30975 9571
rect 31033 9537 31067 9571
rect 31861 9537 31895 9571
rect 35633 9537 35667 9571
rect 36369 9537 36403 9571
rect 36558 9537 36592 9571
rect 37749 9537 37783 9571
rect 38209 9537 38243 9571
rect 5825 9469 5859 9503
rect 7113 9469 7147 9503
rect 7389 9469 7423 9503
rect 7481 9469 7515 9503
rect 7573 9469 7607 9503
rect 7757 9469 7791 9503
rect 10333 9469 10367 9503
rect 20085 9469 20119 9503
rect 23581 9469 23615 9503
rect 23857 9469 23891 9503
rect 24133 9469 24167 9503
rect 25605 9469 25639 9503
rect 26249 9469 26283 9503
rect 32965 9469 32999 9503
rect 33609 9469 33643 9503
rect 35357 9469 35391 9503
rect 35817 9469 35851 9503
rect 37841 9469 37875 9503
rect 38117 9469 38151 9503
rect 38669 9469 38703 9503
rect 40417 9469 40451 9503
rect 7021 9401 7055 9435
rect 8585 9401 8619 9435
rect 21281 9401 21315 9435
rect 26525 9401 26559 9435
rect 26985 9401 27019 9435
rect 36185 9401 36219 9435
rect 2513 9333 2547 9367
rect 5273 9333 5307 9367
rect 5825 9333 5859 9367
rect 6193 9333 6227 9367
rect 6469 9333 6503 9367
rect 8033 9333 8067 9367
rect 10149 9333 10183 9367
rect 10241 9333 10275 9367
rect 21649 9333 21683 9367
rect 21833 9333 21867 9367
rect 25697 9333 25731 9367
rect 27997 9333 28031 9367
rect 30757 9333 30791 9367
rect 4537 9129 4571 9163
rect 6469 9129 6503 9163
rect 6653 9129 6687 9163
rect 9045 9129 9079 9163
rect 9768 9129 9802 9163
rect 12173 9129 12207 9163
rect 17588 9129 17622 9163
rect 19257 9129 19291 9163
rect 21741 9129 21775 9163
rect 21925 9129 21959 9163
rect 22569 9129 22603 9163
rect 22753 9129 22787 9163
rect 24593 9129 24627 9163
rect 32229 9129 32263 9163
rect 32781 9129 32815 9163
rect 38577 9129 38611 9163
rect 5273 9061 5307 9095
rect 19993 9061 20027 9095
rect 22293 9061 22327 9095
rect 37657 9061 37691 9095
rect 1409 8993 1443 9027
rect 3157 8993 3191 9027
rect 3617 8993 3651 9027
rect 4629 8993 4663 9027
rect 5549 8993 5583 9027
rect 5917 8993 5951 9027
rect 6009 8993 6043 9027
rect 6837 8993 6871 9027
rect 7297 8993 7331 9027
rect 9505 8993 9539 9027
rect 12725 8993 12759 9027
rect 13001 8993 13035 9027
rect 17325 8993 17359 9027
rect 19441 8993 19475 9027
rect 20453 8993 20487 9027
rect 21833 8993 21867 9027
rect 25145 8993 25179 9027
rect 25237 8993 25271 9027
rect 27077 8993 27111 9027
rect 29745 8993 29779 9027
rect 32137 8993 32171 9027
rect 36645 8993 36679 9027
rect 37749 8993 37783 9027
rect 3433 8925 3467 8959
rect 4445 8925 4479 8959
rect 4813 8925 4847 8959
rect 5273 8925 5307 8959
rect 5457 8925 5491 8959
rect 6285 8925 6319 8959
rect 6469 8925 6503 8959
rect 6929 8925 6963 8959
rect 8217 8925 8251 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 11345 8925 11379 8959
rect 11989 8925 12023 8959
rect 12081 8925 12115 8959
rect 12265 8925 12299 8959
rect 13093 8925 13127 8959
rect 19533 8925 19567 8959
rect 20361 8925 20395 8959
rect 21465 8925 21499 8959
rect 22109 8925 22143 8959
rect 24777 8925 24811 8959
rect 24869 8925 24903 8959
rect 29837 8925 29871 8959
rect 32656 8925 32690 8959
rect 32873 8925 32907 8959
rect 33265 8925 33299 8959
rect 36185 8925 36219 8959
rect 36277 8925 36311 8959
rect 37105 8925 37139 8959
rect 37289 8925 37323 8959
rect 37473 8925 37507 8959
rect 38485 8925 38519 8959
rect 38669 8925 38703 8959
rect 1685 8857 1719 8891
rect 3249 8857 3283 8891
rect 4537 8857 4571 8891
rect 6193 8857 6227 8891
rect 19809 8857 19843 8891
rect 19901 8857 19935 8891
rect 21557 8857 21591 8891
rect 21741 8857 21775 8891
rect 22385 8857 22419 8891
rect 22601 8857 22635 8891
rect 26801 8857 26835 8891
rect 30113 8857 30147 8891
rect 30205 8857 30239 8891
rect 33057 8857 33091 8891
rect 33149 8857 33183 8891
rect 36553 8857 36587 8891
rect 37381 8857 37415 8891
rect 3801 8789 3835 8823
rect 4997 8789 5031 8823
rect 8769 8789 8803 8823
rect 11253 8789 11287 8823
rect 19073 8789 19107 8823
rect 25329 8789 25363 8823
rect 29561 8789 29595 8823
rect 32597 8789 32631 8823
rect 33425 8789 33459 8823
rect 36001 8789 36035 8823
rect 38393 8789 38427 8823
rect 6193 8585 6227 8619
rect 6377 8585 6411 8619
rect 10793 8585 10827 8619
rect 10885 8585 10919 8619
rect 11805 8585 11839 8619
rect 13553 8585 13587 8619
rect 21097 8585 21131 8619
rect 22293 8585 22327 8619
rect 22385 8585 22419 8619
rect 22477 8585 22511 8619
rect 23305 8585 23339 8619
rect 26433 8585 26467 8619
rect 27353 8585 27387 8619
rect 37105 8585 37139 8619
rect 9597 8517 9631 8551
rect 11345 8517 11379 8551
rect 11713 8517 11747 8551
rect 13001 8517 13035 8551
rect 18153 8517 18187 8551
rect 22109 8517 22143 8551
rect 29745 8517 29779 8551
rect 34253 8517 34287 8551
rect 38853 8517 38887 8551
rect 1777 8449 1811 8483
rect 2973 8449 3007 8483
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 6929 8449 6963 8483
rect 9229 8449 9263 8483
rect 9505 8449 9539 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 10149 8449 10183 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 11069 8449 11103 8483
rect 11161 8449 11195 8483
rect 11897 8449 11931 8483
rect 12449 8449 12483 8483
rect 12541 8449 12575 8483
rect 12817 8449 12851 8483
rect 13093 8449 13127 8483
rect 13185 8449 13219 8483
rect 22937 8449 22971 8483
rect 25145 8449 25179 8483
rect 25329 8449 25363 8483
rect 25421 8449 25455 8483
rect 25513 8449 25547 8483
rect 26985 8449 27019 8483
rect 27169 8449 27203 8483
rect 30021 8449 30055 8483
rect 32137 8449 32171 8483
rect 36001 8449 36035 8483
rect 36185 8449 36219 8483
rect 36737 8449 36771 8483
rect 36921 8449 36955 8483
rect 39129 8449 39163 8483
rect 1869 8381 1903 8415
rect 2881 8381 2915 8415
rect 3249 8381 3283 8415
rect 5917 8381 5951 8415
rect 8953 8381 8987 8415
rect 9965 8381 9999 8415
rect 12081 8381 12115 8415
rect 12265 8381 12299 8415
rect 12357 8381 12391 8415
rect 15025 8381 15059 8415
rect 15301 8381 15335 8415
rect 18889 8381 18923 8415
rect 19349 8381 19383 8415
rect 19625 8381 19659 8415
rect 22845 8381 22879 8415
rect 25789 8381 25823 8415
rect 28273 8381 28307 8415
rect 30665 8381 30699 8415
rect 32413 8381 32447 8415
rect 33977 8381 34011 8415
rect 35725 8381 35759 8415
rect 39221 8381 39255 8415
rect 39773 8381 39807 8415
rect 2145 8313 2179 8347
rect 7481 8313 7515 8347
rect 9321 8313 9355 8347
rect 10333 8313 10367 8347
rect 11529 8313 11563 8347
rect 13369 8313 13403 8347
rect 22661 8313 22695 8347
rect 25697 8313 25731 8347
rect 37381 8313 37415 8347
rect 2237 8245 2271 8279
rect 4721 8245 4755 8279
rect 6009 8245 6043 8279
rect 6561 8245 6595 8279
rect 11253 8245 11287 8279
rect 12725 8245 12759 8279
rect 30113 8245 30147 8279
rect 33885 8245 33919 8279
rect 36001 8245 36035 8279
rect 3157 8041 3191 8075
rect 3433 8041 3467 8075
rect 4077 8041 4111 8075
rect 8585 8041 8619 8075
rect 8769 8041 8803 8075
rect 9505 8041 9539 8075
rect 10333 8041 10367 8075
rect 19073 8041 19107 8075
rect 19901 8041 19935 8075
rect 25421 8041 25455 8075
rect 26985 8041 27019 8075
rect 29377 8041 29411 8075
rect 32137 8041 32171 8075
rect 33333 8041 33367 8075
rect 38761 8041 38795 8075
rect 9229 7973 9263 8007
rect 25605 7973 25639 8007
rect 32045 7973 32079 8007
rect 37381 7973 37415 8007
rect 10609 7905 10643 7939
rect 11161 7905 11195 7939
rect 11345 7905 11379 7939
rect 13829 7905 13863 7939
rect 19257 7905 19291 7939
rect 24501 7905 24535 7939
rect 29101 7905 29135 7939
rect 31585 7905 31619 7939
rect 32689 7905 32723 7939
rect 33885 7905 33919 7939
rect 35633 7905 35667 7939
rect 1409 7837 1443 7871
rect 3801 7837 3835 7871
rect 4169 7837 4203 7871
rect 8953 7837 8987 7871
rect 9045 7837 9079 7871
rect 9321 7837 9355 7871
rect 9505 7837 9539 7871
rect 10333 7837 10367 7871
rect 10517 7837 10551 7871
rect 11069 7837 11103 7871
rect 11437 7837 11471 7871
rect 11713 7837 11747 7871
rect 11805 7837 11839 7871
rect 18521 7837 18555 7871
rect 18889 7837 18923 7871
rect 19993 7837 20027 7871
rect 20269 7837 20303 7871
rect 20361 7837 20395 7871
rect 20913 7837 20947 7871
rect 24593 7837 24627 7871
rect 25697 7837 25731 7871
rect 26709 7837 26743 7871
rect 26801 7837 26835 7871
rect 26985 7837 27019 7871
rect 27077 7837 27111 7871
rect 27261 7837 27295 7871
rect 29009 7837 29043 7871
rect 31309 7837 31343 7871
rect 31677 7837 31711 7871
rect 32321 7837 32355 7871
rect 32413 7837 32447 7871
rect 38393 7837 38427 7871
rect 38669 7837 38703 7871
rect 38853 7837 38887 7871
rect 1685 7769 1719 7803
rect 3401 7769 3435 7803
rect 3617 7769 3651 7803
rect 8401 7769 8435 7803
rect 8601 7769 8635 7803
rect 9229 7769 9263 7803
rect 10977 7769 11011 7803
rect 13553 7769 13587 7803
rect 18705 7769 18739 7803
rect 18797 7769 18831 7803
rect 20177 7769 20211 7803
rect 25237 7769 25271 7803
rect 26433 7769 26467 7803
rect 31033 7769 31067 7803
rect 32781 7769 32815 7803
rect 35909 7769 35943 7803
rect 3249 7701 3283 7735
rect 3893 7701 3927 7735
rect 3985 7701 4019 7735
rect 10885 7701 10919 7735
rect 11621 7701 11655 7735
rect 12081 7701 12115 7735
rect 20545 7701 20579 7735
rect 20729 7701 20763 7735
rect 24961 7701 24995 7735
rect 25437 7701 25471 7735
rect 27169 7701 27203 7735
rect 29561 7701 29595 7735
rect 1777 7497 1811 7531
rect 11529 7497 11563 7531
rect 12449 7497 12483 7531
rect 13001 7497 13035 7531
rect 28549 7497 28583 7531
rect 30665 7497 30699 7531
rect 32505 7497 32539 7531
rect 34453 7497 34487 7531
rect 34713 7497 34747 7531
rect 35817 7497 35851 7531
rect 2237 7429 2271 7463
rect 12633 7429 12667 7463
rect 19717 7429 19751 7463
rect 20729 7429 20763 7463
rect 21281 7429 21315 7463
rect 24317 7429 24351 7463
rect 24409 7429 24443 7463
rect 28181 7429 28215 7463
rect 30849 7429 30883 7463
rect 34253 7429 34287 7463
rect 35265 7429 35299 7463
rect 36001 7429 36035 7463
rect 36185 7429 36219 7463
rect 37473 7429 37507 7463
rect 38209 7429 38243 7463
rect 38669 7429 38703 7463
rect 1685 7361 1719 7395
rect 1869 7361 1903 7395
rect 1961 7361 1995 7395
rect 2053 7361 2087 7395
rect 11713 7361 11747 7395
rect 12357 7361 12391 7395
rect 12725 7361 12759 7395
rect 12817 7361 12851 7395
rect 13093 7361 13127 7395
rect 13277 7361 13311 7395
rect 19257 7361 19291 7395
rect 19349 7361 19383 7395
rect 24133 7361 24167 7395
rect 24501 7361 24535 7395
rect 25513 7361 25547 7395
rect 26249 7361 26283 7395
rect 27261 7361 27295 7395
rect 27537 7361 27571 7395
rect 27905 7361 27939 7395
rect 28089 7361 28123 7395
rect 28365 7361 28399 7395
rect 29377 7361 29411 7395
rect 29561 7361 29595 7395
rect 29653 7361 29687 7395
rect 29745 7361 29779 7395
rect 30757 7361 30791 7395
rect 30941 7361 30975 7395
rect 31125 7361 31159 7395
rect 32137 7361 32171 7395
rect 32230 7361 32264 7395
rect 33885 7361 33919 7395
rect 33977 7361 34011 7395
rect 34161 7361 34195 7395
rect 34897 7361 34931 7395
rect 34989 7361 35023 7395
rect 35357 7361 35391 7395
rect 35449 7361 35483 7395
rect 35633 7361 35667 7395
rect 36461 7361 36495 7395
rect 36645 7361 36679 7395
rect 36737 7361 36771 7395
rect 36829 7361 36863 7395
rect 38485 7361 38519 7395
rect 38761 7361 38795 7395
rect 11897 7293 11931 7327
rect 13001 7293 13035 7327
rect 13185 7293 13219 7327
rect 19625 7293 19659 7327
rect 20177 7293 20211 7327
rect 23305 7293 23339 7327
rect 23581 7293 23615 7327
rect 24777 7293 24811 7327
rect 26065 7293 26099 7327
rect 27169 7293 27203 7327
rect 27629 7293 27663 7327
rect 27721 7293 27755 7327
rect 29285 7293 29319 7327
rect 30021 7293 30055 7327
rect 31217 7293 31251 7327
rect 31309 7293 31343 7327
rect 31401 7293 31435 7327
rect 31585 7293 31619 7327
rect 38301 7293 38335 7327
rect 2237 7225 2271 7259
rect 12633 7225 12667 7259
rect 21005 7225 21039 7259
rect 24685 7225 24719 7259
rect 28641 7225 28675 7259
rect 29929 7225 29963 7259
rect 34161 7225 34195 7259
rect 38945 7225 38979 7259
rect 19073 7157 19107 7191
rect 21833 7157 21867 7191
rect 25421 7157 25455 7191
rect 26985 7157 27019 7191
rect 34437 7157 34471 7191
rect 34621 7157 34655 7191
rect 36369 7157 36403 7191
rect 37013 7157 37047 7191
rect 6653 6953 6687 6987
rect 8585 6953 8619 6987
rect 8769 6953 8803 6987
rect 8953 6953 8987 6987
rect 10412 6953 10446 6987
rect 11897 6953 11931 6987
rect 19625 6953 19659 6987
rect 21109 6953 21143 6987
rect 24409 6953 24443 6987
rect 25893 6953 25927 6987
rect 26512 6953 26546 6987
rect 28917 6953 28951 6987
rect 29561 6953 29595 6987
rect 33044 6953 33078 6987
rect 36461 6953 36495 6987
rect 37197 6953 37231 6987
rect 7113 6885 7147 6919
rect 7849 6885 7883 6919
rect 31033 6885 31067 6919
rect 31585 6885 31619 6919
rect 3525 6817 3559 6851
rect 5273 6817 5307 6851
rect 6837 6817 6871 6851
rect 7665 6817 7699 6851
rect 8217 6817 8251 6851
rect 9045 6817 9079 6851
rect 10149 6817 10183 6851
rect 21373 6817 21407 6851
rect 21465 6817 21499 6851
rect 26157 6817 26191 6851
rect 26249 6817 26283 6851
rect 30481 6817 30515 6851
rect 32781 6817 32815 6851
rect 34529 6817 34563 6851
rect 34897 6817 34931 6851
rect 35909 6817 35943 6851
rect 36277 6817 36311 6851
rect 2605 6749 2639 6783
rect 2789 6749 2823 6783
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 3341 6749 3375 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 4629 6749 4663 6783
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 6469 6749 6503 6783
rect 6653 6749 6687 6783
rect 6929 6749 6963 6783
rect 7205 6749 7239 6783
rect 7481 6749 7515 6783
rect 9229 6749 9263 6783
rect 23765 6749 23799 6783
rect 23857 6749 23891 6783
rect 24133 6749 24167 6783
rect 28273 6749 28307 6783
rect 29745 6749 29779 6783
rect 29929 6749 29963 6783
rect 30113 6749 30147 6783
rect 30573 6749 30607 6783
rect 31401 6749 31435 6783
rect 36001 6749 36035 6783
rect 36369 6749 36403 6783
rect 37013 6749 37047 6783
rect 37749 6749 37783 6783
rect 38853 6749 38887 6783
rect 2973 6681 3007 6715
rect 3157 6681 3191 6715
rect 5825 6681 5859 6715
rect 7297 6681 7331 6715
rect 8401 6681 8435 6715
rect 8617 6681 8651 6715
rect 8953 6681 8987 6715
rect 21741 6681 21775 6715
rect 24225 6681 24259 6715
rect 29837 6681 29871 6715
rect 31217 6681 31251 6715
rect 37933 6681 37967 6715
rect 38301 6681 38335 6715
rect 38485 6681 38519 6715
rect 2697 6613 2731 6647
rect 3893 6613 3927 6647
rect 5641 6613 5675 6647
rect 5917 6613 5951 6647
rect 7757 6613 7791 6647
rect 9413 6613 9447 6647
rect 23213 6613 23247 6647
rect 23581 6613 23615 6647
rect 27997 6613 28031 6647
rect 30205 6613 30239 6647
rect 31309 6613 31343 6647
rect 35541 6613 35575 6647
rect 35725 6613 35759 6647
rect 6745 6409 6779 6443
rect 10609 6409 10643 6443
rect 11069 6409 11103 6443
rect 20177 6409 20211 6443
rect 24961 6409 24995 6443
rect 26985 6409 27019 6443
rect 36921 6409 36955 6443
rect 1685 6341 1719 6375
rect 3493 6341 3527 6375
rect 3709 6341 3743 6375
rect 6377 6341 6411 6375
rect 6593 6341 6627 6375
rect 7113 6341 7147 6375
rect 10517 6341 10551 6375
rect 18705 6341 18739 6375
rect 20821 6341 20855 6375
rect 21189 6341 21223 6375
rect 25145 6341 25179 6375
rect 28457 6341 28491 6375
rect 30941 6341 30975 6375
rect 32689 6341 32723 6375
rect 35449 6341 35483 6375
rect 1409 6273 1443 6307
rect 3893 6273 3927 6307
rect 4077 6273 4111 6307
rect 4169 6273 4203 6307
rect 8861 6273 8895 6307
rect 9321 6273 9355 6307
rect 9873 6273 9907 6307
rect 11253 6273 11287 6307
rect 18429 6273 18463 6307
rect 22017 6273 22051 6307
rect 23213 6273 23247 6307
rect 25513 6273 25547 6307
rect 29101 6273 29135 6307
rect 29377 6273 29411 6307
rect 30481 6273 30515 6307
rect 30757 6273 30791 6307
rect 30849 6273 30883 6307
rect 31125 6273 31159 6307
rect 31585 6273 31619 6307
rect 31677 6273 31711 6307
rect 31769 6273 31803 6307
rect 31953 6273 31987 6307
rect 32413 6273 32447 6307
rect 32781 6273 32815 6307
rect 34989 6273 35023 6307
rect 35173 6273 35207 6307
rect 37289 6273 37323 6307
rect 3157 6205 3191 6239
rect 3985 6205 4019 6239
rect 4445 6205 4479 6239
rect 6837 6205 6871 6239
rect 8953 6205 8987 6239
rect 23489 6205 23523 6239
rect 28733 6205 28767 6239
rect 29009 6205 29043 6239
rect 29469 6205 29503 6239
rect 29929 6205 29963 6239
rect 32321 6205 32355 6239
rect 34713 6205 34747 6239
rect 9229 6137 9263 6171
rect 31401 6137 31435 6171
rect 37473 6137 37507 6171
rect 3341 6069 3375 6103
rect 3525 6069 3559 6103
rect 5917 6069 5951 6103
rect 6561 6069 6595 6103
rect 8585 6069 8619 6103
rect 22661 6069 22695 6103
rect 28825 6069 28859 6103
rect 30573 6069 30607 6103
rect 32137 6069 32171 6103
rect 33241 6069 33275 6103
rect 3525 5865 3559 5899
rect 3801 5865 3835 5899
rect 9045 5865 9079 5899
rect 9321 5865 9355 5899
rect 21833 5865 21867 5899
rect 22569 5865 22603 5899
rect 31309 5865 31343 5899
rect 33241 5865 33275 5899
rect 35909 5865 35943 5899
rect 41981 5865 42015 5899
rect 5733 5797 5767 5831
rect 1777 5729 1811 5763
rect 2053 5729 2087 5763
rect 4077 5729 4111 5763
rect 4629 5729 4663 5763
rect 5917 5729 5951 5763
rect 10793 5729 10827 5763
rect 11069 5729 11103 5763
rect 22753 5729 22787 5763
rect 29561 5729 29595 5763
rect 29837 5729 29871 5763
rect 31677 5729 31711 5763
rect 33149 5729 33183 5763
rect 33793 5729 33827 5763
rect 37381 5729 37415 5763
rect 37657 5729 37691 5763
rect 4169 5661 4203 5695
rect 5457 5661 5491 5695
rect 5733 5661 5767 5695
rect 8769 5661 8803 5695
rect 8953 5661 8987 5695
rect 9137 5661 9171 5695
rect 22385 5661 22419 5695
rect 22845 5661 22879 5695
rect 23213 5661 23247 5695
rect 31401 5661 31435 5695
rect 34713 5661 34747 5695
rect 5365 5593 5399 5627
rect 6193 5593 6227 5627
rect 23121 5593 23155 5627
rect 42073 5593 42107 5627
rect 5549 5525 5583 5559
rect 7665 5525 7699 5559
rect 8125 5525 8159 5559
rect 35357 5525 35391 5559
rect 3249 5321 3283 5355
rect 5549 5321 5583 5355
rect 9597 5321 9631 5355
rect 29929 5321 29963 5355
rect 32137 5321 32171 5355
rect 34713 5321 34747 5355
rect 22201 5253 22235 5287
rect 22293 5253 22327 5287
rect 30665 5253 30699 5287
rect 30849 5253 30883 5287
rect 31033 5253 31067 5287
rect 34989 5253 35023 5287
rect 35081 5253 35115 5287
rect 3157 5185 3191 5219
rect 3341 5185 3375 5219
rect 3801 5185 3835 5219
rect 5825 5185 5859 5219
rect 6745 5185 6779 5219
rect 7849 5185 7883 5219
rect 22109 5185 22143 5219
rect 22477 5185 22511 5219
rect 28181 5185 28215 5219
rect 30297 5185 30331 5219
rect 34897 5185 34931 5219
rect 35265 5185 35299 5219
rect 4077 5117 4111 5151
rect 5917 5117 5951 5151
rect 6193 5117 6227 5151
rect 7297 5117 7331 5151
rect 8125 5117 8159 5151
rect 28457 5117 28491 5151
rect 32781 5117 32815 5151
rect 21925 5049 21959 5083
rect 4905 4777 4939 4811
rect 5641 4777 5675 4811
rect 7205 4777 7239 4811
rect 8033 4777 8067 4811
rect 32965 4777 32999 4811
rect 6193 4709 6227 4743
rect 5549 4641 5583 4675
rect 8493 4641 8527 4675
rect 31217 4641 31251 4675
rect 31493 4641 31527 4675
rect 5825 4573 5859 4607
rect 5917 4573 5951 4607
rect 8401 4573 8435 4607
rect 6009 4505 6043 4539
rect 7481 4505 7515 4539
rect 11713 2397 11747 2431
rect 11897 2261 11931 2295
<< metal1 >>
rect 1104 43546 42504 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 35594 43546
rect 35646 43494 35658 43546
rect 35710 43494 35722 43546
rect 35774 43494 35786 43546
rect 35838 43494 35850 43546
rect 35902 43494 42504 43546
rect 1104 43472 42504 43494
rect 20254 43392 20260 43444
rect 20312 43392 20318 43444
rect 20530 43392 20536 43444
rect 20588 43432 20594 43444
rect 20809 43435 20867 43441
rect 20809 43432 20821 43435
rect 20588 43404 20821 43432
rect 20588 43392 20594 43404
rect 20809 43401 20821 43404
rect 20855 43401 20867 43435
rect 20809 43395 20867 43401
rect 21542 43392 21548 43444
rect 21600 43392 21606 43444
rect 22738 43392 22744 43444
rect 22796 43392 22802 43444
rect 24026 43392 24032 43444
rect 24084 43392 24090 43444
rect 21634 43364 21640 43376
rect 21284 43336 21640 43364
rect 19886 43256 19892 43308
rect 19944 43296 19950 43308
rect 20073 43299 20131 43305
rect 20073 43296 20085 43299
rect 19944 43268 20085 43296
rect 19944 43256 19950 43268
rect 20073 43265 20085 43268
rect 20119 43265 20131 43299
rect 20073 43259 20131 43265
rect 20898 43256 20904 43308
rect 20956 43296 20962 43308
rect 20993 43299 21051 43305
rect 20993 43296 21005 43299
rect 20956 43268 21005 43296
rect 20956 43256 20962 43268
rect 20993 43265 21005 43268
rect 21039 43265 21051 43299
rect 20993 43259 21051 43265
rect 21082 43256 21088 43308
rect 21140 43256 21146 43308
rect 21284 43305 21312 43336
rect 21634 43324 21640 43336
rect 21692 43324 21698 43376
rect 21269 43299 21327 43305
rect 21269 43265 21281 43299
rect 21315 43265 21327 43299
rect 21269 43259 21327 43265
rect 21361 43299 21419 43305
rect 21361 43265 21373 43299
rect 21407 43265 21419 43299
rect 21361 43259 21419 43265
rect 22925 43299 22983 43305
rect 22925 43265 22937 43299
rect 22971 43296 22983 43299
rect 23106 43296 23112 43308
rect 22971 43268 23112 43296
rect 22971 43265 22983 43268
rect 22925 43259 22983 43265
rect 21174 43188 21180 43240
rect 21232 43228 21238 43240
rect 21376 43228 21404 43259
rect 23106 43256 23112 43268
rect 23164 43256 23170 43308
rect 23750 43256 23756 43308
rect 23808 43296 23814 43308
rect 24213 43299 24271 43305
rect 24213 43296 24225 43299
rect 23808 43268 24225 43296
rect 23808 43256 23814 43268
rect 24213 43265 24225 43268
rect 24259 43265 24271 43299
rect 24213 43259 24271 43265
rect 21232 43200 21404 43228
rect 21232 43188 21238 43200
rect 26234 43188 26240 43240
rect 26292 43228 26298 43240
rect 26421 43231 26479 43237
rect 26421 43228 26433 43231
rect 26292 43200 26433 43228
rect 26292 43188 26298 43200
rect 26421 43197 26433 43200
rect 26467 43197 26479 43231
rect 26421 43191 26479 43197
rect 33870 43188 33876 43240
rect 33928 43228 33934 43240
rect 34333 43231 34391 43237
rect 34333 43228 34345 43231
rect 33928 43200 34345 43228
rect 33928 43188 33934 43200
rect 34333 43197 34345 43200
rect 34379 43197 34391 43231
rect 34333 43191 34391 43197
rect 21177 43095 21235 43101
rect 21177 43061 21189 43095
rect 21223 43092 21235 43095
rect 21542 43092 21548 43104
rect 21223 43064 21548 43092
rect 21223 43061 21235 43064
rect 21177 43055 21235 43061
rect 21542 43052 21548 43064
rect 21600 43052 21606 43104
rect 25866 43052 25872 43104
rect 25924 43052 25930 43104
rect 33778 43052 33784 43104
rect 33836 43052 33842 43104
rect 1104 43002 42504 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 42504 43002
rect 1104 42928 42504 42950
rect 32388 42891 32446 42897
rect 32388 42857 32400 42891
rect 32434 42888 32446 42891
rect 33134 42888 33140 42900
rect 32434 42860 33140 42888
rect 32434 42857 32446 42860
rect 32388 42851 32446 42857
rect 33134 42848 33140 42860
rect 33192 42848 33198 42900
rect 33870 42848 33876 42900
rect 33928 42848 33934 42900
rect 17862 42780 17868 42832
rect 17920 42820 17926 42832
rect 17920 42792 20668 42820
rect 17920 42780 17926 42792
rect 19904 42761 19932 42792
rect 20640 42761 20668 42792
rect 23566 42780 23572 42832
rect 23624 42820 23630 42832
rect 23624 42792 26648 42820
rect 23624 42780 23630 42792
rect 25792 42761 25820 42792
rect 26620 42761 26648 42792
rect 19889 42755 19947 42761
rect 19889 42721 19901 42755
rect 19935 42721 19947 42755
rect 19889 42715 19947 42721
rect 20625 42755 20683 42761
rect 20625 42721 20637 42755
rect 20671 42721 20683 42755
rect 20625 42715 20683 42721
rect 25777 42755 25835 42761
rect 25777 42721 25789 42755
rect 25823 42721 25835 42755
rect 25777 42715 25835 42721
rect 26605 42755 26663 42761
rect 26605 42721 26617 42755
rect 26651 42721 26663 42755
rect 26605 42715 26663 42721
rect 27065 42755 27123 42761
rect 27065 42721 27077 42755
rect 27111 42752 27123 42755
rect 29546 42752 29552 42764
rect 27111 42724 29552 42752
rect 27111 42721 27123 42724
rect 27065 42715 27123 42721
rect 29546 42712 29552 42724
rect 29604 42712 29610 42764
rect 31297 42755 31355 42761
rect 31297 42721 31309 42755
rect 31343 42752 31355 42755
rect 31754 42752 31760 42764
rect 31343 42724 31760 42752
rect 31343 42721 31355 42724
rect 31297 42715 31355 42721
rect 31754 42712 31760 42724
rect 31812 42752 31818 42764
rect 31941 42755 31999 42761
rect 31941 42752 31953 42755
rect 31812 42724 31953 42752
rect 31812 42712 31818 42724
rect 31941 42721 31953 42724
rect 31987 42721 31999 42755
rect 34330 42752 34336 42764
rect 31941 42715 31999 42721
rect 33520 42724 34336 42752
rect 33520 42696 33548 42724
rect 34330 42712 34336 42724
rect 34388 42712 34394 42764
rect 19705 42687 19763 42693
rect 19705 42653 19717 42687
rect 19751 42684 19763 42687
rect 20162 42684 20168 42696
rect 19751 42656 20168 42684
rect 19751 42653 19763 42656
rect 19705 42647 19763 42653
rect 20162 42644 20168 42656
rect 20220 42644 20226 42696
rect 20441 42687 20499 42693
rect 20441 42653 20453 42687
rect 20487 42684 20499 42687
rect 20901 42687 20959 42693
rect 20901 42684 20913 42687
rect 20487 42656 20913 42684
rect 20487 42653 20499 42656
rect 20441 42647 20499 42653
rect 20901 42653 20913 42656
rect 20947 42653 20959 42687
rect 20901 42647 20959 42653
rect 21450 42644 21456 42696
rect 21508 42644 21514 42696
rect 21729 42687 21787 42693
rect 21729 42653 21741 42687
rect 21775 42653 21787 42687
rect 23934 42684 23940 42696
rect 23138 42656 23940 42684
rect 21729 42647 21787 42653
rect 19426 42576 19432 42628
rect 19484 42616 19490 42628
rect 21744 42616 21772 42647
rect 23934 42644 23940 42656
rect 23992 42644 23998 42696
rect 24213 42687 24271 42693
rect 24213 42653 24225 42687
rect 24259 42684 24271 42687
rect 24670 42684 24676 42696
rect 24259 42656 24676 42684
rect 24259 42653 24271 42656
rect 24213 42647 24271 42653
rect 24670 42644 24676 42656
rect 24728 42644 24734 42696
rect 25593 42687 25651 42693
rect 25593 42653 25605 42687
rect 25639 42684 25651 42687
rect 25866 42684 25872 42696
rect 25639 42656 25872 42684
rect 25639 42653 25651 42656
rect 25593 42647 25651 42653
rect 25866 42644 25872 42656
rect 25924 42644 25930 42696
rect 32122 42644 32128 42696
rect 32180 42644 32186 42696
rect 33502 42644 33508 42696
rect 33560 42644 33566 42696
rect 33962 42644 33968 42696
rect 34020 42684 34026 42696
rect 34701 42687 34759 42693
rect 34701 42684 34713 42687
rect 34020 42656 34713 42684
rect 34020 42644 34026 42656
rect 34701 42653 34713 42656
rect 34747 42653 34759 42687
rect 34701 42647 34759 42653
rect 19484 42588 21772 42616
rect 19484 42576 19490 42588
rect 22002 42576 22008 42628
rect 22060 42576 22066 42628
rect 23290 42576 23296 42628
rect 23348 42616 23354 42628
rect 23569 42619 23627 42625
rect 23569 42616 23581 42619
rect 23348 42588 23581 42616
rect 23348 42576 23354 42588
rect 23569 42585 23581 42588
rect 23615 42585 23627 42619
rect 23569 42579 23627 42585
rect 27341 42619 27399 42625
rect 27341 42585 27353 42619
rect 27387 42616 27399 42619
rect 27614 42616 27620 42628
rect 27387 42588 27620 42616
rect 27387 42585 27399 42588
rect 27341 42579 27399 42585
rect 27614 42576 27620 42588
rect 27672 42576 27678 42628
rect 28718 42616 28724 42628
rect 28566 42588 28724 42616
rect 28718 42576 28724 42588
rect 28776 42576 28782 42628
rect 29822 42576 29828 42628
rect 29880 42576 29886 42628
rect 30466 42576 30472 42628
rect 30524 42576 30530 42628
rect 33704 42588 34008 42616
rect 19245 42551 19303 42557
rect 19245 42517 19257 42551
rect 19291 42548 19303 42551
rect 19518 42548 19524 42560
rect 19291 42520 19524 42548
rect 19291 42517 19303 42520
rect 19245 42511 19303 42517
rect 19518 42508 19524 42520
rect 19576 42508 19582 42560
rect 19610 42508 19616 42560
rect 19668 42508 19674 42560
rect 19794 42508 19800 42560
rect 19852 42548 19858 42560
rect 20073 42551 20131 42557
rect 20073 42548 20085 42551
rect 19852 42520 20085 42548
rect 19852 42508 19858 42520
rect 20073 42517 20085 42520
rect 20119 42517 20131 42551
rect 20073 42511 20131 42517
rect 20438 42508 20444 42560
rect 20496 42548 20502 42560
rect 20533 42551 20591 42557
rect 20533 42548 20545 42551
rect 20496 42520 20545 42548
rect 20496 42508 20502 42520
rect 20533 42517 20545 42520
rect 20579 42517 20591 42551
rect 20533 42511 20591 42517
rect 23474 42508 23480 42560
rect 23532 42508 23538 42560
rect 24578 42508 24584 42560
rect 24636 42548 24642 42560
rect 25225 42551 25283 42557
rect 25225 42548 25237 42551
rect 24636 42520 25237 42548
rect 24636 42508 24642 42520
rect 25225 42517 25237 42520
rect 25271 42517 25283 42551
rect 25225 42511 25283 42517
rect 25685 42551 25743 42557
rect 25685 42517 25697 42551
rect 25731 42548 25743 42551
rect 25866 42548 25872 42560
rect 25731 42520 25872 42548
rect 25731 42517 25743 42520
rect 25685 42511 25743 42517
rect 25866 42508 25872 42520
rect 25924 42508 25930 42560
rect 26050 42508 26056 42560
rect 26108 42508 26114 42560
rect 26418 42508 26424 42560
rect 26476 42508 26482 42560
rect 26513 42551 26571 42557
rect 26513 42517 26525 42551
rect 26559 42548 26571 42551
rect 26786 42548 26792 42560
rect 26559 42520 26792 42548
rect 26559 42517 26571 42520
rect 26513 42511 26571 42517
rect 26786 42508 26792 42520
rect 26844 42508 26850 42560
rect 28813 42551 28871 42557
rect 28813 42517 28825 42551
rect 28859 42548 28871 42551
rect 28994 42548 29000 42560
rect 28859 42520 29000 42548
rect 28859 42517 28871 42520
rect 28813 42511 28871 42517
rect 28994 42508 29000 42520
rect 29052 42508 29058 42560
rect 31386 42508 31392 42560
rect 31444 42508 31450 42560
rect 33226 42508 33232 42560
rect 33284 42548 33290 42560
rect 33704 42548 33732 42588
rect 33980 42557 34008 42588
rect 34054 42576 34060 42628
rect 34112 42576 34118 42628
rect 34146 42576 34152 42628
rect 34204 42616 34210 42628
rect 34241 42619 34299 42625
rect 34241 42616 34253 42619
rect 34204 42588 34253 42616
rect 34204 42576 34210 42588
rect 34241 42585 34253 42588
rect 34287 42585 34299 42619
rect 34241 42579 34299 42585
rect 33284 42520 33732 42548
rect 33965 42551 34023 42557
rect 33284 42508 33290 42520
rect 33965 42517 33977 42551
rect 34011 42517 34023 42551
rect 33965 42511 34023 42517
rect 35342 42508 35348 42560
rect 35400 42508 35406 42560
rect 1104 42458 42504 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 35594 42458
rect 35646 42406 35658 42458
rect 35710 42406 35722 42458
rect 35774 42406 35786 42458
rect 35838 42406 35850 42458
rect 35902 42406 42504 42458
rect 1104 42384 42504 42406
rect 21177 42347 21235 42353
rect 21177 42313 21189 42347
rect 21223 42344 21235 42347
rect 21450 42344 21456 42356
rect 21223 42316 21456 42344
rect 21223 42313 21235 42316
rect 21177 42307 21235 42313
rect 21450 42304 21456 42316
rect 21508 42304 21514 42356
rect 26053 42347 26111 42353
rect 22204 42316 24348 42344
rect 19705 42279 19763 42285
rect 19705 42245 19717 42279
rect 19751 42276 19763 42279
rect 19794 42276 19800 42288
rect 19751 42248 19800 42276
rect 19751 42245 19763 42248
rect 19705 42239 19763 42245
rect 19794 42236 19800 42248
rect 19852 42236 19858 42288
rect 20254 42236 20260 42288
rect 20312 42236 20318 42288
rect 21082 42236 21088 42288
rect 21140 42276 21146 42288
rect 21269 42279 21327 42285
rect 21269 42276 21281 42279
rect 21140 42248 21281 42276
rect 21140 42236 21146 42248
rect 21269 42245 21281 42248
rect 21315 42245 21327 42279
rect 21269 42239 21327 42245
rect 19426 42168 19432 42220
rect 19484 42168 19490 42220
rect 21453 42211 21511 42217
rect 21453 42177 21465 42211
rect 21499 42208 21511 42211
rect 21634 42208 21640 42220
rect 21499 42180 21640 42208
rect 21499 42177 21511 42180
rect 21453 42171 21511 42177
rect 21634 42168 21640 42180
rect 21692 42168 21698 42220
rect 22204 42217 22232 42316
rect 23934 42276 23940 42288
rect 23690 42248 23940 42276
rect 23934 42236 23940 42248
rect 23992 42236 23998 42288
rect 24320 42220 24348 42316
rect 26053 42313 26065 42347
rect 26099 42344 26111 42347
rect 26234 42344 26240 42356
rect 26099 42316 26240 42344
rect 26099 42313 26111 42316
rect 26053 42307 26111 42313
rect 26234 42304 26240 42316
rect 26292 42304 26298 42356
rect 26418 42304 26424 42356
rect 26476 42344 26482 42356
rect 26789 42347 26847 42353
rect 26789 42344 26801 42347
rect 26476 42316 26801 42344
rect 26476 42304 26482 42316
rect 26789 42313 26801 42316
rect 26835 42313 26847 42347
rect 26789 42307 26847 42313
rect 27614 42304 27620 42356
rect 27672 42304 27678 42356
rect 29822 42304 29828 42356
rect 29880 42344 29886 42356
rect 29917 42347 29975 42353
rect 29917 42344 29929 42347
rect 29880 42316 29929 42344
rect 29880 42304 29886 42316
rect 29917 42313 29929 42316
rect 29963 42313 29975 42347
rect 29917 42307 29975 42313
rect 30285 42347 30343 42353
rect 30285 42313 30297 42347
rect 30331 42344 30343 42347
rect 31386 42344 31392 42356
rect 30331 42316 31392 42344
rect 30331 42313 30343 42316
rect 30285 42307 30343 42313
rect 31386 42304 31392 42316
rect 31444 42304 31450 42356
rect 31478 42304 31484 42356
rect 31536 42344 31542 42356
rect 31536 42316 32904 42344
rect 31536 42304 31542 42316
rect 24578 42236 24584 42288
rect 24636 42236 24642 42288
rect 26252 42276 26280 42304
rect 26878 42276 26884 42288
rect 26252 42248 26884 42276
rect 26878 42236 26884 42248
rect 26936 42276 26942 42288
rect 31113 42279 31171 42285
rect 26936 42248 27200 42276
rect 26936 42236 26942 42248
rect 22189 42211 22247 42217
rect 22189 42177 22201 42211
rect 22235 42177 22247 42211
rect 22189 42171 22247 42177
rect 24302 42168 24308 42220
rect 24360 42168 24366 42220
rect 25682 42168 25688 42220
rect 25740 42168 25746 42220
rect 26694 42168 26700 42220
rect 26752 42208 26758 42220
rect 27172 42217 27200 42248
rect 31113 42245 31125 42279
rect 31159 42276 31171 42279
rect 31159 42248 31800 42276
rect 31159 42245 31171 42248
rect 31113 42239 31171 42245
rect 31772 42220 31800 42248
rect 26973 42211 27031 42217
rect 26973 42208 26985 42211
rect 26752 42180 26985 42208
rect 26752 42168 26758 42180
rect 26973 42177 26985 42180
rect 27019 42177 27031 42211
rect 26973 42171 27031 42177
rect 27157 42211 27215 42217
rect 27157 42177 27169 42211
rect 27203 42177 27215 42211
rect 27157 42171 27215 42177
rect 27985 42211 28043 42217
rect 27985 42177 27997 42211
rect 28031 42208 28043 42211
rect 28445 42211 28503 42217
rect 28445 42208 28457 42211
rect 28031 42180 28457 42208
rect 28031 42177 28043 42180
rect 27985 42171 28043 42177
rect 28445 42177 28457 42180
rect 28491 42177 28503 42211
rect 28445 42171 28503 42177
rect 28994 42168 29000 42220
rect 29052 42168 29058 42220
rect 30834 42168 30840 42220
rect 30892 42208 30898 42220
rect 30929 42211 30987 42217
rect 30929 42208 30941 42211
rect 30892 42180 30941 42208
rect 30892 42168 30898 42180
rect 30929 42177 30941 42180
rect 30975 42177 30987 42211
rect 30929 42171 30987 42177
rect 31202 42168 31208 42220
rect 31260 42168 31266 42220
rect 31389 42214 31447 42217
rect 31312 42211 31447 42214
rect 31312 42186 31401 42211
rect 31312 42152 31340 42186
rect 31389 42177 31401 42186
rect 31435 42177 31447 42211
rect 31389 42171 31447 42177
rect 31481 42211 31539 42217
rect 31481 42177 31493 42211
rect 31527 42177 31539 42211
rect 31481 42171 31539 42177
rect 22462 42100 22468 42152
rect 22520 42100 22526 42152
rect 26234 42100 26240 42152
rect 26292 42100 26298 42152
rect 27706 42100 27712 42152
rect 27764 42140 27770 42152
rect 28077 42143 28135 42149
rect 28077 42140 28089 42143
rect 27764 42112 28089 42140
rect 27764 42100 27770 42112
rect 28077 42109 28089 42112
rect 28123 42109 28135 42143
rect 28077 42103 28135 42109
rect 28169 42143 28227 42149
rect 28169 42109 28181 42143
rect 28215 42109 28227 42143
rect 28169 42103 28227 42109
rect 27890 42032 27896 42084
rect 27948 42072 27954 42084
rect 28184 42072 28212 42103
rect 30098 42100 30104 42152
rect 30156 42140 30162 42152
rect 30377 42143 30435 42149
rect 30377 42140 30389 42143
rect 30156 42112 30389 42140
rect 30156 42100 30162 42112
rect 30377 42109 30389 42112
rect 30423 42109 30435 42143
rect 30377 42103 30435 42109
rect 30469 42143 30527 42149
rect 30469 42109 30481 42143
rect 30515 42109 30527 42143
rect 30469 42103 30527 42109
rect 30745 42143 30803 42149
rect 30745 42109 30757 42143
rect 30791 42140 30803 42143
rect 31294 42140 31300 42152
rect 30791 42112 31300 42140
rect 30791 42109 30803 42112
rect 30745 42103 30803 42109
rect 30484 42072 30512 42103
rect 31294 42100 31300 42112
rect 31352 42100 31358 42152
rect 31496 42140 31524 42171
rect 31570 42168 31576 42220
rect 31628 42168 31634 42220
rect 31754 42168 31760 42220
rect 31812 42168 31818 42220
rect 32876 42217 32904 42316
rect 33134 42304 33140 42356
rect 33192 42304 33198 42356
rect 33505 42347 33563 42353
rect 33505 42313 33517 42347
rect 33551 42344 33563 42347
rect 33778 42344 33784 42356
rect 33551 42316 33784 42344
rect 33551 42313 33563 42316
rect 33505 42307 33563 42313
rect 33778 42304 33784 42316
rect 33836 42304 33842 42356
rect 33962 42304 33968 42356
rect 34020 42304 34026 42356
rect 32953 42279 33011 42285
rect 32953 42245 32965 42279
rect 32999 42276 33011 42279
rect 34146 42276 34152 42288
rect 32999 42248 34152 42276
rect 32999 42245 33011 42248
rect 32953 42239 33011 42245
rect 34146 42236 34152 42248
rect 34204 42236 34210 42288
rect 32861 42211 32919 42217
rect 32861 42177 32873 42211
rect 32907 42177 32919 42211
rect 32861 42171 32919 42177
rect 33045 42211 33103 42217
rect 33045 42177 33057 42211
rect 33091 42208 33103 42211
rect 33870 42208 33876 42220
rect 33091 42180 33876 42208
rect 33091 42177 33103 42180
rect 33045 42171 33103 42177
rect 33870 42168 33876 42180
rect 33928 42168 33934 42220
rect 34330 42168 34336 42220
rect 34388 42168 34394 42220
rect 31846 42140 31852 42152
rect 31496 42112 31852 42140
rect 31846 42100 31852 42112
rect 31904 42100 31910 42152
rect 33594 42100 33600 42152
rect 33652 42100 33658 42152
rect 33689 42143 33747 42149
rect 33689 42109 33701 42143
rect 33735 42109 33747 42143
rect 33689 42103 33747 42109
rect 30650 42072 30656 42084
rect 27948 42044 30656 42072
rect 27948 42032 27954 42044
rect 30650 42032 30656 42044
rect 30708 42072 30714 42084
rect 33704 42072 33732 42103
rect 34698 42100 34704 42152
rect 34756 42140 34762 42152
rect 35437 42143 35495 42149
rect 35437 42140 35449 42143
rect 34756 42112 35449 42140
rect 34756 42100 34762 42112
rect 35437 42109 35449 42112
rect 35483 42109 35495 42143
rect 35437 42103 35495 42109
rect 35713 42143 35771 42149
rect 35713 42109 35725 42143
rect 35759 42140 35771 42143
rect 35759 42112 35894 42140
rect 35759 42109 35771 42112
rect 35713 42103 35771 42109
rect 30708 42044 33732 42072
rect 35866 42072 35894 42112
rect 37458 42100 37464 42152
rect 37516 42140 37522 42152
rect 38289 42143 38347 42149
rect 38289 42140 38301 42143
rect 37516 42112 38301 42140
rect 37516 42100 37522 42112
rect 38289 42109 38301 42112
rect 38335 42109 38347 42143
rect 38289 42103 38347 42109
rect 38562 42100 38568 42152
rect 38620 42140 38626 42152
rect 38841 42143 38899 42149
rect 38841 42140 38853 42143
rect 38620 42112 38853 42140
rect 38620 42100 38626 42112
rect 38841 42109 38853 42112
rect 38887 42109 38899 42143
rect 38841 42103 38899 42109
rect 35986 42072 35992 42084
rect 35866 42044 35992 42072
rect 30708 42032 30714 42044
rect 35986 42032 35992 42044
rect 36044 42032 36050 42084
rect 21637 42007 21695 42013
rect 21637 41973 21649 42007
rect 21683 42004 21695 42007
rect 21910 42004 21916 42016
rect 21683 41976 21916 42004
rect 21683 41973 21695 41976
rect 21637 41967 21695 41973
rect 21910 41964 21916 41976
rect 21968 41964 21974 42016
rect 22554 41964 22560 42016
rect 22612 42004 22618 42016
rect 23937 42007 23995 42013
rect 23937 42004 23949 42007
rect 22612 41976 23949 42004
rect 22612 41964 22618 41976
rect 23937 41973 23949 41976
rect 23983 42004 23995 42007
rect 24670 42004 24676 42016
rect 23983 41976 24676 42004
rect 23983 41973 23995 41976
rect 23937 41967 23995 41973
rect 24670 41964 24676 41976
rect 24728 41964 24734 42016
rect 27062 41964 27068 42016
rect 27120 41964 27126 42016
rect 31205 42007 31263 42013
rect 31205 41973 31217 42007
rect 31251 42004 31263 42007
rect 31570 42004 31576 42016
rect 31251 41976 31576 42004
rect 31251 41973 31263 41976
rect 31205 41967 31263 41973
rect 31570 41964 31576 41976
rect 31628 41964 31634 42016
rect 31665 42007 31723 42013
rect 31665 41973 31677 42007
rect 31711 42004 31723 42007
rect 31846 42004 31852 42016
rect 31711 41976 31852 42004
rect 31711 41973 31723 41976
rect 31665 41967 31723 41973
rect 31846 41964 31852 41976
rect 31904 41964 31910 42016
rect 37734 41964 37740 42016
rect 37792 41964 37798 42016
rect 39482 41964 39488 42016
rect 39540 41964 39546 42016
rect 1104 41914 42504 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 42504 41914
rect 1104 41840 42504 41862
rect 19610 41760 19616 41812
rect 19668 41800 19674 41812
rect 21085 41803 21143 41809
rect 21085 41800 21097 41803
rect 19668 41772 21097 41800
rect 19668 41760 19674 41772
rect 21085 41769 21097 41772
rect 21131 41769 21143 41803
rect 21085 41763 21143 41769
rect 22462 41760 22468 41812
rect 22520 41800 22526 41812
rect 22649 41803 22707 41809
rect 22649 41800 22661 41803
rect 22520 41772 22661 41800
rect 22520 41760 22526 41772
rect 22649 41769 22661 41772
rect 22695 41769 22707 41803
rect 22649 41763 22707 41769
rect 23934 41760 23940 41812
rect 23992 41800 23998 41812
rect 25682 41800 25688 41812
rect 23992 41772 25688 41800
rect 23992 41760 23998 41772
rect 25682 41760 25688 41772
rect 25740 41760 25746 41812
rect 26234 41760 26240 41812
rect 26292 41800 26298 41812
rect 26513 41803 26571 41809
rect 26513 41800 26525 41803
rect 26292 41772 26525 41800
rect 26292 41760 26298 41772
rect 26513 41769 26525 41772
rect 26559 41769 26571 41803
rect 26513 41763 26571 41769
rect 28718 41760 28724 41812
rect 28776 41800 28782 41812
rect 30466 41800 30472 41812
rect 28776 41772 30472 41800
rect 28776 41760 28782 41772
rect 30466 41760 30472 41772
rect 30524 41760 30530 41812
rect 31202 41760 31208 41812
rect 31260 41800 31266 41812
rect 31478 41800 31484 41812
rect 31260 41772 31484 41800
rect 31260 41760 31266 41772
rect 31478 41760 31484 41772
rect 31536 41760 31542 41812
rect 34054 41760 34060 41812
rect 34112 41760 34118 41812
rect 34698 41760 34704 41812
rect 34756 41760 34762 41812
rect 23566 41732 23572 41744
rect 23216 41704 23572 41732
rect 16853 41667 16911 41673
rect 16853 41633 16865 41667
rect 16899 41664 16911 41667
rect 16899 41636 19288 41664
rect 16899 41633 16911 41636
rect 16853 41627 16911 41633
rect 19260 41605 19288 41636
rect 19518 41624 19524 41676
rect 19576 41624 19582 41676
rect 20993 41667 21051 41673
rect 20993 41633 21005 41667
rect 21039 41664 21051 41667
rect 21082 41664 21088 41676
rect 21039 41636 21088 41664
rect 21039 41633 21051 41636
rect 20993 41627 21051 41633
rect 21082 41624 21088 41636
rect 21140 41624 21146 41676
rect 21450 41624 21456 41676
rect 21508 41664 21514 41676
rect 23216 41673 23244 41704
rect 23566 41692 23572 41704
rect 23624 41692 23630 41744
rect 24578 41692 24584 41744
rect 24636 41732 24642 41744
rect 24673 41735 24731 41741
rect 24673 41732 24685 41735
rect 24636 41704 24685 41732
rect 24636 41692 24642 41704
rect 24673 41701 24685 41704
rect 24719 41701 24731 41735
rect 24673 41695 24731 41701
rect 28074 41692 28080 41744
rect 28132 41732 28138 41744
rect 28445 41735 28503 41741
rect 28445 41732 28457 41735
rect 28132 41704 28457 41732
rect 28132 41692 28138 41704
rect 28445 41701 28457 41704
rect 28491 41701 28503 41735
rect 28445 41695 28503 41701
rect 28994 41692 29000 41744
rect 29052 41692 29058 41744
rect 31110 41692 31116 41744
rect 31168 41732 31174 41744
rect 31573 41735 31631 41741
rect 31573 41732 31585 41735
rect 31168 41704 31585 41732
rect 31168 41692 31174 41704
rect 31573 41701 31585 41704
rect 31619 41701 31631 41735
rect 31573 41695 31631 41701
rect 31662 41692 31668 41744
rect 31720 41732 31726 41744
rect 31720 41704 33456 41732
rect 31720 41692 31726 41704
rect 23201 41667 23259 41673
rect 21508 41636 21864 41664
rect 21508 41624 21514 41636
rect 19245 41599 19303 41605
rect 19245 41565 19257 41599
rect 19291 41565 19303 41599
rect 21100 41596 21128 41624
rect 21836 41605 21864 41636
rect 23201 41633 23213 41667
rect 23247 41633 23259 41667
rect 23201 41627 23259 41633
rect 23474 41624 23480 41676
rect 23532 41664 23538 41676
rect 23842 41664 23848 41676
rect 23532 41636 23848 41664
rect 23532 41624 23538 41636
rect 23842 41624 23848 41636
rect 23900 41664 23906 41676
rect 24029 41667 24087 41673
rect 24029 41664 24041 41667
rect 23900 41636 24041 41664
rect 23900 41624 23906 41636
rect 24029 41633 24041 41636
rect 24075 41633 24087 41667
rect 24029 41627 24087 41633
rect 24302 41624 24308 41676
rect 24360 41664 24366 41676
rect 24765 41667 24823 41673
rect 24765 41664 24777 41667
rect 24360 41636 24777 41664
rect 24360 41624 24366 41636
rect 24765 41633 24777 41636
rect 24811 41633 24823 41667
rect 24765 41627 24823 41633
rect 25041 41667 25099 41673
rect 25041 41633 25053 41667
rect 25087 41664 25099 41667
rect 26050 41664 26056 41676
rect 25087 41636 26056 41664
rect 25087 41633 25099 41636
rect 25041 41627 25099 41633
rect 26050 41624 26056 41636
rect 26108 41624 26114 41676
rect 29012 41664 29040 41692
rect 28092 41636 29040 41664
rect 21637 41599 21695 41605
rect 21637 41596 21649 41599
rect 21100 41568 21649 41596
rect 19245 41559 19303 41565
rect 21637 41565 21649 41568
rect 21683 41565 21695 41599
rect 21637 41559 21695 41565
rect 21821 41599 21879 41605
rect 21821 41565 21833 41599
rect 21867 41565 21879 41599
rect 21821 41559 21879 41565
rect 17126 41488 17132 41540
rect 17184 41488 17190 41540
rect 19260 41528 19288 41559
rect 21910 41556 21916 41608
rect 21968 41556 21974 41608
rect 22554 41556 22560 41608
rect 22612 41556 22618 41608
rect 23017 41599 23075 41605
rect 23017 41565 23029 41599
rect 23063 41596 23075 41599
rect 23290 41596 23296 41608
rect 23063 41568 23296 41596
rect 23063 41565 23075 41568
rect 23017 41559 23075 41565
rect 23290 41556 23296 41568
rect 23348 41556 23354 41608
rect 24394 41556 24400 41608
rect 24452 41556 24458 41608
rect 24670 41556 24676 41608
rect 24728 41556 24734 41608
rect 26878 41556 26884 41608
rect 26936 41596 26942 41608
rect 26973 41599 27031 41605
rect 26973 41596 26985 41599
rect 26936 41568 26985 41596
rect 26936 41556 26942 41568
rect 26973 41565 26985 41568
rect 27019 41565 27031 41599
rect 26973 41559 27031 41565
rect 19426 41528 19432 41540
rect 18354 41500 19196 41528
rect 19260 41500 19432 41528
rect 18598 41420 18604 41472
rect 18656 41420 18662 41472
rect 19168 41460 19196 41500
rect 19426 41488 19432 41500
rect 19484 41488 19490 41540
rect 19978 41528 19984 41540
rect 19904 41500 19984 41528
rect 19904 41460 19932 41500
rect 19978 41488 19984 41500
rect 20036 41488 20042 41540
rect 21542 41488 21548 41540
rect 21600 41528 21606 41540
rect 22097 41531 22155 41537
rect 22097 41528 22109 41531
rect 21600 41500 22109 41528
rect 21600 41488 21606 41500
rect 22097 41497 22109 41500
rect 22143 41497 22155 41531
rect 22097 41491 22155 41497
rect 22281 41531 22339 41537
rect 22281 41497 22293 41531
rect 22327 41528 22339 41531
rect 22370 41528 22376 41540
rect 22327 41500 22376 41528
rect 22327 41497 22339 41500
rect 22281 41491 22339 41497
rect 22370 41488 22376 41500
rect 22428 41488 22434 41540
rect 22465 41531 22523 41537
rect 22465 41497 22477 41531
rect 22511 41528 22523 41531
rect 22511 41500 22876 41528
rect 22511 41497 22523 41500
rect 22465 41491 22523 41497
rect 20254 41460 20260 41472
rect 19168 41432 20260 41460
rect 20254 41420 20260 41432
rect 20312 41420 20318 41472
rect 21082 41420 21088 41472
rect 21140 41460 21146 41472
rect 21821 41463 21879 41469
rect 21821 41460 21833 41463
rect 21140 41432 21833 41460
rect 21140 41420 21146 41432
rect 21821 41429 21833 41432
rect 21867 41429 21879 41463
rect 21821 41423 21879 41429
rect 22554 41420 22560 41472
rect 22612 41420 22618 41472
rect 22848 41460 22876 41500
rect 22922 41488 22928 41540
rect 22980 41528 22986 41540
rect 23109 41531 23167 41537
rect 23109 41528 23121 41531
rect 22980 41500 23121 41528
rect 22980 41488 22986 41500
rect 23109 41497 23121 41500
rect 23155 41497 23167 41531
rect 23566 41528 23572 41540
rect 23109 41491 23167 41497
rect 23400 41500 23572 41528
rect 23400 41460 23428 41500
rect 23566 41488 23572 41500
rect 23624 41528 23630 41540
rect 24489 41531 24547 41537
rect 24489 41528 24501 41531
rect 23624 41500 24501 41528
rect 23624 41488 23630 41500
rect 24489 41497 24501 41500
rect 24535 41497 24547 41531
rect 24489 41491 24547 41497
rect 25682 41488 25688 41540
rect 25740 41488 25746 41540
rect 26694 41528 26700 41540
rect 26344 41500 26700 41528
rect 22848 41432 23428 41460
rect 23474 41420 23480 41472
rect 23532 41420 23538 41472
rect 24762 41420 24768 41472
rect 24820 41460 24826 41472
rect 26344 41460 26372 41500
rect 26694 41488 26700 41500
rect 26752 41528 26758 41540
rect 26789 41531 26847 41537
rect 26789 41528 26801 41531
rect 26752 41500 26801 41528
rect 26752 41488 26758 41500
rect 26789 41497 26801 41500
rect 26835 41497 26847 41531
rect 28092 41528 28120 41636
rect 28166 41556 28172 41608
rect 28224 41596 28230 41608
rect 28828 41605 28856 41636
rect 29546 41624 29552 41676
rect 29604 41664 29610 41676
rect 29730 41664 29736 41676
rect 29604 41636 29736 41664
rect 29604 41624 29610 41636
rect 29730 41624 29736 41636
rect 29788 41624 29794 41676
rect 31294 41624 31300 41676
rect 31352 41664 31358 41676
rect 31352 41636 31708 41664
rect 31352 41624 31358 41636
rect 28537 41599 28595 41605
rect 28537 41596 28549 41599
rect 28224 41568 28549 41596
rect 28224 41556 28230 41568
rect 28537 41565 28549 41568
rect 28583 41565 28595 41599
rect 28537 41559 28595 41565
rect 28813 41599 28871 41605
rect 28813 41565 28825 41599
rect 28859 41565 28871 41599
rect 28813 41559 28871 41565
rect 28997 41599 29055 41605
rect 28997 41565 29009 41599
rect 29043 41596 29055 41599
rect 29270 41596 29276 41608
rect 29043 41568 29276 41596
rect 29043 41565 29055 41568
rect 28997 41559 29055 41565
rect 29270 41556 29276 41568
rect 29328 41556 29334 41608
rect 31478 41556 31484 41608
rect 31536 41596 31542 41608
rect 31680 41605 31708 41636
rect 31754 41624 31760 41676
rect 31812 41664 31818 41676
rect 32858 41664 32864 41676
rect 31812 41636 32864 41664
rect 31812 41624 31818 41636
rect 32858 41624 32864 41636
rect 32916 41664 32922 41676
rect 33045 41667 33103 41673
rect 33045 41664 33057 41667
rect 32916 41636 33057 41664
rect 32916 41624 32922 41636
rect 33045 41633 33057 41636
rect 33091 41633 33103 41667
rect 33045 41627 33103 41633
rect 33137 41667 33195 41673
rect 33137 41633 33149 41667
rect 33183 41664 33195 41667
rect 33318 41664 33324 41676
rect 33183 41636 33324 41664
rect 33183 41633 33195 41636
rect 33137 41627 33195 41633
rect 33318 41624 33324 41636
rect 33376 41624 33382 41676
rect 31573 41599 31631 41605
rect 31573 41596 31585 41599
rect 31536 41568 31585 41596
rect 31536 41556 31542 41568
rect 31573 41565 31585 41568
rect 31619 41565 31631 41599
rect 31573 41559 31631 41565
rect 31665 41599 31723 41605
rect 31665 41565 31677 41599
rect 31711 41565 31723 41599
rect 31665 41559 31723 41565
rect 31846 41556 31852 41608
rect 31904 41556 31910 41608
rect 32953 41599 33011 41605
rect 32953 41565 32965 41599
rect 32999 41565 33011 41599
rect 32953 41559 33011 41565
rect 28445 41531 28503 41537
rect 28445 41528 28457 41531
rect 28092 41500 28457 41528
rect 26789 41491 26847 41497
rect 28445 41497 28457 41500
rect 28491 41497 28503 41531
rect 28721 41531 28779 41537
rect 28721 41528 28733 41531
rect 28445 41491 28503 41497
rect 28552 41500 28733 41528
rect 24820 41432 26372 41460
rect 24820 41420 24826 41432
rect 26602 41420 26608 41472
rect 26660 41420 26666 41472
rect 28261 41463 28319 41469
rect 28261 41429 28273 41463
rect 28307 41460 28319 41463
rect 28552 41460 28580 41500
rect 28721 41497 28733 41500
rect 28767 41497 28779 41531
rect 28721 41491 28779 41497
rect 28307 41432 28580 41460
rect 28307 41429 28319 41432
rect 28261 41423 28319 41429
rect 28626 41420 28632 41472
rect 28684 41420 28690 41472
rect 28736 41460 28764 41491
rect 29178 41488 29184 41540
rect 29236 41528 29242 41540
rect 29236 41500 29960 41528
rect 29236 41488 29242 41500
rect 29365 41463 29423 41469
rect 29365 41460 29377 41463
rect 28736 41432 29377 41460
rect 29365 41429 29377 41432
rect 29411 41429 29423 41463
rect 29932 41460 29960 41500
rect 30006 41488 30012 41540
rect 30064 41488 30070 41540
rect 30466 41488 30472 41540
rect 30524 41488 30530 41540
rect 32968 41528 32996 41559
rect 33226 41556 33232 41608
rect 33284 41556 33290 41608
rect 33428 41596 33456 41704
rect 33870 41664 33876 41676
rect 33704 41636 33876 41664
rect 33704 41605 33732 41636
rect 33870 41624 33876 41636
rect 33928 41624 33934 41676
rect 34072 41664 34100 41760
rect 34422 41692 34428 41744
rect 34480 41692 34486 41744
rect 35345 41667 35403 41673
rect 34072 41636 34284 41664
rect 33689 41599 33747 41605
rect 33428 41568 33548 41596
rect 33410 41528 33416 41540
rect 32968 41500 33416 41528
rect 33410 41488 33416 41500
rect 33468 41488 33474 41540
rect 33520 41528 33548 41568
rect 33689 41565 33701 41599
rect 33735 41565 33747 41599
rect 33689 41559 33747 41565
rect 34146 41556 34152 41608
rect 34204 41556 34210 41608
rect 34256 41605 34284 41636
rect 35345 41633 35357 41667
rect 35391 41664 35403 41667
rect 38010 41664 38016 41676
rect 35391 41636 38016 41664
rect 35391 41633 35403 41636
rect 35345 41627 35403 41633
rect 38010 41624 38016 41636
rect 38068 41624 38074 41676
rect 39022 41624 39028 41676
rect 39080 41664 39086 41676
rect 39669 41667 39727 41673
rect 39669 41664 39681 41667
rect 39080 41636 39681 41664
rect 39080 41624 39086 41636
rect 39669 41633 39681 41636
rect 39715 41633 39727 41667
rect 39669 41627 39727 41633
rect 34241 41599 34299 41605
rect 34241 41565 34253 41599
rect 34287 41565 34299 41599
rect 34241 41559 34299 41565
rect 37458 41556 37464 41608
rect 37516 41556 37522 41608
rect 33873 41531 33931 41537
rect 33873 41528 33885 41531
rect 33520 41500 33885 41528
rect 33873 41497 33885 41500
rect 33919 41497 33931 41531
rect 33873 41491 33931 41497
rect 33962 41488 33968 41540
rect 34020 41528 34026 41540
rect 34425 41531 34483 41537
rect 34425 41528 34437 41531
rect 34020 41500 34437 41528
rect 34020 41488 34026 41500
rect 34425 41497 34437 41500
rect 34471 41497 34483 41531
rect 34425 41491 34483 41497
rect 35069 41531 35127 41537
rect 35069 41497 35081 41531
rect 35115 41528 35127 41531
rect 35342 41528 35348 41540
rect 35115 41500 35348 41528
rect 35115 41497 35127 41500
rect 35069 41491 35127 41497
rect 35342 41488 35348 41500
rect 35400 41488 35406 41540
rect 37553 41531 37611 41537
rect 37553 41497 37565 41531
rect 37599 41528 37611 41531
rect 37642 41528 37648 41540
rect 37599 41500 37648 41528
rect 37599 41497 37611 41500
rect 37553 41491 37611 41497
rect 37642 41488 37648 41500
rect 37700 41488 37706 41540
rect 37737 41531 37795 41537
rect 37737 41497 37749 41531
rect 37783 41528 37795 41531
rect 37826 41528 37832 41540
rect 37783 41500 37832 41528
rect 37783 41497 37795 41500
rect 37737 41491 37795 41497
rect 37826 41488 37832 41500
rect 37884 41488 37890 41540
rect 38102 41488 38108 41540
rect 38160 41528 38166 41540
rect 38160 41500 38226 41528
rect 38160 41488 38166 41500
rect 39390 41488 39396 41540
rect 39448 41488 39454 41540
rect 30834 41460 30840 41472
rect 29932 41432 30840 41460
rect 29365 41423 29423 41429
rect 30834 41420 30840 41432
rect 30892 41420 30898 41472
rect 31478 41420 31484 41472
rect 31536 41460 31542 41472
rect 31662 41460 31668 41472
rect 31536 41432 31668 41460
rect 31536 41420 31542 41432
rect 31662 41420 31668 41432
rect 31720 41420 31726 41472
rect 32766 41420 32772 41472
rect 32824 41420 32830 41472
rect 35158 41420 35164 41472
rect 35216 41420 35222 41472
rect 37458 41420 37464 41472
rect 37516 41420 37522 41472
rect 37918 41420 37924 41472
rect 37976 41420 37982 41472
rect 1104 41370 42504 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 35594 41370
rect 35646 41318 35658 41370
rect 35710 41318 35722 41370
rect 35774 41318 35786 41370
rect 35838 41318 35850 41370
rect 35902 41318 42504 41370
rect 1104 41296 42504 41318
rect 17126 41216 17132 41268
rect 17184 41256 17190 41268
rect 17497 41259 17555 41265
rect 17497 41256 17509 41259
rect 17184 41228 17509 41256
rect 17184 41216 17190 41228
rect 17497 41225 17509 41228
rect 17543 41225 17555 41259
rect 17497 41219 17555 41225
rect 17604 41228 21680 41256
rect 17218 41188 17224 41200
rect 16040 41160 17224 41188
rect 16040 41061 16068 41160
rect 17218 41148 17224 41160
rect 17276 41188 17282 41200
rect 17604 41188 17632 41228
rect 17276 41160 17632 41188
rect 20272 41160 20668 41188
rect 17276 41148 17282 41160
rect 16117 41123 16175 41129
rect 16117 41089 16129 41123
rect 16163 41120 16175 41123
rect 17865 41123 17923 41129
rect 16163 41092 16896 41120
rect 16163 41089 16175 41092
rect 16117 41083 16175 41089
rect 16868 41064 16896 41092
rect 17865 41089 17877 41123
rect 17911 41120 17923 41123
rect 18598 41120 18604 41132
rect 17911 41092 18604 41120
rect 17911 41089 17923 41092
rect 17865 41083 17923 41089
rect 18598 41080 18604 41092
rect 18656 41120 18662 41132
rect 18782 41120 18788 41132
rect 18656 41092 18788 41120
rect 18656 41080 18662 41092
rect 18782 41080 18788 41092
rect 18840 41080 18846 41132
rect 20272 41129 20300 41160
rect 20257 41123 20315 41129
rect 20257 41089 20269 41123
rect 20303 41089 20315 41123
rect 20257 41083 20315 41089
rect 20533 41123 20591 41129
rect 20533 41089 20545 41123
rect 20579 41089 20591 41123
rect 20640 41120 20668 41160
rect 21652 41132 21680 41228
rect 22002 41216 22008 41268
rect 22060 41256 22066 41268
rect 22465 41259 22523 41265
rect 22465 41256 22477 41259
rect 22060 41228 22477 41256
rect 22060 41216 22066 41228
rect 22465 41225 22477 41228
rect 22511 41225 22523 41259
rect 22465 41219 22523 41225
rect 23477 41259 23535 41265
rect 23477 41225 23489 41259
rect 23523 41256 23535 41259
rect 23566 41256 23572 41268
rect 23523 41228 23572 41256
rect 23523 41225 23535 41228
rect 23477 41219 23535 41225
rect 23566 41216 23572 41228
rect 23624 41216 23630 41268
rect 26142 41256 26148 41268
rect 25976 41228 26148 41256
rect 22066 41160 23704 41188
rect 21082 41120 21088 41132
rect 20640 41092 21088 41120
rect 20533 41083 20591 41089
rect 16025 41055 16083 41061
rect 16025 41021 16037 41055
rect 16071 41021 16083 41055
rect 16025 41015 16083 41021
rect 16850 41012 16856 41064
rect 16908 41012 16914 41064
rect 17770 41012 17776 41064
rect 17828 41052 17834 41064
rect 17957 41055 18015 41061
rect 17957 41052 17969 41055
rect 17828 41024 17969 41052
rect 17828 41012 17834 41024
rect 17957 41021 17969 41024
rect 18003 41021 18015 41055
rect 17957 41015 18015 41021
rect 18046 41012 18052 41064
rect 18104 41012 18110 41064
rect 20548 41052 20576 41083
rect 21082 41080 21088 41092
rect 21140 41080 21146 41132
rect 21177 41123 21235 41129
rect 21177 41089 21189 41123
rect 21223 41089 21235 41123
rect 21177 41083 21235 41089
rect 21269 41123 21327 41129
rect 21269 41089 21281 41123
rect 21315 41120 21327 41123
rect 21453 41123 21511 41129
rect 21315 41092 21404 41120
rect 21315 41089 21327 41092
rect 21269 41083 21327 41089
rect 21192 41052 21220 41083
rect 20548 41024 21312 41052
rect 21284 40996 21312 41024
rect 16485 40987 16543 40993
rect 16485 40953 16497 40987
rect 16531 40984 16543 40987
rect 18874 40984 18880 40996
rect 16531 40956 18880 40984
rect 16531 40953 16543 40956
rect 16485 40947 16543 40953
rect 18874 40944 18880 40956
rect 18932 40944 18938 40996
rect 20346 40944 20352 40996
rect 20404 40944 20410 40996
rect 20441 40987 20499 40993
rect 20441 40953 20453 40987
rect 20487 40984 20499 40987
rect 20530 40984 20536 40996
rect 20487 40956 20536 40984
rect 20487 40953 20499 40956
rect 20441 40947 20499 40953
rect 20530 40944 20536 40956
rect 20588 40944 20594 40996
rect 20806 40944 20812 40996
rect 20864 40944 20870 40996
rect 21266 40944 21272 40996
rect 21324 40944 21330 40996
rect 21376 40984 21404 41092
rect 21453 41089 21465 41123
rect 21499 41089 21511 41123
rect 21453 41083 21511 41089
rect 21468 41052 21496 41083
rect 21542 41080 21548 41132
rect 21600 41080 21606 41132
rect 21634 41080 21640 41132
rect 21692 41120 21698 41132
rect 22066 41120 22094 41160
rect 21692 41092 22094 41120
rect 22833 41123 22891 41129
rect 21692 41080 21698 41092
rect 22833 41089 22845 41123
rect 22879 41120 22891 41123
rect 23474 41120 23480 41132
rect 22879 41092 23480 41120
rect 22879 41089 22891 41092
rect 22833 41083 22891 41089
rect 23474 41080 23480 41092
rect 23532 41080 23538 41132
rect 23676 41129 23704 41160
rect 23842 41148 23848 41200
rect 23900 41148 23906 41200
rect 25976 41197 26004 41228
rect 26142 41216 26148 41228
rect 26200 41216 26206 41268
rect 26234 41216 26240 41268
rect 26292 41256 26298 41268
rect 27985 41259 28043 41265
rect 26292 41228 26464 41256
rect 26292 41216 26298 41228
rect 26436 41197 26464 41228
rect 27985 41225 27997 41259
rect 28031 41256 28043 41259
rect 28166 41256 28172 41268
rect 28031 41228 28172 41256
rect 28031 41225 28043 41228
rect 27985 41219 28043 41225
rect 28166 41216 28172 41228
rect 28224 41216 28230 41268
rect 28258 41216 28264 41268
rect 28316 41256 28322 41268
rect 28902 41256 28908 41268
rect 28316 41228 28908 41256
rect 28316 41216 28322 41228
rect 28902 41216 28908 41228
rect 28960 41216 28966 41268
rect 30834 41216 30840 41268
rect 30892 41256 30898 41268
rect 31478 41256 31484 41268
rect 30892 41228 31484 41256
rect 30892 41216 30898 41228
rect 31478 41216 31484 41228
rect 31536 41216 31542 41268
rect 33594 41216 33600 41268
rect 33652 41256 33658 41268
rect 34333 41259 34391 41265
rect 34333 41256 34345 41259
rect 33652 41228 34345 41256
rect 33652 41216 33658 41228
rect 34333 41225 34345 41228
rect 34379 41225 34391 41259
rect 34333 41219 34391 41225
rect 35158 41216 35164 41268
rect 35216 41216 35222 41268
rect 37645 41259 37703 41265
rect 37645 41225 37657 41259
rect 37691 41256 37703 41259
rect 37734 41256 37740 41268
rect 37691 41228 37740 41256
rect 37691 41225 37703 41228
rect 37645 41219 37703 41225
rect 37734 41216 37740 41228
rect 37792 41216 37798 41268
rect 39209 41259 39267 41265
rect 39209 41225 39221 41259
rect 39255 41256 39267 41259
rect 39390 41256 39396 41268
rect 39255 41228 39396 41256
rect 39255 41225 39267 41228
rect 39209 41219 39267 41225
rect 39390 41216 39396 41228
rect 39448 41216 39454 41268
rect 39482 41216 39488 41268
rect 39540 41256 39546 41268
rect 39577 41259 39635 41265
rect 39577 41256 39589 41259
rect 39540 41228 39589 41256
rect 39540 41216 39546 41228
rect 39577 41225 39589 41228
rect 39623 41225 39635 41259
rect 39577 41219 39635 41225
rect 25961 41191 26019 41197
rect 25961 41157 25973 41191
rect 26007 41157 26019 41191
rect 26421 41191 26479 41197
rect 26421 41188 26433 41191
rect 25961 41151 26019 41157
rect 26068 41160 26433 41188
rect 23661 41123 23719 41129
rect 23661 41089 23673 41123
rect 23707 41089 23719 41123
rect 23860 41120 23888 41148
rect 23937 41123 23995 41129
rect 23937 41120 23949 41123
rect 23860 41092 23949 41120
rect 23661 41083 23719 41089
rect 23937 41089 23949 41092
rect 23983 41089 23995 41123
rect 23937 41083 23995 41089
rect 24121 41123 24179 41129
rect 24121 41089 24133 41123
rect 24167 41120 24179 41123
rect 24762 41120 24768 41132
rect 24167 41092 24768 41120
rect 24167 41089 24179 41092
rect 24121 41083 24179 41089
rect 21910 41052 21916 41064
rect 21468 41024 21916 41052
rect 21910 41012 21916 41024
rect 21968 41012 21974 41064
rect 22738 41012 22744 41064
rect 22796 41052 22802 41064
rect 22925 41055 22983 41061
rect 22925 41052 22937 41055
rect 22796 41024 22937 41052
rect 22796 41012 22802 41024
rect 22925 41021 22937 41024
rect 22971 41021 22983 41055
rect 22925 41015 22983 41021
rect 23109 41055 23167 41061
rect 23109 41021 23121 41055
rect 23155 41052 23167 41055
rect 23566 41052 23572 41064
rect 23155 41024 23572 41052
rect 23155 41021 23167 41024
rect 23109 41015 23167 41021
rect 23566 41012 23572 41024
rect 23624 41012 23630 41064
rect 23676 41052 23704 41083
rect 24136 41052 24164 41083
rect 24762 41080 24768 41092
rect 24820 41080 24826 41132
rect 26068 41129 26096 41160
rect 26421 41157 26433 41160
rect 26467 41157 26479 41191
rect 29178 41188 29184 41200
rect 26421 41151 26479 41157
rect 28000 41160 29184 41188
rect 25777 41123 25835 41129
rect 25777 41089 25789 41123
rect 25823 41089 25835 41123
rect 25777 41083 25835 41089
rect 26053 41123 26111 41129
rect 26053 41089 26065 41123
rect 26099 41089 26111 41123
rect 26053 41083 26111 41089
rect 26145 41123 26203 41129
rect 26145 41089 26157 41123
rect 26191 41089 26203 41123
rect 26145 41083 26203 41089
rect 23676 41024 24164 41052
rect 21450 40984 21456 40996
rect 21376 40956 21456 40984
rect 21450 40944 21456 40956
rect 21508 40944 21514 40996
rect 22370 40944 22376 40996
rect 22428 40984 22434 40996
rect 24029 40987 24087 40993
rect 24029 40984 24041 40987
rect 22428 40956 24041 40984
rect 22428 40944 22434 40956
rect 24029 40953 24041 40956
rect 24075 40984 24087 40987
rect 24394 40984 24400 40996
rect 24075 40956 24400 40984
rect 24075 40953 24087 40956
rect 24029 40947 24087 40953
rect 24394 40944 24400 40956
rect 24452 40944 24458 40996
rect 25792 40984 25820 41083
rect 26160 40984 26188 41083
rect 26234 41080 26240 41132
rect 26292 41120 26298 41132
rect 26602 41120 26608 41132
rect 26292 41092 26608 41120
rect 26292 41080 26298 41092
rect 26602 41080 26608 41092
rect 26660 41080 26666 41132
rect 27798 41080 27804 41132
rect 27856 41080 27862 41132
rect 28000 41129 28028 41160
rect 29178 41148 29184 41160
rect 29236 41148 29242 41200
rect 31849 41191 31907 41197
rect 31849 41157 31861 41191
rect 31895 41188 31907 41191
rect 31895 41160 32352 41188
rect 31895 41157 31907 41160
rect 31849 41151 31907 41157
rect 27985 41123 28043 41129
rect 27985 41089 27997 41123
rect 28031 41089 28043 41123
rect 27985 41083 28043 41089
rect 28074 41080 28080 41132
rect 28132 41120 28138 41132
rect 28261 41123 28319 41129
rect 28261 41120 28273 41123
rect 28132 41092 28273 41120
rect 28132 41080 28138 41092
rect 28261 41089 28273 41092
rect 28307 41089 28319 41123
rect 28261 41083 28319 41089
rect 28534 41080 28540 41132
rect 28592 41080 28598 41132
rect 28721 41123 28779 41129
rect 28721 41089 28733 41123
rect 28767 41089 28779 41123
rect 28721 41083 28779 41089
rect 28350 41012 28356 41064
rect 28408 41012 28414 41064
rect 28445 41055 28503 41061
rect 28445 41021 28457 41055
rect 28491 41021 28503 41055
rect 28445 41015 28503 41021
rect 27062 40984 27068 40996
rect 25792 40956 27068 40984
rect 27062 40944 27068 40956
rect 27120 40944 27126 40996
rect 28077 40987 28135 40993
rect 28077 40953 28089 40987
rect 28123 40984 28135 40987
rect 28258 40984 28264 40996
rect 28123 40956 28264 40984
rect 28123 40953 28135 40956
rect 28077 40947 28135 40953
rect 28258 40944 28264 40956
rect 28316 40944 28322 40996
rect 28460 40928 28488 41015
rect 28736 40984 28764 41083
rect 28902 41080 28908 41132
rect 28960 41120 28966 41132
rect 28960 41080 28994 41120
rect 29086 41080 29092 41132
rect 29144 41120 29150 41132
rect 29730 41120 29736 41132
rect 29144 41092 29736 41120
rect 29144 41080 29150 41092
rect 29730 41080 29736 41092
rect 29788 41120 29794 41132
rect 30101 41123 30159 41129
rect 30101 41120 30113 41123
rect 29788 41092 30113 41120
rect 29788 41080 29794 41092
rect 30101 41089 30113 41092
rect 30147 41089 30159 41123
rect 30101 41083 30159 41089
rect 30926 41080 30932 41132
rect 30984 41080 30990 41132
rect 31570 41080 31576 41132
rect 31628 41080 31634 41132
rect 31754 41080 31760 41132
rect 31812 41080 31818 41132
rect 32324 41129 32352 41160
rect 32858 41148 32864 41200
rect 32916 41188 32922 41200
rect 34701 41191 34759 41197
rect 32916 41160 33548 41188
rect 32916 41148 32922 41160
rect 31941 41123 31999 41129
rect 31941 41089 31953 41123
rect 31987 41120 31999 41123
rect 32309 41123 32367 41129
rect 31987 41092 32260 41120
rect 31987 41089 31999 41092
rect 31941 41083 31999 41089
rect 28966 41052 28994 41080
rect 28966 41024 31754 41052
rect 31110 40984 31116 40996
rect 28736 40956 31116 40984
rect 31110 40944 31116 40956
rect 31168 40944 31174 40996
rect 31726 40984 31754 41024
rect 32232 40984 32260 41092
rect 32309 41089 32321 41123
rect 32355 41089 32367 41123
rect 32309 41083 32367 41089
rect 33134 41080 33140 41132
rect 33192 41080 33198 41132
rect 33226 41080 33232 41132
rect 33284 41120 33290 41132
rect 33321 41123 33379 41129
rect 33321 41120 33333 41123
rect 33284 41092 33333 41120
rect 33284 41080 33290 41092
rect 33321 41089 33333 41092
rect 33367 41089 33379 41123
rect 33321 41083 33379 41089
rect 33410 41080 33416 41132
rect 33468 41080 33474 41132
rect 33520 41129 33548 41160
rect 34701 41157 34713 41191
rect 34747 41188 34759 41191
rect 34790 41188 34796 41200
rect 34747 41160 34796 41188
rect 34747 41157 34759 41160
rect 34701 41151 34759 41157
rect 34790 41148 34796 41160
rect 34848 41188 34854 41200
rect 35621 41191 35679 41197
rect 35621 41188 35633 41191
rect 34848 41160 35633 41188
rect 34848 41148 34854 41160
rect 35621 41157 35633 41160
rect 35667 41157 35679 41191
rect 35621 41151 35679 41157
rect 36817 41191 36875 41197
rect 36817 41157 36829 41191
rect 36863 41188 36875 41191
rect 37366 41188 37372 41200
rect 36863 41160 37372 41188
rect 36863 41157 36875 41160
rect 36817 41151 36875 41157
rect 37366 41148 37372 41160
rect 37424 41188 37430 41200
rect 37550 41188 37556 41200
rect 37424 41160 37556 41188
rect 37424 41148 37430 41160
rect 37550 41148 37556 41160
rect 37608 41148 37614 41200
rect 37826 41148 37832 41200
rect 37884 41148 37890 41200
rect 37918 41148 37924 41200
rect 37976 41188 37982 41200
rect 38562 41188 38568 41200
rect 37976 41160 38568 41188
rect 37976 41148 37982 41160
rect 33505 41123 33563 41129
rect 33505 41089 33517 41123
rect 33551 41089 33563 41123
rect 33505 41083 33563 41089
rect 33597 41123 33655 41129
rect 33597 41089 33609 41123
rect 33643 41120 33655 41123
rect 35434 41120 35440 41132
rect 33643 41092 33677 41120
rect 34808 41092 35440 41120
rect 33643 41089 33655 41092
rect 33597 41083 33655 41089
rect 32401 41055 32459 41061
rect 32401 41021 32413 41055
rect 32447 41052 32459 41055
rect 33042 41052 33048 41064
rect 32447 41024 33048 41052
rect 32447 41021 32459 41024
rect 32401 41015 32459 41021
rect 33042 41012 33048 41024
rect 33100 41012 33106 41064
rect 33428 41052 33456 41080
rect 33612 41052 33640 41083
rect 34422 41052 34428 41064
rect 33428 41024 34428 41052
rect 34422 41012 34428 41024
rect 34480 41012 34486 41064
rect 34808 41061 34836 41092
rect 35434 41080 35440 41092
rect 35492 41120 35498 41132
rect 35529 41123 35587 41129
rect 35529 41120 35541 41123
rect 35492 41092 35541 41120
rect 35492 41080 35498 41092
rect 35529 41089 35541 41092
rect 35575 41089 35587 41123
rect 35529 41083 35587 41089
rect 37001 41123 37059 41129
rect 37001 41089 37013 41123
rect 37047 41089 37059 41123
rect 37001 41083 37059 41089
rect 37093 41123 37151 41129
rect 37093 41089 37105 41123
rect 37139 41120 37151 41123
rect 37844 41120 37872 41148
rect 38120 41129 38148 41160
rect 38562 41148 38568 41160
rect 38620 41188 38626 41200
rect 40037 41191 40095 41197
rect 40037 41188 40049 41191
rect 38620 41160 40049 41188
rect 38620 41148 38626 41160
rect 40037 41157 40049 41160
rect 40083 41157 40095 41191
rect 40037 41151 40095 41157
rect 38105 41123 38163 41129
rect 37139 41092 37964 41120
rect 37139 41089 37151 41092
rect 37093 41083 37151 41089
rect 34793 41055 34851 41061
rect 34793 41021 34805 41055
rect 34839 41021 34851 41055
rect 34793 41015 34851 41021
rect 34885 41055 34943 41061
rect 34885 41021 34897 41055
rect 34931 41021 34943 41055
rect 34885 41015 34943 41021
rect 35713 41055 35771 41061
rect 35713 41021 35725 41055
rect 35759 41021 35771 41055
rect 35713 41015 35771 41021
rect 33318 40984 33324 40996
rect 31726 40956 33324 40984
rect 33318 40944 33324 40956
rect 33376 40984 33382 40996
rect 33413 40987 33471 40993
rect 33413 40984 33425 40987
rect 33376 40956 33425 40984
rect 33376 40944 33382 40956
rect 33413 40953 33425 40956
rect 33459 40953 33471 40987
rect 33413 40947 33471 40953
rect 34698 40944 34704 40996
rect 34756 40984 34762 40996
rect 34900 40984 34928 41015
rect 35728 40984 35756 41015
rect 37016 40984 37044 41083
rect 37737 41055 37795 41061
rect 37737 41021 37749 41055
rect 37783 41021 37795 41055
rect 37737 41015 37795 41021
rect 37752 40984 37780 41015
rect 37826 41012 37832 41064
rect 37884 41012 37890 41064
rect 37936 41052 37964 41092
rect 38105 41089 38117 41123
rect 38151 41089 38163 41123
rect 38105 41083 38163 41089
rect 38286 41080 38292 41132
rect 38344 41080 38350 41132
rect 38749 41123 38807 41129
rect 38749 41089 38761 41123
rect 38795 41120 38807 41123
rect 39574 41120 39580 41132
rect 38795 41092 39580 41120
rect 38795 41089 38807 41092
rect 38749 41083 38807 41089
rect 39574 41080 39580 41092
rect 39632 41080 39638 41132
rect 40218 41080 40224 41132
rect 40276 41080 40282 41132
rect 38197 41055 38255 41061
rect 38197 41052 38209 41055
rect 37936 41024 38209 41052
rect 38197 41021 38209 41024
rect 38243 41021 38255 41055
rect 38197 41015 38255 41021
rect 38838 41012 38844 41064
rect 38896 41012 38902 41064
rect 39025 41055 39083 41061
rect 39025 41021 39037 41055
rect 39071 41021 39083 41055
rect 39025 41015 39083 41021
rect 38381 40987 38439 40993
rect 38381 40984 38393 40987
rect 34756 40956 35756 40984
rect 36740 40956 36952 40984
rect 37016 40956 37412 40984
rect 37752 40956 38393 40984
rect 34756 40944 34762 40956
rect 17034 40876 17040 40928
rect 17092 40916 17098 40928
rect 17405 40919 17463 40925
rect 17405 40916 17417 40919
rect 17092 40888 17417 40916
rect 17092 40876 17098 40888
rect 17405 40885 17417 40888
rect 17451 40885 17463 40919
rect 17405 40879 17463 40885
rect 20717 40919 20775 40925
rect 20717 40885 20729 40919
rect 20763 40916 20775 40919
rect 21174 40916 21180 40928
rect 20763 40888 21180 40916
rect 20763 40885 20775 40888
rect 20717 40879 20775 40885
rect 21174 40876 21180 40888
rect 21232 40876 21238 40928
rect 26050 40876 26056 40928
rect 26108 40876 26114 40928
rect 26418 40876 26424 40928
rect 26476 40876 26482 40928
rect 28442 40876 28448 40928
rect 28500 40876 28506 40928
rect 28626 40876 28632 40928
rect 28684 40916 28690 40928
rect 29270 40916 29276 40928
rect 28684 40888 29276 40916
rect 28684 40876 28690 40888
rect 29270 40876 29276 40888
rect 29328 40876 29334 40928
rect 30466 40876 30472 40928
rect 30524 40916 30530 40928
rect 31021 40919 31079 40925
rect 31021 40916 31033 40919
rect 30524 40888 31033 40916
rect 30524 40876 30530 40888
rect 31021 40885 31033 40888
rect 31067 40885 31079 40919
rect 31021 40879 31079 40885
rect 32582 40876 32588 40928
rect 32640 40876 32646 40928
rect 33781 40919 33839 40925
rect 33781 40885 33793 40919
rect 33827 40916 33839 40919
rect 36740 40916 36768 40956
rect 33827 40888 36768 40916
rect 33827 40885 33839 40888
rect 33781 40879 33839 40885
rect 36814 40876 36820 40928
rect 36872 40876 36878 40928
rect 36924 40916 36952 40956
rect 37182 40916 37188 40928
rect 36924 40888 37188 40916
rect 37182 40876 37188 40888
rect 37240 40876 37246 40928
rect 37274 40876 37280 40928
rect 37332 40876 37338 40928
rect 37384 40916 37412 40956
rect 38381 40953 38393 40956
rect 38427 40953 38439 40987
rect 39040 40984 39068 41015
rect 39298 41012 39304 41064
rect 39356 41052 39362 41064
rect 39669 41055 39727 41061
rect 39669 41052 39681 41055
rect 39356 41024 39681 41052
rect 39356 41012 39362 41024
rect 39669 41021 39681 41024
rect 39715 41021 39727 41055
rect 39669 41015 39727 41021
rect 39761 41055 39819 41061
rect 39761 41021 39773 41055
rect 39807 41052 39819 41055
rect 40126 41052 40132 41064
rect 39807 41024 40132 41052
rect 39807 41021 39819 41024
rect 39761 41015 39819 41021
rect 40126 41012 40132 41024
rect 40184 41012 40190 41064
rect 39850 40984 39856 40996
rect 39040 40956 39856 40984
rect 38381 40947 38439 40953
rect 39850 40944 39856 40956
rect 39908 40944 39914 40996
rect 37642 40916 37648 40928
rect 37384 40888 37648 40916
rect 37642 40876 37648 40888
rect 37700 40916 37706 40928
rect 40405 40919 40463 40925
rect 40405 40916 40417 40919
rect 37700 40888 40417 40916
rect 37700 40876 37706 40888
rect 40405 40885 40417 40888
rect 40451 40885 40463 40919
rect 40405 40879 40463 40885
rect 1104 40826 42504 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 42504 40826
rect 1104 40752 42504 40774
rect 16850 40672 16856 40724
rect 16908 40712 16914 40724
rect 17129 40715 17187 40721
rect 17129 40712 17141 40715
rect 16908 40684 17141 40712
rect 16908 40672 16914 40684
rect 17129 40681 17141 40684
rect 17175 40681 17187 40715
rect 17129 40675 17187 40681
rect 17770 40672 17776 40724
rect 17828 40672 17834 40724
rect 18601 40715 18659 40721
rect 18601 40681 18613 40715
rect 18647 40712 18659 40715
rect 20346 40712 20352 40724
rect 18647 40684 20352 40712
rect 18647 40681 18659 40684
rect 18601 40675 18659 40681
rect 20346 40672 20352 40684
rect 20404 40672 20410 40724
rect 24949 40715 25007 40721
rect 24949 40681 24961 40715
rect 24995 40712 25007 40715
rect 24995 40684 27660 40712
rect 24995 40681 25007 40684
rect 24949 40675 25007 40681
rect 19429 40647 19487 40653
rect 19429 40613 19441 40647
rect 19475 40644 19487 40647
rect 20530 40644 20536 40656
rect 19475 40616 20536 40644
rect 19475 40613 19487 40616
rect 19429 40607 19487 40613
rect 20530 40604 20536 40616
rect 20588 40644 20594 40656
rect 21177 40647 21235 40653
rect 21177 40644 21189 40647
rect 20588 40616 21189 40644
rect 20588 40604 20594 40616
rect 21177 40613 21189 40616
rect 21223 40613 21235 40647
rect 21177 40607 21235 40613
rect 26050 40604 26056 40656
rect 26108 40604 26114 40656
rect 17402 40536 17408 40588
rect 17460 40576 17466 40588
rect 18325 40579 18383 40585
rect 18325 40576 18337 40579
rect 17460 40548 18337 40576
rect 17460 40536 17466 40548
rect 18325 40545 18337 40548
rect 18371 40545 18383 40579
rect 18325 40539 18383 40545
rect 14734 40468 14740 40520
rect 14792 40508 14798 40520
rect 15381 40511 15439 40517
rect 15381 40508 15393 40511
rect 14792 40480 15393 40508
rect 14792 40468 14798 40480
rect 15381 40477 15393 40480
rect 15427 40477 15439 40511
rect 15381 40471 15439 40477
rect 18782 40468 18788 40520
rect 18840 40468 18846 40520
rect 18874 40468 18880 40520
rect 18932 40468 18938 40520
rect 20548 40517 20576 40604
rect 21085 40579 21143 40585
rect 21085 40576 21097 40579
rect 20732 40548 21097 40576
rect 20732 40517 20760 40548
rect 21085 40545 21097 40548
rect 21131 40545 21143 40579
rect 21085 40539 21143 40545
rect 21453 40579 21511 40585
rect 21453 40545 21465 40579
rect 21499 40576 21511 40579
rect 24854 40576 24860 40588
rect 21499 40548 24860 40576
rect 21499 40545 21511 40548
rect 21453 40539 21511 40545
rect 24854 40536 24860 40548
rect 24912 40576 24918 40588
rect 25317 40579 25375 40585
rect 25317 40576 25329 40579
rect 24912 40548 25329 40576
rect 24912 40536 24918 40548
rect 25317 40545 25329 40548
rect 25363 40545 25375 40579
rect 25317 40539 25375 40545
rect 19245 40511 19303 40517
rect 19245 40477 19257 40511
rect 19291 40477 19303 40511
rect 19429 40511 19487 40517
rect 19429 40508 19441 40511
rect 19245 40471 19303 40477
rect 19352 40480 19441 40508
rect 15654 40400 15660 40452
rect 15712 40400 15718 40452
rect 16114 40400 16120 40452
rect 16172 40400 16178 40452
rect 18601 40443 18659 40449
rect 18601 40409 18613 40443
rect 18647 40440 18659 40443
rect 18690 40440 18696 40452
rect 18647 40412 18696 40440
rect 18647 40409 18659 40412
rect 18601 40403 18659 40409
rect 18690 40400 18696 40412
rect 18748 40400 18754 40452
rect 18800 40440 18828 40468
rect 19260 40440 19288 40471
rect 18800 40412 19288 40440
rect 17770 40332 17776 40384
rect 17828 40372 17834 40384
rect 18141 40375 18199 40381
rect 18141 40372 18153 40375
rect 17828 40344 18153 40372
rect 17828 40332 17834 40344
rect 18141 40341 18153 40344
rect 18187 40341 18199 40375
rect 18141 40335 18199 40341
rect 18230 40332 18236 40384
rect 18288 40332 18294 40384
rect 18874 40332 18880 40384
rect 18932 40372 18938 40384
rect 19352 40372 19380 40480
rect 19429 40477 19441 40480
rect 19475 40477 19487 40511
rect 19429 40471 19487 40477
rect 20533 40511 20591 40517
rect 20533 40477 20545 40511
rect 20579 40477 20591 40511
rect 20533 40471 20591 40477
rect 20717 40511 20775 40517
rect 20717 40477 20729 40511
rect 20763 40477 20775 40511
rect 20717 40471 20775 40477
rect 20809 40511 20867 40517
rect 20809 40477 20821 40511
rect 20855 40477 20867 40511
rect 20809 40471 20867 40477
rect 19518 40400 19524 40452
rect 19576 40400 19582 40452
rect 20257 40443 20315 40449
rect 20257 40409 20269 40443
rect 20303 40409 20315 40443
rect 20257 40403 20315 40409
rect 18932 40344 19380 40372
rect 18932 40332 18938 40344
rect 19426 40332 19432 40384
rect 19484 40372 19490 40384
rect 20272 40372 20300 40403
rect 20346 40400 20352 40452
rect 20404 40440 20410 40452
rect 20732 40440 20760 40471
rect 20404 40412 20760 40440
rect 20824 40440 20852 40471
rect 20990 40468 20996 40520
rect 21048 40468 21054 40520
rect 21266 40468 21272 40520
rect 21324 40468 21330 40520
rect 22554 40508 22560 40520
rect 22066 40480 22560 40508
rect 22066 40440 22094 40480
rect 22554 40468 22560 40480
rect 22612 40508 22618 40520
rect 22771 40511 22829 40517
rect 22771 40508 22783 40511
rect 22612 40480 22783 40508
rect 22612 40468 22618 40480
rect 22771 40477 22783 40480
rect 22817 40477 22829 40511
rect 22771 40471 22829 40477
rect 22925 40511 22983 40517
rect 22925 40477 22937 40511
rect 22971 40508 22983 40511
rect 24578 40508 24584 40520
rect 22971 40480 24584 40508
rect 22971 40477 22983 40480
rect 22925 40471 22983 40477
rect 24578 40468 24584 40480
rect 24636 40468 24642 40520
rect 25130 40468 25136 40520
rect 25188 40468 25194 40520
rect 25225 40511 25283 40517
rect 25225 40477 25237 40511
rect 25271 40477 25283 40511
rect 25225 40471 25283 40477
rect 20824 40412 22094 40440
rect 24596 40440 24624 40468
rect 25240 40440 25268 40471
rect 25406 40468 25412 40520
rect 25464 40468 25470 40520
rect 25593 40511 25651 40517
rect 25593 40477 25605 40511
rect 25639 40508 25651 40511
rect 26068 40508 26096 40604
rect 25639 40480 26096 40508
rect 25639 40477 25651 40480
rect 25593 40471 25651 40477
rect 26418 40468 26424 40520
rect 26476 40508 26482 40520
rect 27632 40517 27660 40684
rect 27890 40672 27896 40724
rect 27948 40712 27954 40724
rect 28166 40712 28172 40724
rect 27948 40684 28172 40712
rect 27948 40672 27954 40684
rect 28166 40672 28172 40684
rect 28224 40672 28230 40724
rect 28644 40684 28856 40712
rect 28644 40644 28672 40684
rect 28460 40616 28672 40644
rect 28460 40585 28488 40616
rect 28718 40604 28724 40656
rect 28776 40604 28782 40656
rect 28828 40644 28856 40684
rect 30006 40672 30012 40724
rect 30064 40712 30070 40724
rect 30101 40715 30159 40721
rect 30101 40712 30113 40715
rect 30064 40684 30113 40712
rect 30064 40672 30070 40684
rect 30101 40681 30113 40684
rect 30147 40681 30159 40715
rect 30101 40675 30159 40681
rect 31478 40672 31484 40724
rect 31536 40712 31542 40724
rect 34698 40712 34704 40724
rect 31536 40684 34704 40712
rect 31536 40672 31542 40684
rect 34698 40672 34704 40684
rect 34756 40672 34762 40724
rect 36252 40715 36310 40721
rect 36252 40681 36264 40715
rect 36298 40712 36310 40715
rect 37274 40712 37280 40724
rect 36298 40684 37280 40712
rect 36298 40681 36310 40684
rect 36252 40675 36310 40681
rect 37274 40672 37280 40684
rect 37332 40672 37338 40724
rect 37366 40672 37372 40724
rect 37424 40712 37430 40724
rect 37737 40715 37795 40721
rect 37737 40712 37749 40715
rect 37424 40684 37749 40712
rect 37424 40672 37430 40684
rect 37737 40681 37749 40684
rect 37783 40681 37795 40715
rect 37737 40675 37795 40681
rect 38286 40672 38292 40724
rect 38344 40712 38350 40724
rect 40034 40712 40040 40724
rect 38344 40684 40040 40712
rect 38344 40672 38350 40684
rect 40034 40672 40040 40684
rect 40092 40712 40098 40724
rect 40218 40712 40224 40724
rect 40092 40684 40224 40712
rect 40092 40672 40098 40684
rect 40218 40672 40224 40684
rect 40276 40672 40282 40724
rect 31021 40647 31079 40653
rect 31021 40644 31033 40647
rect 28828 40616 31033 40644
rect 31021 40613 31033 40616
rect 31067 40613 31079 40647
rect 31021 40607 31079 40613
rect 31110 40604 31116 40656
rect 31168 40604 31174 40656
rect 33042 40604 33048 40656
rect 33100 40604 33106 40656
rect 38010 40604 38016 40656
rect 38068 40644 38074 40656
rect 40126 40644 40132 40656
rect 38068 40616 40132 40644
rect 38068 40604 38074 40616
rect 40126 40604 40132 40616
rect 40184 40604 40190 40656
rect 28445 40579 28503 40585
rect 28445 40545 28457 40579
rect 28491 40545 28503 40579
rect 28445 40539 28503 40545
rect 28534 40536 28540 40588
rect 28592 40576 28598 40588
rect 28592 40548 29316 40576
rect 28592 40536 28598 40548
rect 27433 40511 27491 40517
rect 27433 40508 27445 40511
rect 26476 40480 27445 40508
rect 26476 40468 26482 40480
rect 27433 40477 27445 40480
rect 27479 40477 27491 40511
rect 27433 40471 27491 40477
rect 27617 40511 27675 40517
rect 27617 40477 27629 40511
rect 27663 40508 27675 40511
rect 27798 40508 27804 40520
rect 27663 40480 27804 40508
rect 27663 40477 27675 40480
rect 27617 40471 27675 40477
rect 24596 40412 25268 40440
rect 27448 40440 27476 40471
rect 27798 40468 27804 40480
rect 27856 40468 27862 40520
rect 27982 40508 27988 40520
rect 27943 40480 27988 40508
rect 27982 40468 27988 40480
rect 28040 40468 28046 40520
rect 28074 40468 28080 40520
rect 28132 40468 28138 40520
rect 28353 40511 28411 40517
rect 28353 40477 28365 40511
rect 28399 40508 28411 40511
rect 28813 40511 28871 40517
rect 28813 40508 28825 40511
rect 28399 40480 28825 40508
rect 28399 40477 28411 40480
rect 28353 40471 28411 40477
rect 28813 40477 28825 40480
rect 28859 40477 28871 40511
rect 28813 40471 28871 40477
rect 28902 40468 28908 40520
rect 28960 40508 28966 40520
rect 29288 40517 29316 40548
rect 30650 40536 30656 40588
rect 30708 40536 30714 40588
rect 31481 40579 31539 40585
rect 31481 40545 31493 40579
rect 31527 40576 31539 40579
rect 31754 40576 31760 40588
rect 31527 40548 31760 40576
rect 31527 40545 31539 40548
rect 31481 40539 31539 40545
rect 31754 40536 31760 40548
rect 31812 40536 31818 40588
rect 32858 40536 32864 40588
rect 32916 40536 32922 40588
rect 35986 40536 35992 40588
rect 36044 40576 36050 40588
rect 36044 40548 39252 40576
rect 36044 40536 36050 40548
rect 39224 40520 39252 40548
rect 28997 40511 29055 40517
rect 28997 40508 29009 40511
rect 28960 40480 29009 40508
rect 28960 40468 28966 40480
rect 28997 40477 29009 40480
rect 29043 40477 29055 40511
rect 28997 40471 29055 40477
rect 29089 40511 29147 40517
rect 29089 40477 29101 40511
rect 29135 40477 29147 40511
rect 29089 40471 29147 40477
rect 29181 40511 29239 40517
rect 29181 40477 29193 40511
rect 29227 40477 29239 40511
rect 29181 40471 29239 40477
rect 29273 40511 29331 40517
rect 29273 40477 29285 40511
rect 29319 40477 29331 40511
rect 29273 40471 29331 40477
rect 29104 40440 29132 40471
rect 27448 40412 29132 40440
rect 20404 40400 20410 40412
rect 28368 40384 28396 40412
rect 19484 40344 20300 40372
rect 20625 40375 20683 40381
rect 19484 40332 19490 40344
rect 20625 40341 20637 40375
rect 20671 40372 20683 40375
rect 20714 40372 20720 40384
rect 20671 40344 20720 40372
rect 20671 40341 20683 40344
rect 20625 40335 20683 40341
rect 20714 40332 20720 40344
rect 20772 40332 20778 40384
rect 22554 40332 22560 40384
rect 22612 40332 22618 40384
rect 25961 40375 26019 40381
rect 25961 40341 25973 40375
rect 26007 40372 26019 40375
rect 26050 40372 26056 40384
rect 26007 40344 26056 40372
rect 26007 40341 26019 40344
rect 25961 40335 26019 40341
rect 26050 40332 26056 40344
rect 26108 40332 26114 40384
rect 27525 40375 27583 40381
rect 27525 40341 27537 40375
rect 27571 40372 27583 40375
rect 27614 40372 27620 40384
rect 27571 40344 27620 40372
rect 27571 40341 27583 40344
rect 27525 40335 27583 40341
rect 27614 40332 27620 40344
rect 27672 40332 27678 40384
rect 27709 40375 27767 40381
rect 27709 40341 27721 40375
rect 27755 40372 27767 40375
rect 27890 40372 27896 40384
rect 27755 40344 27896 40372
rect 27755 40341 27767 40344
rect 27709 40335 27767 40341
rect 27890 40332 27896 40344
rect 27948 40332 27954 40384
rect 28350 40332 28356 40384
rect 28408 40332 28414 40384
rect 28902 40332 28908 40384
rect 28960 40372 28966 40384
rect 29196 40372 29224 40471
rect 30466 40468 30472 40520
rect 30524 40468 30530 40520
rect 32766 40468 32772 40520
rect 32824 40468 32830 40520
rect 33226 40468 33232 40520
rect 33284 40517 33290 40520
rect 33284 40511 33317 40517
rect 33305 40477 33317 40511
rect 33284 40471 33317 40477
rect 33284 40468 33290 40471
rect 33410 40468 33416 40520
rect 33468 40468 33474 40520
rect 39206 40468 39212 40520
rect 39264 40468 39270 40520
rect 38102 40440 38108 40452
rect 37490 40412 38108 40440
rect 38102 40400 38108 40412
rect 38160 40440 38166 40452
rect 40126 40440 40132 40452
rect 38160 40412 40132 40440
rect 38160 40400 38166 40412
rect 40126 40400 40132 40412
rect 40184 40400 40190 40452
rect 28960 40344 29224 40372
rect 28960 40332 28966 40344
rect 30558 40332 30564 40384
rect 30616 40332 30622 40384
rect 32398 40332 32404 40384
rect 32456 40332 32462 40384
rect 1104 40282 42504 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 35594 40282
rect 35646 40230 35658 40282
rect 35710 40230 35722 40282
rect 35774 40230 35786 40282
rect 35838 40230 35850 40282
rect 35902 40230 42504 40282
rect 1104 40208 42504 40230
rect 15654 40128 15660 40180
rect 15712 40168 15718 40180
rect 16669 40171 16727 40177
rect 16669 40168 16681 40171
rect 15712 40140 16681 40168
rect 15712 40128 15718 40140
rect 16669 40137 16681 40140
rect 16715 40137 16727 40171
rect 16669 40131 16727 40137
rect 17034 40128 17040 40180
rect 17092 40128 17098 40180
rect 17129 40171 17187 40177
rect 17129 40137 17141 40171
rect 17175 40168 17187 40171
rect 17497 40171 17555 40177
rect 17497 40168 17509 40171
rect 17175 40140 17509 40168
rect 17175 40137 17187 40140
rect 17129 40131 17187 40137
rect 17497 40137 17509 40140
rect 17543 40137 17555 40171
rect 17497 40131 17555 40137
rect 17865 40171 17923 40177
rect 17865 40137 17877 40171
rect 17911 40168 17923 40171
rect 18230 40168 18236 40180
rect 17911 40140 18236 40168
rect 17911 40137 17923 40140
rect 17865 40131 17923 40137
rect 18230 40128 18236 40140
rect 18288 40128 18294 40180
rect 23293 40171 23351 40177
rect 23293 40137 23305 40171
rect 23339 40168 23351 40171
rect 24394 40168 24400 40180
rect 23339 40140 24400 40168
rect 23339 40137 23351 40140
rect 23293 40131 23351 40137
rect 24394 40128 24400 40140
rect 24452 40128 24458 40180
rect 27982 40128 27988 40180
rect 28040 40168 28046 40180
rect 28534 40168 28540 40180
rect 28040 40140 28540 40168
rect 28040 40128 28046 40140
rect 28534 40128 28540 40140
rect 28592 40128 28598 40180
rect 32858 40128 32864 40180
rect 32916 40168 32922 40180
rect 36449 40171 36507 40177
rect 36449 40168 36461 40171
rect 32916 40140 36461 40168
rect 32916 40128 32922 40140
rect 36449 40137 36461 40140
rect 36495 40137 36507 40171
rect 36449 40131 36507 40137
rect 39298 40128 39304 40180
rect 39356 40128 39362 40180
rect 39574 40128 39580 40180
rect 39632 40168 39638 40180
rect 39761 40171 39819 40177
rect 39761 40168 39773 40171
rect 39632 40140 39773 40168
rect 39632 40128 39638 40140
rect 39761 40137 39773 40140
rect 39807 40137 39819 40171
rect 39761 40131 39819 40137
rect 17770 40060 17776 40112
rect 17828 40100 17834 40112
rect 17957 40103 18015 40109
rect 17957 40100 17969 40103
rect 17828 40072 17969 40100
rect 17828 40060 17834 40072
rect 17957 40069 17969 40072
rect 18003 40069 18015 40103
rect 18782 40100 18788 40112
rect 17957 40063 18015 40069
rect 18524 40072 18788 40100
rect 18524 40041 18552 40072
rect 18782 40060 18788 40072
rect 18840 40060 18846 40112
rect 21174 40060 21180 40112
rect 21232 40100 21238 40112
rect 21232 40072 22048 40100
rect 21232 40060 21238 40072
rect 18509 40035 18567 40041
rect 18509 40001 18521 40035
rect 18555 40001 18567 40035
rect 18509 39995 18567 40001
rect 19426 39992 19432 40044
rect 19484 40032 19490 40044
rect 19613 40035 19671 40041
rect 19613 40032 19625 40035
rect 19484 40004 19625 40032
rect 19484 39992 19490 40004
rect 19613 40001 19625 40004
rect 19659 40001 19671 40035
rect 19613 39995 19671 40001
rect 20714 39992 20720 40044
rect 20772 39992 20778 40044
rect 22020 40041 22048 40072
rect 23382 40060 23388 40112
rect 23440 40060 23446 40112
rect 24872 40072 25176 40100
rect 24872 40044 24900 40072
rect 22005 40035 22063 40041
rect 22005 40001 22017 40035
rect 22051 40001 22063 40035
rect 22005 39995 22063 40001
rect 22094 39992 22100 40044
rect 22152 40032 22158 40044
rect 22925 40035 22983 40041
rect 22925 40032 22937 40035
rect 22152 40004 22937 40032
rect 22152 39992 22158 40004
rect 22925 40001 22937 40004
rect 22971 40001 22983 40035
rect 22925 39995 22983 40001
rect 24213 40035 24271 40041
rect 24213 40001 24225 40035
rect 24259 40032 24271 40035
rect 24302 40032 24308 40044
rect 24259 40004 24308 40032
rect 24259 40001 24271 40004
rect 24213 39995 24271 40001
rect 24302 39992 24308 40004
rect 24360 39992 24366 40044
rect 24578 39992 24584 40044
rect 24636 39992 24642 40044
rect 24765 40035 24823 40041
rect 24765 40001 24777 40035
rect 24811 40032 24823 40035
rect 24854 40032 24860 40044
rect 24811 40004 24860 40032
rect 24811 40001 24823 40004
rect 24765 39995 24823 40001
rect 24854 39992 24860 40004
rect 24912 39992 24918 40044
rect 25148 40041 25176 40072
rect 27614 40060 27620 40112
rect 27672 40100 27678 40112
rect 27672 40072 28028 40100
rect 27672 40060 27678 40072
rect 25041 40035 25099 40041
rect 25041 40001 25053 40035
rect 25087 40001 25099 40035
rect 25041 39995 25099 40001
rect 25133 40035 25191 40041
rect 25133 40001 25145 40035
rect 25179 40001 25191 40035
rect 25133 39995 25191 40001
rect 17310 39924 17316 39976
rect 17368 39964 17374 39976
rect 17862 39964 17868 39976
rect 17368 39936 17868 39964
rect 17368 39924 17374 39936
rect 17862 39924 17868 39936
rect 17920 39924 17926 39976
rect 18049 39967 18107 39973
rect 18049 39933 18061 39967
rect 18095 39933 18107 39967
rect 18049 39927 18107 39933
rect 18601 39967 18659 39973
rect 18601 39933 18613 39967
rect 18647 39964 18659 39967
rect 18874 39964 18880 39976
rect 18647 39936 18880 39964
rect 18647 39933 18659 39936
rect 18601 39927 18659 39933
rect 17402 39856 17408 39908
rect 17460 39896 17466 39908
rect 18064 39896 18092 39927
rect 18874 39924 18880 39936
rect 18932 39924 18938 39976
rect 20806 39924 20812 39976
rect 20864 39924 20870 39976
rect 21913 39967 21971 39973
rect 21913 39933 21925 39967
rect 21959 39964 21971 39967
rect 22554 39964 22560 39976
rect 21959 39936 22560 39964
rect 21959 39933 21971 39936
rect 21913 39927 21971 39933
rect 22554 39924 22560 39936
rect 22612 39924 22618 39976
rect 23014 39924 23020 39976
rect 23072 39924 23078 39976
rect 17460 39868 18092 39896
rect 17460 39856 17466 39868
rect 21082 39856 21088 39908
rect 21140 39896 21146 39908
rect 24596 39896 24624 39992
rect 25056 39964 25084 39995
rect 25222 39992 25228 40044
rect 25280 40032 25286 40044
rect 28000 40041 28028 40072
rect 32398 40060 32404 40112
rect 32456 40060 32462 40112
rect 33134 40060 33140 40112
rect 33192 40100 33198 40112
rect 33192 40072 36584 40100
rect 33192 40060 33198 40072
rect 25317 40035 25375 40041
rect 25317 40032 25329 40035
rect 25280 40004 25329 40032
rect 25280 39992 25286 40004
rect 25317 40001 25329 40004
rect 25363 40001 25375 40035
rect 25317 39995 25375 40001
rect 25501 40035 25559 40041
rect 25501 40001 25513 40035
rect 25547 40032 25559 40035
rect 25961 40035 26019 40041
rect 25961 40032 25973 40035
rect 25547 40004 25973 40032
rect 25547 40001 25559 40004
rect 25501 39995 25559 40001
rect 25961 40001 25973 40004
rect 26007 40001 26019 40035
rect 25961 39995 26019 40001
rect 27985 40035 28043 40041
rect 27985 40001 27997 40035
rect 28031 40001 28043 40035
rect 27985 39995 28043 40001
rect 31021 40035 31079 40041
rect 31021 40001 31033 40035
rect 31067 40032 31079 40035
rect 31110 40032 31116 40044
rect 31067 40004 31116 40032
rect 31067 40001 31079 40004
rect 31021 39995 31079 40001
rect 31110 39992 31116 40004
rect 31168 39992 31174 40044
rect 32030 39992 32036 40044
rect 32088 40032 32094 40044
rect 32125 40035 32183 40041
rect 32125 40032 32137 40035
rect 32088 40004 32137 40032
rect 32088 39992 32094 40004
rect 32125 40001 32137 40004
rect 32171 40001 32183 40035
rect 32125 39995 32183 40001
rect 32217 40035 32275 40041
rect 32217 40001 32229 40035
rect 32263 40001 32275 40035
rect 32217 39995 32275 40001
rect 36556 40032 36584 40072
rect 36814 40060 36820 40112
rect 36872 40100 36878 40112
rect 36909 40103 36967 40109
rect 36909 40100 36921 40103
rect 36872 40072 36921 40100
rect 36872 40060 36878 40072
rect 36909 40069 36921 40072
rect 36955 40069 36967 40103
rect 36909 40063 36967 40069
rect 38286 40060 38292 40112
rect 38344 40060 38350 40112
rect 38838 40060 38844 40112
rect 38896 40100 38902 40112
rect 39669 40103 39727 40109
rect 39669 40100 39681 40103
rect 38896 40072 39681 40100
rect 38896 40060 38902 40072
rect 39669 40069 39681 40072
rect 39715 40069 39727 40103
rect 39669 40063 39727 40069
rect 37458 40032 37464 40044
rect 36556 40004 37464 40032
rect 25056 39936 25360 39964
rect 25332 39908 25360 39936
rect 26050 39924 26056 39976
rect 26108 39924 26114 39976
rect 26789 39967 26847 39973
rect 26789 39933 26801 39967
rect 26835 39964 26847 39967
rect 26970 39964 26976 39976
rect 26835 39936 26976 39964
rect 26835 39933 26847 39936
rect 26789 39927 26847 39933
rect 26970 39924 26976 39936
rect 27028 39924 27034 39976
rect 27890 39924 27896 39976
rect 27948 39924 27954 39976
rect 25225 39899 25283 39905
rect 21140 39868 22968 39896
rect 24596 39868 24900 39896
rect 21140 39856 21146 39868
rect 18782 39788 18788 39840
rect 18840 39828 18846 39840
rect 18877 39831 18935 39837
rect 18877 39828 18889 39831
rect 18840 39800 18889 39828
rect 18840 39788 18846 39800
rect 18877 39797 18889 39800
rect 18923 39797 18935 39831
rect 18877 39791 18935 39797
rect 22094 39788 22100 39840
rect 22152 39828 22158 39840
rect 22940 39837 22968 39868
rect 22373 39831 22431 39837
rect 22373 39828 22385 39831
rect 22152 39800 22385 39828
rect 22152 39788 22158 39800
rect 22373 39797 22385 39800
rect 22419 39797 22431 39831
rect 22373 39791 22431 39797
rect 22925 39831 22983 39837
rect 22925 39797 22937 39831
rect 22971 39797 22983 39831
rect 22925 39791 22983 39797
rect 24762 39788 24768 39840
rect 24820 39788 24826 39840
rect 24872 39828 24900 39868
rect 25225 39865 25237 39899
rect 25271 39865 25283 39899
rect 25225 39859 25283 39865
rect 25240 39828 25268 39859
rect 25314 39856 25320 39908
rect 25372 39856 25378 39908
rect 28350 39856 28356 39908
rect 28408 39856 28414 39908
rect 30837 39899 30895 39905
rect 30837 39865 30849 39899
rect 30883 39896 30895 39899
rect 32232 39896 32260 39995
rect 32490 39896 32496 39908
rect 30883 39868 32496 39896
rect 30883 39865 30895 39868
rect 30837 39859 30895 39865
rect 32490 39856 32496 39868
rect 32548 39856 32554 39908
rect 36556 39905 36584 40004
rect 37458 39992 37464 40004
rect 37516 39992 37522 40044
rect 39117 39967 39175 39973
rect 39117 39933 39129 39967
rect 39163 39964 39175 39967
rect 39206 39964 39212 39976
rect 39163 39936 39212 39964
rect 39163 39933 39175 39936
rect 39117 39927 39175 39933
rect 39206 39924 39212 39936
rect 39264 39924 39270 39976
rect 39850 39924 39856 39976
rect 39908 39924 39914 39976
rect 36541 39899 36599 39905
rect 36541 39865 36553 39899
rect 36587 39865 36599 39899
rect 36541 39859 36599 39865
rect 24872 39800 25268 39828
rect 32398 39788 32404 39840
rect 32456 39788 32462 39840
rect 32674 39788 32680 39840
rect 32732 39828 32738 39840
rect 35342 39828 35348 39840
rect 32732 39800 35348 39828
rect 32732 39788 32738 39800
rect 35342 39788 35348 39800
rect 35400 39788 35406 39840
rect 1104 39738 42504 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 42504 39738
rect 1104 39664 42504 39686
rect 30009 39627 30067 39633
rect 30009 39593 30021 39627
rect 30055 39624 30067 39627
rect 30098 39624 30104 39636
rect 30055 39596 30104 39624
rect 30055 39593 30067 39596
rect 30009 39587 30067 39593
rect 30098 39584 30104 39596
rect 30156 39584 30162 39636
rect 30558 39584 30564 39636
rect 30616 39624 30622 39636
rect 30837 39627 30895 39633
rect 30837 39624 30849 39627
rect 30616 39596 30849 39624
rect 30616 39584 30622 39596
rect 30837 39593 30849 39596
rect 30883 39593 30895 39627
rect 30837 39587 30895 39593
rect 32030 39584 32036 39636
rect 32088 39624 32094 39636
rect 32125 39627 32183 39633
rect 32125 39624 32137 39627
rect 32088 39596 32137 39624
rect 32088 39584 32094 39596
rect 32125 39593 32137 39596
rect 32171 39593 32183 39627
rect 32125 39587 32183 39593
rect 32214 39584 32220 39636
rect 32272 39624 32278 39636
rect 32582 39624 32588 39636
rect 32272 39596 32588 39624
rect 32272 39584 32278 39596
rect 32582 39584 32588 39596
rect 32640 39624 32646 39636
rect 32861 39627 32919 39633
rect 32861 39624 32873 39627
rect 32640 39596 32873 39624
rect 32640 39584 32646 39596
rect 32861 39593 32873 39596
rect 32907 39593 32919 39627
rect 32861 39587 32919 39593
rect 33502 39584 33508 39636
rect 33560 39624 33566 39636
rect 34882 39624 34888 39636
rect 33560 39596 34888 39624
rect 33560 39584 33566 39596
rect 34882 39584 34888 39596
rect 34940 39584 34946 39636
rect 35250 39584 35256 39636
rect 35308 39624 35314 39636
rect 35621 39627 35679 39633
rect 35621 39624 35633 39627
rect 35308 39596 35633 39624
rect 35308 39584 35314 39596
rect 35621 39593 35633 39596
rect 35667 39593 35679 39627
rect 35621 39587 35679 39593
rect 24578 39516 24584 39568
rect 24636 39556 24642 39568
rect 31110 39556 31116 39568
rect 24636 39528 31116 39556
rect 24636 39516 24642 39528
rect 31110 39516 31116 39528
rect 31168 39556 31174 39568
rect 34517 39559 34575 39565
rect 31168 39528 34284 39556
rect 31168 39516 31174 39528
rect 18782 39448 18788 39500
rect 18840 39448 18846 39500
rect 22186 39448 22192 39500
rect 22244 39488 22250 39500
rect 22925 39491 22983 39497
rect 22925 39488 22937 39491
rect 22244 39460 22937 39488
rect 22244 39448 22250 39460
rect 22925 39457 22937 39460
rect 22971 39457 22983 39491
rect 24596 39488 24624 39516
rect 22925 39451 22983 39457
rect 23952 39460 24624 39488
rect 24857 39491 24915 39497
rect 18690 39380 18696 39432
rect 18748 39380 18754 39432
rect 22094 39380 22100 39432
rect 22152 39420 22158 39432
rect 22649 39423 22707 39429
rect 22649 39420 22661 39423
rect 22152 39392 22661 39420
rect 22152 39380 22158 39392
rect 22649 39389 22661 39392
rect 22695 39389 22707 39423
rect 22649 39383 22707 39389
rect 22741 39423 22799 39429
rect 22741 39389 22753 39423
rect 22787 39389 22799 39423
rect 22741 39383 22799 39389
rect 22833 39423 22891 39429
rect 22833 39389 22845 39423
rect 22879 39420 22891 39423
rect 23952 39420 23980 39460
rect 24857 39457 24869 39491
rect 24903 39488 24915 39491
rect 25593 39491 25651 39497
rect 25593 39488 25605 39491
rect 24903 39460 25605 39488
rect 24903 39457 24915 39460
rect 24857 39451 24915 39457
rect 25593 39457 25605 39460
rect 25639 39457 25651 39491
rect 25593 39451 25651 39457
rect 30653 39491 30711 39497
rect 30653 39457 30665 39491
rect 30699 39488 30711 39491
rect 30834 39488 30840 39500
rect 30699 39460 30840 39488
rect 30699 39457 30711 39460
rect 30653 39451 30711 39457
rect 30834 39448 30840 39460
rect 30892 39488 30898 39500
rect 31478 39488 31484 39500
rect 30892 39460 31484 39488
rect 30892 39448 30898 39460
rect 31478 39448 31484 39460
rect 31536 39448 31542 39500
rect 32030 39448 32036 39500
rect 32088 39488 32094 39500
rect 32493 39491 32551 39497
rect 32493 39488 32505 39491
rect 32088 39460 32505 39488
rect 32088 39448 32094 39460
rect 32493 39457 32505 39460
rect 32539 39457 32551 39491
rect 32493 39451 32551 39457
rect 32674 39448 32680 39500
rect 32732 39448 32738 39500
rect 34256 39488 34284 39528
rect 34517 39525 34529 39559
rect 34563 39525 34575 39559
rect 34517 39519 34575 39525
rect 34532 39488 34560 39519
rect 34606 39516 34612 39568
rect 34664 39556 34670 39568
rect 34664 39528 35756 39556
rect 34664 39516 34670 39528
rect 35253 39491 35311 39497
rect 34256 39460 34376 39488
rect 34532 39460 35020 39488
rect 22879 39392 23980 39420
rect 24029 39423 24087 39429
rect 22879 39389 22891 39392
rect 22833 39383 22891 39389
rect 24029 39389 24041 39423
rect 24075 39420 24087 39423
rect 24302 39420 24308 39432
rect 24075 39392 24308 39420
rect 24075 39389 24087 39392
rect 24029 39383 24087 39389
rect 21818 39312 21824 39364
rect 21876 39352 21882 39364
rect 22756 39352 22784 39383
rect 24302 39380 24308 39392
rect 24360 39380 24366 39432
rect 24762 39380 24768 39432
rect 24820 39380 24826 39432
rect 25222 39380 25228 39432
rect 25280 39380 25286 39432
rect 25314 39380 25320 39432
rect 25372 39420 25378 39432
rect 31757 39423 31815 39429
rect 25372 39392 25417 39420
rect 25372 39380 25378 39392
rect 31757 39389 31769 39423
rect 31803 39420 31815 39423
rect 31846 39420 31852 39432
rect 31803 39392 31852 39420
rect 31803 39389 31815 39392
rect 31757 39383 31815 39389
rect 31846 39380 31852 39392
rect 31904 39420 31910 39432
rect 32214 39420 32220 39432
rect 31904 39392 32220 39420
rect 31904 39380 31910 39392
rect 32214 39380 32220 39392
rect 32272 39380 32278 39432
rect 32306 39380 32312 39432
rect 32364 39420 32370 39432
rect 32401 39423 32459 39429
rect 32401 39420 32413 39423
rect 32364 39392 32413 39420
rect 32364 39380 32370 39392
rect 32401 39389 32413 39392
rect 32447 39389 32459 39423
rect 32401 39383 32459 39389
rect 21876 39324 22784 39352
rect 30377 39355 30435 39361
rect 21876 39312 21882 39324
rect 30377 39321 30389 39355
rect 30423 39352 30435 39355
rect 30926 39352 30932 39364
rect 30423 39324 30932 39352
rect 30423 39321 30435 39324
rect 30377 39315 30435 39321
rect 30926 39312 30932 39324
rect 30984 39352 30990 39364
rect 31297 39355 31355 39361
rect 31297 39352 31309 39355
rect 30984 39324 31309 39352
rect 30984 39312 30990 39324
rect 31297 39321 31309 39324
rect 31343 39321 31355 39355
rect 31297 39315 31355 39321
rect 31938 39312 31944 39364
rect 31996 39352 32002 39364
rect 32416 39352 32444 39383
rect 32582 39380 32588 39432
rect 32640 39380 32646 39432
rect 32861 39423 32919 39429
rect 32861 39389 32873 39423
rect 32907 39389 32919 39423
rect 32861 39383 32919 39389
rect 32953 39423 33011 39429
rect 32953 39389 32965 39423
rect 32999 39389 33011 39423
rect 32953 39383 33011 39389
rect 32876 39352 32904 39383
rect 31996 39324 32352 39352
rect 32416 39324 32904 39352
rect 31996 39312 32002 39324
rect 19061 39287 19119 39293
rect 19061 39253 19073 39287
rect 19107 39284 19119 39287
rect 19702 39284 19708 39296
rect 19107 39256 19708 39284
rect 19107 39253 19119 39256
rect 19061 39247 19119 39253
rect 19702 39244 19708 39256
rect 19760 39244 19766 39296
rect 22465 39287 22523 39293
rect 22465 39253 22477 39287
rect 22511 39284 22523 39287
rect 22646 39284 22652 39296
rect 22511 39256 22652 39284
rect 22511 39253 22523 39256
rect 22465 39247 22523 39253
rect 22646 39244 22652 39256
rect 22704 39244 22710 39296
rect 25133 39287 25191 39293
rect 25133 39253 25145 39287
rect 25179 39284 25191 39287
rect 25590 39284 25596 39296
rect 25179 39256 25596 39284
rect 25179 39253 25191 39256
rect 25133 39247 25191 39253
rect 25590 39244 25596 39256
rect 25648 39244 25654 39296
rect 30469 39287 30527 39293
rect 30469 39253 30481 39287
rect 30515 39284 30527 39287
rect 30558 39284 30564 39296
rect 30515 39256 30564 39284
rect 30515 39253 30527 39256
rect 30469 39247 30527 39253
rect 30558 39244 30564 39256
rect 30616 39284 30622 39296
rect 31205 39287 31263 39293
rect 31205 39284 31217 39287
rect 30616 39256 31217 39284
rect 30616 39244 30622 39256
rect 31205 39253 31217 39256
rect 31251 39253 31263 39287
rect 31205 39247 31263 39253
rect 32214 39244 32220 39296
rect 32272 39244 32278 39296
rect 32324 39284 32352 39324
rect 32968 39284 32996 39383
rect 34238 39380 34244 39432
rect 34296 39380 34302 39432
rect 34348 39429 34376 39460
rect 34333 39423 34391 39429
rect 34333 39389 34345 39423
rect 34379 39389 34391 39423
rect 34333 39383 34391 39389
rect 34440 39392 34744 39420
rect 34440 39352 34468 39392
rect 34348 39324 34468 39352
rect 34348 39296 34376 39324
rect 34514 39312 34520 39364
rect 34572 39312 34578 39364
rect 34716 39352 34744 39392
rect 34790 39380 34796 39432
rect 34848 39420 34854 39432
rect 34992 39429 35020 39460
rect 35253 39457 35265 39491
rect 35299 39488 35311 39491
rect 35342 39488 35348 39500
rect 35299 39460 35348 39488
rect 35299 39457 35311 39460
rect 35253 39451 35311 39457
rect 35342 39448 35348 39460
rect 35400 39448 35406 39500
rect 34885 39423 34943 39429
rect 34885 39420 34897 39423
rect 34848 39392 34897 39420
rect 34848 39380 34854 39392
rect 34885 39389 34897 39392
rect 34931 39389 34943 39423
rect 34885 39383 34943 39389
rect 34977 39423 35035 39429
rect 34977 39389 34989 39423
rect 35023 39389 35035 39423
rect 35621 39423 35679 39429
rect 35621 39420 35633 39423
rect 34977 39383 35035 39389
rect 35084 39392 35633 39420
rect 35084 39352 35112 39392
rect 35621 39389 35633 39392
rect 35667 39389 35679 39423
rect 35728 39420 35756 39528
rect 38562 39516 38568 39568
rect 38620 39556 38626 39568
rect 39393 39559 39451 39565
rect 39393 39556 39405 39559
rect 38620 39528 39405 39556
rect 38620 39516 38626 39528
rect 39393 39525 39405 39528
rect 39439 39525 39451 39559
rect 39393 39519 39451 39525
rect 40218 39448 40224 39500
rect 40276 39488 40282 39500
rect 40405 39491 40463 39497
rect 40405 39488 40417 39491
rect 40276 39460 40417 39488
rect 40276 39448 40282 39460
rect 40405 39457 40417 39460
rect 40451 39457 40463 39491
rect 40405 39451 40463 39457
rect 35805 39423 35863 39429
rect 35805 39420 35817 39423
rect 35728 39392 35817 39420
rect 35621 39383 35679 39389
rect 35805 39389 35817 39392
rect 35851 39389 35863 39423
rect 35805 39383 35863 39389
rect 34716 39324 35112 39352
rect 35158 39312 35164 39364
rect 35216 39352 35222 39364
rect 35345 39355 35403 39361
rect 35345 39352 35357 39355
rect 35216 39324 35357 39352
rect 35216 39312 35222 39324
rect 35345 39321 35357 39324
rect 35391 39321 35403 39355
rect 35636 39352 35664 39383
rect 36814 39380 36820 39432
rect 36872 39420 36878 39432
rect 37277 39423 37335 39429
rect 37277 39420 37289 39423
rect 36872 39392 37289 39420
rect 36872 39380 36878 39392
rect 37277 39389 37289 39392
rect 37323 39389 37335 39423
rect 37277 39383 37335 39389
rect 36630 39352 36636 39364
rect 35636 39324 36636 39352
rect 35345 39315 35403 39321
rect 36630 39312 36636 39324
rect 36688 39312 36694 39364
rect 37292 39352 37320 39383
rect 37366 39380 37372 39432
rect 37424 39420 37430 39432
rect 37461 39423 37519 39429
rect 37461 39420 37473 39423
rect 37424 39392 37473 39420
rect 37424 39380 37430 39392
rect 37461 39389 37473 39392
rect 37507 39389 37519 39423
rect 37461 39383 37519 39389
rect 39666 39380 39672 39432
rect 39724 39380 39730 39432
rect 40954 39420 40960 39432
rect 40144 39392 40960 39420
rect 38194 39352 38200 39364
rect 37292 39324 38200 39352
rect 38194 39312 38200 39324
rect 38252 39312 38258 39364
rect 39390 39312 39396 39364
rect 39448 39352 39454 39364
rect 40144 39352 40172 39392
rect 40954 39380 40960 39392
rect 41012 39420 41018 39432
rect 41233 39423 41291 39429
rect 41233 39420 41245 39423
rect 41012 39392 41245 39420
rect 41012 39380 41018 39392
rect 41233 39389 41245 39392
rect 41279 39389 41291 39423
rect 41233 39383 41291 39389
rect 42150 39380 42156 39432
rect 42208 39380 42214 39432
rect 39448 39324 40172 39352
rect 40221 39355 40279 39361
rect 39448 39312 39454 39324
rect 40221 39321 40233 39355
rect 40267 39352 40279 39355
rect 40681 39355 40739 39361
rect 40681 39352 40693 39355
rect 40267 39324 40693 39352
rect 40267 39321 40279 39324
rect 40221 39315 40279 39321
rect 40681 39321 40693 39324
rect 40727 39321 40739 39355
rect 40681 39315 40739 39321
rect 32324 39256 32996 39284
rect 33229 39287 33287 39293
rect 33229 39253 33241 39287
rect 33275 39284 33287 39287
rect 34330 39284 34336 39296
rect 33275 39256 34336 39284
rect 33275 39253 33287 39256
rect 33229 39247 33287 39253
rect 34330 39244 34336 39256
rect 34388 39244 34394 39296
rect 34422 39244 34428 39296
rect 34480 39284 34486 39296
rect 34701 39287 34759 39293
rect 34701 39284 34713 39287
rect 34480 39256 34713 39284
rect 34480 39244 34486 39256
rect 34701 39253 34713 39256
rect 34747 39253 34759 39287
rect 34701 39247 34759 39253
rect 35434 39244 35440 39296
rect 35492 39244 35498 39296
rect 37369 39287 37427 39293
rect 37369 39253 37381 39287
rect 37415 39284 37427 39287
rect 37642 39284 37648 39296
rect 37415 39256 37648 39284
rect 37415 39253 37427 39256
rect 37369 39247 37427 39253
rect 37642 39244 37648 39256
rect 37700 39244 37706 39296
rect 39574 39244 39580 39296
rect 39632 39244 39638 39296
rect 39758 39244 39764 39296
rect 39816 39284 39822 39296
rect 39853 39287 39911 39293
rect 39853 39284 39865 39287
rect 39816 39256 39865 39284
rect 39816 39244 39822 39256
rect 39853 39253 39865 39256
rect 39899 39253 39911 39287
rect 39853 39247 39911 39253
rect 40310 39244 40316 39296
rect 40368 39244 40374 39296
rect 41414 39244 41420 39296
rect 41472 39284 41478 39296
rect 41509 39287 41567 39293
rect 41509 39284 41521 39287
rect 41472 39256 41521 39284
rect 41472 39244 41478 39256
rect 41509 39253 41521 39256
rect 41555 39253 41567 39287
rect 41509 39247 41567 39253
rect 1104 39194 42504 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 42504 39194
rect 1104 39120 42504 39142
rect 17129 39083 17187 39089
rect 17129 39049 17141 39083
rect 17175 39080 17187 39083
rect 17218 39080 17224 39092
rect 17175 39052 17224 39080
rect 17175 39049 17187 39052
rect 17129 39043 17187 39049
rect 17218 39040 17224 39052
rect 17276 39040 17282 39092
rect 17497 39083 17555 39089
rect 17497 39049 17509 39083
rect 17543 39080 17555 39083
rect 18690 39080 18696 39092
rect 17543 39052 18696 39080
rect 17543 39049 17555 39052
rect 17497 39043 17555 39049
rect 18690 39040 18696 39052
rect 18748 39040 18754 39092
rect 23474 39080 23480 39092
rect 19628 39052 20484 39080
rect 16574 38972 16580 39024
rect 16632 39012 16638 39024
rect 17037 39015 17095 39021
rect 17037 39012 17049 39015
rect 16632 38984 17049 39012
rect 16632 38972 16638 38984
rect 17037 38981 17049 38984
rect 17083 39012 17095 39015
rect 17083 38984 18552 39012
rect 17083 38981 17095 38984
rect 17037 38975 17095 38981
rect 14734 38904 14740 38956
rect 14792 38904 14798 38956
rect 16114 38904 16120 38956
rect 16172 38904 16178 38956
rect 18524 38953 18552 38984
rect 19628 38953 19656 39052
rect 20254 39021 20260 39024
rect 20225 39015 20260 39021
rect 20225 39012 20237 39015
rect 19812 38984 20237 39012
rect 18509 38947 18567 38953
rect 18509 38913 18521 38947
rect 18555 38913 18567 38947
rect 19613 38947 19671 38953
rect 19613 38944 19625 38947
rect 18509 38907 18567 38913
rect 18892 38916 19625 38944
rect 15013 38879 15071 38885
rect 15013 38845 15025 38879
rect 15059 38876 15071 38879
rect 16482 38876 16488 38888
rect 15059 38848 16488 38876
rect 15059 38845 15071 38848
rect 15013 38839 15071 38845
rect 16482 38836 16488 38848
rect 16540 38836 16546 38888
rect 16853 38879 16911 38885
rect 16853 38845 16865 38879
rect 16899 38845 16911 38879
rect 16853 38839 16911 38845
rect 18141 38879 18199 38885
rect 18141 38845 18153 38879
rect 18187 38876 18199 38879
rect 18417 38879 18475 38885
rect 18417 38876 18429 38879
rect 18187 38848 18429 38876
rect 18187 38845 18199 38848
rect 18141 38839 18199 38845
rect 18417 38845 18429 38848
rect 18463 38845 18475 38879
rect 18417 38839 18475 38845
rect 16868 38808 16896 38839
rect 18156 38808 18184 38839
rect 16500 38780 18184 38808
rect 16500 38749 16528 38780
rect 16485 38743 16543 38749
rect 16485 38709 16497 38743
rect 16531 38709 16543 38743
rect 16485 38703 16543 38709
rect 17586 38700 17592 38752
rect 17644 38700 17650 38752
rect 18414 38700 18420 38752
rect 18472 38740 18478 38752
rect 18892 38749 18920 38916
rect 19613 38913 19625 38916
rect 19659 38913 19671 38947
rect 19613 38907 19671 38913
rect 19702 38904 19708 38956
rect 19760 38944 19766 38956
rect 19812 38944 19840 38984
rect 20225 38981 20237 38984
rect 20225 38975 20260 38981
rect 20254 38972 20260 38975
rect 20312 38972 20318 39024
rect 20346 38972 20352 39024
rect 20404 39012 20410 39024
rect 20456 39021 20484 39052
rect 22204 39052 23480 39080
rect 20441 39015 20499 39021
rect 20441 39012 20453 39015
rect 20404 38984 20453 39012
rect 20404 38972 20410 38984
rect 20441 38981 20453 38984
rect 20487 38981 20499 39015
rect 20441 38975 20499 38981
rect 21082 38972 21088 39024
rect 21140 39012 21146 39024
rect 21269 39015 21327 39021
rect 21269 39012 21281 39015
rect 21140 38984 21281 39012
rect 21140 38972 21146 38984
rect 21269 38981 21281 38984
rect 21315 38981 21327 39015
rect 21269 38975 21327 38981
rect 22094 38972 22100 39024
rect 22152 38972 22158 39024
rect 19760 38916 19840 38944
rect 19760 38904 19766 38916
rect 20806 38904 20812 38956
rect 20864 38904 20870 38956
rect 21450 38944 21456 38956
rect 20916 38916 21456 38944
rect 19981 38879 20039 38885
rect 19981 38845 19993 38879
rect 20027 38876 20039 38879
rect 20916 38876 20944 38916
rect 21450 38904 21456 38916
rect 21508 38904 21514 38956
rect 21637 38947 21695 38953
rect 21637 38913 21649 38947
rect 21683 38944 21695 38947
rect 21818 38944 21824 38956
rect 21683 38916 21824 38944
rect 21683 38913 21695 38916
rect 21637 38907 21695 38913
rect 21818 38904 21824 38916
rect 21876 38904 21882 38956
rect 22204 38953 22232 39052
rect 23474 39040 23480 39052
rect 23532 39080 23538 39092
rect 24302 39080 24308 39092
rect 23532 39052 24308 39080
rect 23532 39040 23538 39052
rect 24302 39040 24308 39052
rect 24360 39040 24366 39092
rect 25041 39083 25099 39089
rect 25041 39049 25053 39083
rect 25087 39080 25099 39083
rect 25314 39080 25320 39092
rect 25087 39052 25320 39080
rect 25087 39049 25099 39052
rect 25041 39043 25099 39049
rect 25314 39040 25320 39052
rect 25372 39040 25378 39092
rect 28534 39080 28540 39092
rect 28092 39052 28540 39080
rect 23934 39012 23940 39024
rect 23690 38984 23940 39012
rect 23934 38972 23940 38984
rect 23992 38972 23998 39024
rect 24872 38984 25176 39012
rect 24872 38956 24900 38984
rect 21913 38947 21971 38953
rect 21913 38913 21925 38947
rect 21959 38913 21971 38947
rect 21913 38907 21971 38913
rect 22189 38947 22247 38953
rect 22189 38913 22201 38947
rect 22235 38913 22247 38947
rect 22189 38907 22247 38913
rect 24765 38947 24823 38953
rect 24765 38913 24777 38947
rect 24811 38944 24823 38947
rect 24854 38944 24860 38956
rect 24811 38916 24860 38944
rect 24811 38913 24823 38916
rect 24765 38907 24823 38913
rect 21928 38876 21956 38907
rect 24854 38904 24860 38916
rect 24912 38904 24918 38956
rect 24949 38947 25007 38953
rect 24949 38913 24961 38947
rect 24995 38913 25007 38947
rect 24949 38907 25007 38913
rect 20027 38848 20944 38876
rect 21836 38848 21956 38876
rect 20027 38845 20039 38848
rect 19981 38839 20039 38845
rect 19334 38768 19340 38820
rect 19392 38808 19398 38820
rect 20622 38808 20628 38820
rect 19392 38780 20628 38808
rect 19392 38768 19398 38780
rect 20622 38768 20628 38780
rect 20680 38768 20686 38820
rect 18877 38743 18935 38749
rect 18877 38740 18889 38743
rect 18472 38712 18889 38740
rect 18472 38700 18478 38712
rect 18877 38709 18889 38712
rect 18923 38709 18935 38743
rect 18877 38703 18935 38709
rect 20070 38700 20076 38752
rect 20128 38700 20134 38752
rect 20257 38743 20315 38749
rect 20257 38709 20269 38743
rect 20303 38740 20315 38743
rect 20530 38740 20536 38752
rect 20303 38712 20536 38740
rect 20303 38709 20315 38712
rect 20257 38703 20315 38709
rect 20530 38700 20536 38712
rect 20588 38740 20594 38752
rect 21836 38740 21864 38848
rect 22462 38836 22468 38888
rect 22520 38836 22526 38888
rect 24581 38879 24639 38885
rect 24581 38845 24593 38879
rect 24627 38845 24639 38879
rect 24964 38876 24992 38907
rect 25038 38904 25044 38956
rect 25096 38904 25102 38956
rect 25148 38953 25176 38984
rect 25590 38972 25596 39024
rect 25648 38972 25654 39024
rect 25133 38947 25191 38953
rect 25133 38913 25145 38947
rect 25179 38913 25191 38947
rect 25133 38907 25191 38913
rect 25225 38947 25283 38953
rect 25225 38913 25237 38947
rect 25271 38944 25283 38947
rect 25314 38944 25320 38956
rect 25271 38916 25320 38944
rect 25271 38913 25283 38916
rect 25225 38907 25283 38913
rect 25240 38876 25268 38907
rect 25314 38904 25320 38916
rect 25372 38904 25378 38956
rect 25406 38904 25412 38956
rect 25464 38904 25470 38956
rect 28092 38953 28120 39052
rect 28534 39040 28540 39052
rect 28592 39080 28598 39092
rect 29089 39083 29147 39089
rect 28592 39052 28948 39080
rect 28592 39040 28598 39052
rect 28629 39015 28687 39021
rect 28629 38981 28641 39015
rect 28675 39012 28687 39015
rect 28718 39012 28724 39024
rect 28675 38984 28724 39012
rect 28675 38981 28687 38984
rect 28629 38975 28687 38981
rect 28718 38972 28724 38984
rect 28776 38972 28782 39024
rect 25777 38947 25835 38953
rect 25777 38913 25789 38947
rect 25823 38913 25835 38947
rect 28077 38947 28135 38953
rect 28077 38944 28089 38947
rect 25777 38907 25835 38913
rect 26712 38916 28089 38944
rect 24964 38848 25268 38876
rect 24581 38839 24639 38845
rect 23937 38811 23995 38817
rect 23937 38777 23949 38811
rect 23983 38808 23995 38811
rect 24118 38808 24124 38820
rect 23983 38780 24124 38808
rect 23983 38777 23995 38780
rect 23937 38771 23995 38777
rect 24118 38768 24124 38780
rect 24176 38808 24182 38820
rect 24596 38808 24624 38839
rect 24176 38780 24624 38808
rect 24176 38768 24182 38780
rect 25222 38768 25228 38820
rect 25280 38808 25286 38820
rect 25409 38811 25467 38817
rect 25409 38808 25421 38811
rect 25280 38780 25421 38808
rect 25280 38768 25286 38780
rect 25409 38777 25421 38780
rect 25455 38777 25467 38811
rect 25409 38771 25467 38777
rect 20588 38712 21864 38740
rect 22097 38743 22155 38749
rect 20588 38700 20594 38712
rect 22097 38709 22109 38743
rect 22143 38740 22155 38743
rect 22554 38740 22560 38752
rect 22143 38712 22560 38740
rect 22143 38709 22155 38712
rect 22097 38703 22155 38709
rect 22554 38700 22560 38712
rect 22612 38700 22618 38752
rect 24026 38700 24032 38752
rect 24084 38700 24090 38752
rect 24394 38700 24400 38752
rect 24452 38740 24458 38752
rect 25792 38740 25820 38907
rect 26712 38752 26740 38916
rect 28077 38913 28089 38916
rect 28123 38913 28135 38947
rect 28077 38907 28135 38913
rect 28350 38904 28356 38956
rect 28408 38904 28414 38956
rect 28920 38953 28948 39052
rect 29089 39049 29101 39083
rect 29135 39080 29147 39083
rect 31938 39080 31944 39092
rect 29135 39052 31944 39080
rect 29135 39049 29147 39052
rect 29089 39043 29147 39049
rect 30116 38953 30144 39052
rect 31938 39040 31944 39052
rect 31996 39040 32002 39092
rect 32122 39040 32128 39092
rect 32180 39080 32186 39092
rect 33962 39080 33968 39092
rect 32180 39052 33968 39080
rect 32180 39040 32186 39052
rect 33962 39040 33968 39052
rect 34020 39040 34026 39092
rect 36170 39080 36176 39092
rect 34624 39052 36176 39080
rect 30193 39015 30251 39021
rect 30193 38981 30205 39015
rect 30239 39012 30251 39015
rect 34624 39012 34652 39052
rect 36170 39040 36176 39052
rect 36228 39080 36234 39092
rect 36228 39052 36492 39080
rect 36228 39040 36234 39052
rect 30239 38984 30788 39012
rect 30239 38981 30251 38984
rect 30193 38975 30251 38981
rect 30760 38953 30788 38984
rect 33796 38984 34652 39012
rect 28537 38947 28595 38953
rect 28537 38913 28549 38947
rect 28583 38944 28595 38947
rect 28905 38947 28963 38953
rect 28583 38916 28856 38944
rect 28583 38913 28595 38916
rect 28537 38907 28595 38913
rect 28368 38876 28396 38904
rect 28828 38888 28856 38916
rect 28905 38913 28917 38947
rect 28951 38913 28963 38947
rect 28905 38907 28963 38913
rect 30101 38947 30159 38953
rect 30101 38913 30113 38947
rect 30147 38913 30159 38947
rect 30101 38907 30159 38913
rect 30285 38947 30343 38953
rect 30285 38913 30297 38947
rect 30331 38913 30343 38947
rect 30285 38907 30343 38913
rect 30745 38947 30803 38953
rect 30745 38913 30757 38947
rect 30791 38913 30803 38947
rect 30745 38907 30803 38913
rect 31297 38947 31355 38953
rect 31297 38913 31309 38947
rect 31343 38944 31355 38947
rect 31386 38944 31392 38956
rect 31343 38916 31392 38944
rect 31343 38913 31355 38916
rect 31297 38907 31355 38913
rect 28721 38879 28779 38885
rect 28721 38876 28733 38879
rect 28368 38848 28733 38876
rect 28721 38845 28733 38848
rect 28767 38845 28779 38879
rect 28721 38839 28779 38845
rect 28810 38836 28816 38888
rect 28868 38876 28874 38888
rect 30300 38876 30328 38907
rect 31386 38904 31392 38916
rect 31444 38944 31450 38956
rect 31444 38916 32076 38944
rect 31444 38904 31450 38916
rect 28868 38848 30328 38876
rect 28868 38836 28874 38848
rect 30300 38808 30328 38848
rect 30837 38879 30895 38885
rect 30837 38845 30849 38879
rect 30883 38876 30895 38879
rect 31846 38876 31852 38888
rect 30883 38848 31852 38876
rect 30883 38845 30895 38848
rect 30837 38839 30895 38845
rect 31846 38836 31852 38848
rect 31904 38836 31910 38888
rect 28368 38780 28672 38808
rect 30300 38780 31754 38808
rect 24452 38712 25820 38740
rect 25961 38743 26019 38749
rect 24452 38700 24458 38712
rect 25961 38709 25973 38743
rect 26007 38740 26019 38743
rect 26694 38740 26700 38752
rect 26007 38712 26700 38740
rect 26007 38709 26019 38712
rect 25961 38703 26019 38709
rect 26694 38700 26700 38712
rect 26752 38700 26758 38752
rect 26970 38700 26976 38752
rect 27028 38740 27034 38752
rect 28215 38743 28273 38749
rect 28215 38740 28227 38743
rect 27028 38712 28227 38740
rect 27028 38700 27034 38712
rect 28215 38709 28227 38712
rect 28261 38740 28273 38743
rect 28368 38740 28396 38780
rect 28261 38712 28396 38740
rect 28261 38709 28273 38712
rect 28215 38703 28273 38709
rect 28442 38700 28448 38752
rect 28500 38700 28506 38752
rect 28644 38749 28672 38780
rect 28629 38743 28687 38749
rect 28629 38709 28641 38743
rect 28675 38740 28687 38743
rect 28718 38740 28724 38752
rect 28675 38712 28724 38740
rect 28675 38709 28687 38712
rect 28629 38703 28687 38709
rect 28718 38700 28724 38712
rect 28776 38700 28782 38752
rect 30374 38700 30380 38752
rect 30432 38740 30438 38752
rect 30469 38743 30527 38749
rect 30469 38740 30481 38743
rect 30432 38712 30481 38740
rect 30432 38700 30438 38712
rect 30469 38709 30481 38712
rect 30515 38709 30527 38743
rect 30469 38703 30527 38709
rect 31110 38700 31116 38752
rect 31168 38700 31174 38752
rect 31726 38740 31754 38780
rect 31938 38740 31944 38752
rect 31726 38712 31944 38740
rect 31938 38700 31944 38712
rect 31996 38700 32002 38752
rect 32048 38740 32076 38916
rect 32122 38904 32128 38956
rect 32180 38904 32186 38956
rect 33502 38904 33508 38956
rect 33560 38904 33566 38956
rect 32401 38879 32459 38885
rect 32401 38876 32413 38879
rect 32140 38848 32413 38876
rect 32140 38820 32168 38848
rect 32401 38845 32413 38848
rect 32447 38845 32459 38879
rect 32401 38839 32459 38845
rect 32122 38768 32128 38820
rect 32180 38768 32186 38820
rect 33796 38740 33824 38984
rect 34882 38972 34888 39024
rect 34940 38972 34946 39024
rect 33962 38904 33968 38956
rect 34020 38904 34026 38956
rect 36464 38953 36492 39052
rect 40218 39040 40224 39092
rect 40276 39080 40282 39092
rect 40276 39052 40816 39080
rect 40276 39040 40282 39052
rect 38562 39012 38568 39024
rect 38120 38984 38568 39012
rect 38120 38956 38148 38984
rect 38562 38972 38568 38984
rect 38620 39012 38626 39024
rect 39485 39015 39543 39021
rect 38620 38984 38976 39012
rect 38620 38972 38626 38984
rect 36173 38947 36231 38953
rect 36173 38913 36185 38947
rect 36219 38913 36231 38947
rect 36173 38907 36231 38913
rect 36449 38947 36507 38953
rect 36449 38913 36461 38947
rect 36495 38913 36507 38947
rect 36449 38907 36507 38913
rect 34606 38836 34612 38888
rect 34664 38876 34670 38888
rect 35250 38876 35256 38888
rect 34664 38848 35256 38876
rect 34664 38836 34670 38848
rect 35250 38836 35256 38848
rect 35308 38876 35314 38888
rect 36081 38879 36139 38885
rect 36081 38876 36093 38879
rect 35308 38848 36093 38876
rect 35308 38836 35314 38848
rect 36081 38845 36093 38848
rect 36127 38845 36139 38879
rect 36188 38876 36216 38907
rect 36630 38904 36636 38956
rect 36688 38904 36694 38956
rect 37642 38904 37648 38956
rect 37700 38904 37706 38956
rect 38102 38904 38108 38956
rect 38160 38904 38166 38956
rect 38194 38904 38200 38956
rect 38252 38904 38258 38956
rect 38378 38904 38384 38956
rect 38436 38944 38442 38956
rect 38948 38953 38976 38984
rect 39485 38981 39497 39015
rect 39531 39012 39543 39015
rect 39758 39012 39764 39024
rect 39531 38984 39764 39012
rect 39531 38981 39543 38984
rect 39485 38975 39543 38981
rect 39758 38972 39764 38984
rect 39816 38972 39822 39024
rect 40126 38972 40132 39024
rect 40184 38972 40190 39024
rect 40788 39012 40816 39052
rect 40954 39040 40960 39092
rect 41012 39040 41018 39092
rect 41414 39040 41420 39092
rect 41472 39040 41478 39092
rect 41230 39012 41236 39024
rect 40788 38984 41236 39012
rect 41230 38972 41236 38984
rect 41288 39012 41294 39024
rect 41288 38984 41644 39012
rect 41288 38972 41294 38984
rect 38779 38947 38837 38953
rect 38779 38944 38791 38947
rect 38436 38916 38791 38944
rect 38436 38904 38442 38916
rect 38779 38913 38791 38916
rect 38825 38913 38837 38947
rect 38779 38907 38837 38913
rect 38933 38947 38991 38953
rect 38933 38913 38945 38947
rect 38979 38913 38991 38947
rect 38933 38907 38991 38913
rect 36541 38879 36599 38885
rect 36541 38876 36553 38879
rect 36188 38848 36553 38876
rect 36081 38839 36139 38845
rect 36541 38845 36553 38848
rect 36587 38845 36599 38879
rect 36541 38839 36599 38845
rect 37737 38879 37795 38885
rect 37737 38845 37749 38879
rect 37783 38876 37795 38879
rect 38565 38879 38623 38885
rect 38565 38876 38577 38879
rect 37783 38848 38577 38876
rect 37783 38845 37795 38848
rect 37737 38839 37795 38845
rect 38565 38845 38577 38848
rect 38611 38845 38623 38879
rect 38565 38839 38623 38845
rect 35710 38768 35716 38820
rect 35768 38768 35774 38820
rect 36096 38808 36124 38839
rect 39206 38836 39212 38888
rect 39264 38836 39270 38888
rect 41322 38836 41328 38888
rect 41380 38876 41386 38888
rect 41616 38885 41644 38984
rect 41509 38879 41567 38885
rect 41509 38876 41521 38879
rect 41380 38848 41521 38876
rect 41380 38836 41386 38848
rect 41509 38845 41521 38848
rect 41555 38845 41567 38879
rect 41509 38839 41567 38845
rect 41601 38879 41659 38885
rect 41601 38845 41613 38879
rect 41647 38845 41659 38879
rect 41601 38839 41659 38845
rect 37277 38811 37335 38817
rect 37277 38808 37289 38811
rect 36096 38780 37289 38808
rect 37277 38777 37289 38780
rect 37323 38777 37335 38811
rect 37277 38771 37335 38777
rect 37366 38768 37372 38820
rect 37424 38808 37430 38820
rect 38010 38808 38016 38820
rect 37424 38780 38016 38808
rect 37424 38768 37430 38780
rect 38010 38768 38016 38780
rect 38068 38808 38074 38820
rect 38289 38811 38347 38817
rect 38289 38808 38301 38811
rect 38068 38780 38301 38808
rect 38068 38768 38074 38780
rect 38289 38777 38301 38780
rect 38335 38777 38347 38811
rect 38289 38771 38347 38777
rect 32048 38712 33824 38740
rect 33870 38700 33876 38752
rect 33928 38700 33934 38752
rect 34228 38743 34286 38749
rect 34228 38709 34240 38743
rect 34274 38740 34286 38743
rect 34422 38740 34428 38752
rect 34274 38712 34428 38740
rect 34274 38709 34286 38712
rect 34228 38703 34286 38709
rect 34422 38700 34428 38712
rect 34480 38700 34486 38752
rect 34882 38700 34888 38752
rect 34940 38740 34946 38752
rect 35618 38740 35624 38752
rect 34940 38712 35624 38740
rect 34940 38700 34946 38712
rect 35618 38700 35624 38712
rect 35676 38700 35682 38752
rect 35897 38743 35955 38749
rect 35897 38709 35909 38743
rect 35943 38740 35955 38743
rect 35986 38740 35992 38752
rect 35943 38712 35992 38740
rect 35943 38709 35955 38712
rect 35897 38703 35955 38709
rect 35986 38700 35992 38712
rect 36044 38700 36050 38752
rect 37826 38700 37832 38752
rect 37884 38740 37890 38752
rect 37921 38743 37979 38749
rect 37921 38740 37933 38743
rect 37884 38712 37933 38740
rect 37884 38700 37890 38712
rect 37921 38709 37933 38712
rect 37967 38709 37979 38743
rect 37921 38703 37979 38709
rect 41046 38700 41052 38752
rect 41104 38700 41110 38752
rect 1104 38650 42504 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 42504 38650
rect 1104 38576 42504 38598
rect 16482 38496 16488 38548
rect 16540 38536 16546 38548
rect 16669 38539 16727 38545
rect 16669 38536 16681 38539
rect 16540 38508 16681 38536
rect 16540 38496 16546 38508
rect 16669 38505 16681 38508
rect 16715 38505 16727 38539
rect 16669 38499 16727 38505
rect 17402 38496 17408 38548
rect 17460 38536 17466 38548
rect 20990 38536 20996 38548
rect 17460 38508 20996 38536
rect 17460 38496 17466 38508
rect 20990 38496 20996 38508
rect 21048 38496 21054 38548
rect 21450 38496 21456 38548
rect 21508 38536 21514 38548
rect 21508 38508 22140 38536
rect 21508 38496 21514 38508
rect 16574 38428 16580 38480
rect 16632 38428 16638 38480
rect 19705 38471 19763 38477
rect 19705 38437 19717 38471
rect 19751 38468 19763 38471
rect 20257 38471 20315 38477
rect 20257 38468 20269 38471
rect 19751 38440 20269 38468
rect 19751 38437 19763 38440
rect 19705 38431 19763 38437
rect 20257 38437 20269 38440
rect 20303 38437 20315 38471
rect 20257 38431 20315 38437
rect 21266 38428 21272 38480
rect 21324 38468 21330 38480
rect 22005 38471 22063 38477
rect 22005 38468 22017 38471
rect 21324 38440 22017 38468
rect 21324 38428 21330 38440
rect 22005 38437 22017 38440
rect 22051 38437 22063 38471
rect 22112 38468 22140 38508
rect 22462 38496 22468 38548
rect 22520 38496 22526 38548
rect 24854 38496 24860 38548
rect 24912 38496 24918 38548
rect 25314 38496 25320 38548
rect 25372 38536 25378 38548
rect 26053 38539 26111 38545
rect 26053 38536 26065 38539
rect 25372 38508 26065 38536
rect 25372 38496 25378 38508
rect 26053 38505 26065 38508
rect 26099 38505 26111 38539
rect 31846 38536 31852 38548
rect 26053 38499 26111 38505
rect 26151 38508 31852 38536
rect 23014 38468 23020 38480
rect 22112 38440 23020 38468
rect 22005 38431 22063 38437
rect 17310 38360 17316 38412
rect 17368 38360 17374 38412
rect 19613 38403 19671 38409
rect 19613 38369 19625 38403
rect 19659 38400 19671 38403
rect 20070 38400 20076 38412
rect 19659 38372 20076 38400
rect 19659 38369 19671 38372
rect 19613 38363 19671 38369
rect 20070 38360 20076 38372
rect 20128 38360 20134 38412
rect 20993 38403 21051 38409
rect 20993 38400 21005 38403
rect 20364 38372 21005 38400
rect 14826 38292 14832 38344
rect 14884 38292 14890 38344
rect 17494 38292 17500 38344
rect 17552 38292 17558 38344
rect 19334 38292 19340 38344
rect 19392 38332 19398 38344
rect 19521 38335 19579 38341
rect 19521 38332 19533 38335
rect 19392 38304 19533 38332
rect 19392 38292 19398 38304
rect 19521 38301 19533 38304
rect 19567 38301 19579 38335
rect 19521 38295 19579 38301
rect 19797 38335 19855 38341
rect 19797 38301 19809 38335
rect 19843 38332 19855 38335
rect 20364 38332 20392 38372
rect 20993 38369 21005 38372
rect 21039 38369 21051 38403
rect 20993 38363 21051 38369
rect 21082 38360 21088 38412
rect 21140 38400 21146 38412
rect 21545 38403 21603 38409
rect 21545 38400 21557 38403
rect 21140 38372 21557 38400
rect 21140 38360 21146 38372
rect 21545 38369 21557 38372
rect 21591 38400 21603 38403
rect 21591 38372 22048 38400
rect 21591 38369 21603 38372
rect 21545 38363 21603 38369
rect 19843 38304 20392 38332
rect 19843 38301 19855 38304
rect 19797 38295 19855 38301
rect 20530 38292 20536 38344
rect 20588 38332 20594 38344
rect 20588 38304 21404 38332
rect 20588 38292 20594 38304
rect 15102 38224 15108 38276
rect 15160 38224 15166 38276
rect 16114 38224 16120 38276
rect 16172 38224 16178 38276
rect 17037 38267 17095 38273
rect 17037 38233 17049 38267
rect 17083 38264 17095 38267
rect 17586 38264 17592 38276
rect 17083 38236 17592 38264
rect 17083 38233 17095 38236
rect 17037 38227 17095 38233
rect 17586 38224 17592 38236
rect 17644 38224 17650 38276
rect 18138 38224 18144 38276
rect 18196 38264 18202 38276
rect 18417 38267 18475 38273
rect 18417 38264 18429 38267
rect 18196 38236 18429 38264
rect 18196 38224 18202 38236
rect 18417 38233 18429 38236
rect 18463 38233 18475 38267
rect 18417 38227 18475 38233
rect 18782 38224 18788 38276
rect 18840 38224 18846 38276
rect 20254 38224 20260 38276
rect 20312 38224 20318 38276
rect 20346 38224 20352 38276
rect 20404 38264 20410 38276
rect 20441 38267 20499 38273
rect 20441 38264 20453 38267
rect 20404 38236 20453 38264
rect 20404 38224 20410 38236
rect 20441 38233 20453 38236
rect 20487 38233 20499 38267
rect 20441 38227 20499 38233
rect 17126 38156 17132 38208
rect 17184 38156 17190 38208
rect 17678 38156 17684 38208
rect 17736 38156 17742 38208
rect 19058 38156 19064 38208
rect 19116 38196 19122 38208
rect 19337 38199 19395 38205
rect 19337 38196 19349 38199
rect 19116 38168 19349 38196
rect 19116 38156 19122 38168
rect 19337 38165 19349 38168
rect 19383 38165 19395 38199
rect 19337 38159 19395 38165
rect 19702 38156 19708 38208
rect 19760 38196 19766 38208
rect 20548 38196 20576 38292
rect 20625 38267 20683 38273
rect 20625 38233 20637 38267
rect 20671 38233 20683 38267
rect 20625 38227 20683 38233
rect 19760 38168 20576 38196
rect 20640 38196 20668 38227
rect 20714 38224 20720 38276
rect 20772 38264 20778 38276
rect 20809 38267 20867 38273
rect 20809 38264 20821 38267
rect 20772 38236 20821 38264
rect 20772 38224 20778 38236
rect 20809 38233 20821 38236
rect 20855 38233 20867 38267
rect 21376 38264 21404 38304
rect 21450 38292 21456 38344
rect 21508 38332 21514 38344
rect 21637 38335 21695 38341
rect 21637 38332 21649 38335
rect 21508 38304 21649 38332
rect 21508 38292 21514 38304
rect 21637 38301 21649 38304
rect 21683 38301 21695 38335
rect 21637 38295 21695 38301
rect 21729 38335 21787 38341
rect 21729 38301 21741 38335
rect 21775 38301 21787 38335
rect 21729 38295 21787 38301
rect 21821 38335 21879 38341
rect 21821 38301 21833 38335
rect 21867 38332 21879 38335
rect 21910 38332 21916 38344
rect 21867 38304 21916 38332
rect 21867 38301 21879 38304
rect 21821 38295 21879 38301
rect 21744 38264 21772 38295
rect 21910 38292 21916 38304
rect 21968 38292 21974 38344
rect 22020 38341 22048 38372
rect 22296 38341 22324 38440
rect 23014 38428 23020 38440
rect 23072 38428 23078 38480
rect 26151 38468 26179 38508
rect 31846 38496 31852 38508
rect 31904 38496 31910 38548
rect 32122 38496 32128 38548
rect 32180 38496 32186 38548
rect 34149 38539 34207 38545
rect 34149 38505 34161 38539
rect 34195 38536 34207 38539
rect 34238 38536 34244 38548
rect 34195 38508 34244 38536
rect 34195 38505 34207 38508
rect 34149 38499 34207 38505
rect 34238 38496 34244 38508
rect 34296 38496 34302 38548
rect 34790 38496 34796 38548
rect 34848 38536 34854 38548
rect 35253 38539 35311 38545
rect 35253 38536 35265 38539
rect 34848 38508 35265 38536
rect 34848 38496 34854 38508
rect 35253 38505 35265 38508
rect 35299 38505 35311 38539
rect 35253 38499 35311 38505
rect 39574 38496 39580 38548
rect 39632 38536 39638 38548
rect 39853 38539 39911 38545
rect 39853 38536 39865 38539
rect 39632 38508 39865 38536
rect 39632 38496 39638 38508
rect 39853 38505 39865 38508
rect 39899 38505 39911 38539
rect 39853 38499 39911 38505
rect 40126 38496 40132 38548
rect 40184 38536 40190 38548
rect 41138 38536 41144 38548
rect 40184 38508 41144 38536
rect 40184 38496 40190 38508
rect 41138 38496 41144 38508
rect 41196 38536 41202 38548
rect 41414 38536 41420 38548
rect 41196 38508 41420 38536
rect 41196 38496 41202 38508
rect 41414 38496 41420 38508
rect 41472 38496 41478 38548
rect 42150 38496 42156 38548
rect 42208 38496 42214 38548
rect 24780 38440 26179 38468
rect 26973 38471 27031 38477
rect 22646 38360 22652 38412
rect 22704 38360 22710 38412
rect 23109 38403 23167 38409
rect 23109 38369 23121 38403
rect 23155 38400 23167 38403
rect 24026 38400 24032 38412
rect 23155 38372 24032 38400
rect 23155 38369 23167 38372
rect 23109 38363 23167 38369
rect 24026 38360 24032 38372
rect 24084 38360 24090 38412
rect 24780 38400 24808 38440
rect 24320 38372 24808 38400
rect 22005 38335 22063 38341
rect 22005 38301 22017 38335
rect 22051 38301 22063 38335
rect 22005 38295 22063 38301
rect 22281 38335 22339 38341
rect 22281 38301 22293 38335
rect 22327 38301 22339 38335
rect 22281 38295 22339 38301
rect 22554 38292 22560 38344
rect 22612 38332 22618 38344
rect 22741 38335 22799 38341
rect 22741 38332 22753 38335
rect 22612 38304 22753 38332
rect 22612 38292 22618 38304
rect 22741 38301 22753 38304
rect 22787 38301 22799 38335
rect 22741 38295 22799 38301
rect 22830 38292 22836 38344
rect 22888 38332 22894 38344
rect 24320 38332 24348 38372
rect 22888 38304 24348 38332
rect 22888 38292 22894 38304
rect 24394 38292 24400 38344
rect 24452 38292 24458 38344
rect 24578 38292 24584 38344
rect 24636 38292 24642 38344
rect 24780 38341 24808 38372
rect 25317 38403 25375 38409
rect 25317 38369 25329 38403
rect 25363 38400 25375 38403
rect 25590 38400 25596 38412
rect 25363 38372 25596 38400
rect 25363 38369 25375 38372
rect 25317 38363 25375 38369
rect 25590 38360 25596 38372
rect 25648 38360 25654 38412
rect 24765 38335 24823 38341
rect 24765 38301 24777 38335
rect 24811 38301 24823 38335
rect 24765 38295 24823 38301
rect 24949 38335 25007 38341
rect 24949 38301 24961 38335
rect 24995 38332 25007 38335
rect 25038 38332 25044 38344
rect 24995 38304 25044 38332
rect 24995 38301 25007 38304
rect 24949 38295 25007 38301
rect 25038 38292 25044 38304
rect 25096 38292 25102 38344
rect 25884 38341 25912 38440
rect 26973 38437 26985 38471
rect 27019 38468 27031 38471
rect 27246 38468 27252 38480
rect 27019 38440 27252 38468
rect 27019 38437 27031 38440
rect 26973 38431 27031 38437
rect 27246 38428 27252 38440
rect 27304 38428 27310 38480
rect 27540 38440 31754 38468
rect 27540 38412 27568 38440
rect 27341 38403 27399 38409
rect 27341 38400 27353 38403
rect 26712 38372 27353 38400
rect 26712 38344 26740 38372
rect 27341 38369 27353 38372
rect 27387 38369 27399 38403
rect 27341 38363 27399 38369
rect 27522 38360 27528 38412
rect 27580 38360 27586 38412
rect 28169 38403 28227 38409
rect 28169 38369 28181 38403
rect 28215 38400 28227 38403
rect 28350 38400 28356 38412
rect 28215 38372 28356 38400
rect 28215 38369 28227 38372
rect 28169 38363 28227 38369
rect 28350 38360 28356 38372
rect 28408 38360 28414 38412
rect 28626 38360 28632 38412
rect 28684 38360 28690 38412
rect 25225 38335 25283 38341
rect 25225 38301 25237 38335
rect 25271 38301 25283 38335
rect 25225 38295 25283 38301
rect 25869 38335 25927 38341
rect 25869 38301 25881 38335
rect 25915 38301 25927 38335
rect 25869 38295 25927 38301
rect 22189 38267 22247 38273
rect 22189 38264 22201 38267
rect 21376 38236 22201 38264
rect 20809 38227 20867 38233
rect 22189 38233 22201 38236
rect 22235 38233 22247 38267
rect 22189 38227 22247 38233
rect 20990 38196 20996 38208
rect 20640 38168 20996 38196
rect 19760 38156 19766 38168
rect 20990 38156 20996 38168
rect 21048 38156 21054 38208
rect 21174 38156 21180 38208
rect 21232 38196 21238 38208
rect 21361 38199 21419 38205
rect 21361 38196 21373 38199
rect 21232 38168 21373 38196
rect 21232 38156 21238 38168
rect 21361 38165 21373 38168
rect 21407 38165 21419 38199
rect 22204 38196 22232 38227
rect 23014 38224 23020 38276
rect 23072 38224 23078 38276
rect 24489 38267 24547 38273
rect 24489 38233 24501 38267
rect 24535 38264 24547 38267
rect 25240 38264 25268 38295
rect 26694 38292 26700 38344
rect 26752 38292 26758 38344
rect 26970 38292 26976 38344
rect 27028 38332 27034 38344
rect 27249 38335 27307 38341
rect 27249 38332 27261 38335
rect 27028 38304 27261 38332
rect 27028 38292 27034 38304
rect 27249 38301 27261 38304
rect 27295 38301 27307 38335
rect 27249 38295 27307 38301
rect 27433 38335 27491 38341
rect 27433 38301 27445 38335
rect 27479 38301 27491 38335
rect 27433 38295 27491 38301
rect 28077 38335 28135 38341
rect 28077 38301 28089 38335
rect 28123 38332 28135 38335
rect 28258 38332 28264 38344
rect 28123 38304 28264 38332
rect 28123 38301 28135 38304
rect 28077 38295 28135 38301
rect 24535 38236 25268 38264
rect 24535 38233 24547 38236
rect 24489 38227 24547 38233
rect 25682 38224 25688 38276
rect 25740 38224 25746 38276
rect 26789 38267 26847 38273
rect 26789 38233 26801 38267
rect 26835 38264 26847 38267
rect 27448 38264 27476 38295
rect 28258 38292 28264 38304
rect 28316 38292 28322 38344
rect 28442 38292 28448 38344
rect 28500 38332 28506 38344
rect 28721 38335 28779 38341
rect 28721 38332 28733 38335
rect 28500 38304 28733 38332
rect 28500 38292 28506 38304
rect 28721 38301 28733 38304
rect 28767 38301 28779 38335
rect 28721 38295 28779 38301
rect 28810 38264 28816 38276
rect 26835 38236 28816 38264
rect 26835 38233 26847 38236
rect 26789 38227 26847 38233
rect 28810 38224 28816 38236
rect 28868 38224 28874 38276
rect 31726 38264 31754 38440
rect 34514 38428 34520 38480
rect 34572 38468 34578 38480
rect 35066 38468 35072 38480
rect 34572 38440 35072 38468
rect 34572 38428 34578 38440
rect 35066 38428 35072 38440
rect 35124 38428 35130 38480
rect 38194 38428 38200 38480
rect 38252 38428 38258 38480
rect 38378 38428 38384 38480
rect 38436 38468 38442 38480
rect 39393 38471 39451 38477
rect 39393 38468 39405 38471
rect 38436 38440 39405 38468
rect 38436 38428 38442 38440
rect 39393 38437 39405 38440
rect 39439 38437 39451 38471
rect 39393 38431 39451 38437
rect 32214 38360 32220 38412
rect 32272 38400 32278 38412
rect 32309 38403 32367 38409
rect 32309 38400 32321 38403
rect 32272 38372 32321 38400
rect 32272 38360 32278 38372
rect 32309 38369 32321 38372
rect 32355 38369 32367 38403
rect 32309 38363 32367 38369
rect 32674 38360 32680 38412
rect 32732 38360 32738 38412
rect 33962 38360 33968 38412
rect 34020 38400 34026 38412
rect 35345 38403 35403 38409
rect 35345 38400 35357 38403
rect 34020 38372 35357 38400
rect 34020 38360 34026 38372
rect 35345 38369 35357 38372
rect 35391 38369 35403 38403
rect 35345 38363 35403 38369
rect 37093 38403 37151 38409
rect 37093 38369 37105 38403
rect 37139 38369 37151 38403
rect 37093 38363 37151 38369
rect 32398 38292 32404 38344
rect 32456 38292 32462 38344
rect 32692 38264 32720 38360
rect 32769 38335 32827 38341
rect 32769 38301 32781 38335
rect 32815 38332 32827 38335
rect 33870 38332 33876 38344
rect 32815 38304 33876 38332
rect 32815 38301 32827 38304
rect 32769 38295 32827 38301
rect 33870 38292 33876 38304
rect 33928 38292 33934 38344
rect 34238 38292 34244 38344
rect 34296 38332 34302 38344
rect 34296 38304 34744 38332
rect 34296 38292 34302 38304
rect 31726 38236 32720 38264
rect 34330 38224 34336 38276
rect 34388 38224 34394 38276
rect 34517 38267 34575 38273
rect 34517 38233 34529 38267
rect 34563 38264 34575 38267
rect 34606 38264 34612 38276
rect 34563 38236 34612 38264
rect 34563 38233 34575 38236
rect 34517 38227 34575 38233
rect 34606 38224 34612 38236
rect 34664 38224 34670 38276
rect 34716 38264 34744 38304
rect 34790 38292 34796 38344
rect 34848 38292 34854 38344
rect 34882 38292 34888 38344
rect 34940 38292 34946 38344
rect 34977 38335 35035 38341
rect 34977 38301 34989 38335
rect 35023 38301 35035 38335
rect 34977 38295 35035 38301
rect 34992 38264 35020 38295
rect 35066 38292 35072 38344
rect 35124 38292 35130 38344
rect 37108 38332 37136 38363
rect 38010 38360 38016 38412
rect 38068 38400 38074 38412
rect 38289 38403 38347 38409
rect 38289 38400 38301 38403
rect 38068 38372 38301 38400
rect 38068 38360 38074 38372
rect 38289 38369 38301 38372
rect 38335 38369 38347 38403
rect 38289 38363 38347 38369
rect 37734 38332 37740 38344
rect 37108 38304 37740 38332
rect 37734 38292 37740 38304
rect 37792 38292 37798 38344
rect 38102 38292 38108 38344
rect 38160 38292 38166 38344
rect 38396 38341 38424 38428
rect 39206 38360 39212 38412
rect 39264 38400 39270 38412
rect 40405 38403 40463 38409
rect 40405 38400 40417 38403
rect 39264 38372 40417 38400
rect 39264 38360 39270 38372
rect 40405 38369 40417 38372
rect 40451 38369 40463 38403
rect 40405 38363 40463 38369
rect 40681 38403 40739 38409
rect 40681 38369 40693 38403
rect 40727 38400 40739 38403
rect 41046 38400 41052 38412
rect 40727 38372 41052 38400
rect 40727 38369 40739 38372
rect 40681 38363 40739 38369
rect 41046 38360 41052 38372
rect 41104 38360 41110 38412
rect 38381 38335 38439 38341
rect 38381 38301 38393 38335
rect 38427 38301 38439 38335
rect 38381 38295 38439 38301
rect 38565 38335 38623 38341
rect 38565 38301 38577 38335
rect 38611 38332 38623 38335
rect 38654 38332 38660 38344
rect 38611 38304 38660 38332
rect 38611 38301 38623 38304
rect 38565 38295 38623 38301
rect 38654 38292 38660 38304
rect 38712 38292 38718 38344
rect 39390 38292 39396 38344
rect 39448 38292 39454 38344
rect 39485 38335 39543 38341
rect 39485 38301 39497 38335
rect 39531 38332 39543 38335
rect 39574 38332 39580 38344
rect 39531 38304 39580 38332
rect 39531 38301 39543 38304
rect 39485 38295 39543 38301
rect 39574 38292 39580 38304
rect 39632 38292 39638 38344
rect 39666 38292 39672 38344
rect 39724 38292 39730 38344
rect 40034 38292 40040 38344
rect 40092 38292 40098 38344
rect 34716 38236 35020 38264
rect 35621 38267 35679 38273
rect 35621 38233 35633 38267
rect 35667 38233 35679 38267
rect 35621 38227 35679 38233
rect 24578 38196 24584 38208
rect 22204 38168 24584 38196
rect 21361 38159 21419 38165
rect 24578 38156 24584 38168
rect 24636 38156 24642 38208
rect 25590 38156 25596 38208
rect 25648 38156 25654 38208
rect 27065 38199 27123 38205
rect 27065 38165 27077 38199
rect 27111 38196 27123 38199
rect 27154 38196 27160 38208
rect 27111 38168 27160 38196
rect 27111 38165 27123 38168
rect 27065 38159 27123 38165
rect 27154 38156 27160 38168
rect 27212 38156 27218 38208
rect 28442 38156 28448 38208
rect 28500 38156 28506 38208
rect 29089 38199 29147 38205
rect 29089 38165 29101 38199
rect 29135 38196 29147 38199
rect 29546 38196 29552 38208
rect 29135 38168 29552 38196
rect 29135 38165 29147 38168
rect 29089 38159 29147 38165
rect 29546 38156 29552 38168
rect 29604 38156 29610 38208
rect 31938 38156 31944 38208
rect 31996 38196 32002 38208
rect 32582 38196 32588 38208
rect 31996 38168 32588 38196
rect 31996 38156 32002 38168
rect 32582 38156 32588 38168
rect 32640 38196 32646 38208
rect 34882 38196 34888 38208
rect 32640 38168 34888 38196
rect 32640 38156 32646 38168
rect 34882 38156 34888 38168
rect 34940 38156 34946 38208
rect 35434 38156 35440 38208
rect 35492 38196 35498 38208
rect 35636 38196 35664 38227
rect 35710 38224 35716 38276
rect 35768 38264 35774 38276
rect 40221 38267 40279 38273
rect 35768 38236 36110 38264
rect 35768 38224 35774 38236
rect 40221 38233 40233 38267
rect 40267 38233 40279 38267
rect 40221 38227 40279 38233
rect 35492 38168 35664 38196
rect 35492 38156 35498 38168
rect 37182 38156 37188 38208
rect 37240 38156 37246 38208
rect 37918 38156 37924 38208
rect 37976 38156 37982 38208
rect 40126 38156 40132 38208
rect 40184 38196 40190 38208
rect 40236 38196 40264 38227
rect 41138 38224 41144 38276
rect 41196 38224 41202 38276
rect 42150 38196 42156 38208
rect 40184 38168 42156 38196
rect 40184 38156 40190 38168
rect 42150 38156 42156 38168
rect 42208 38156 42214 38208
rect 1104 38106 42504 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 42504 38106
rect 1104 38032 42504 38054
rect 15102 37952 15108 38004
rect 15160 37992 15166 38004
rect 15657 37995 15715 38001
rect 15657 37992 15669 37995
rect 15160 37964 15669 37992
rect 15160 37952 15166 37964
rect 15657 37961 15669 37964
rect 15703 37961 15715 37995
rect 15657 37955 15715 37961
rect 16025 37995 16083 38001
rect 16025 37961 16037 37995
rect 16071 37992 16083 37995
rect 16669 37995 16727 38001
rect 16669 37992 16681 37995
rect 16071 37964 16681 37992
rect 16071 37961 16083 37964
rect 16025 37955 16083 37961
rect 16669 37961 16681 37964
rect 16715 37961 16727 37995
rect 16669 37955 16727 37961
rect 17678 37952 17684 38004
rect 17736 37992 17742 38004
rect 17736 37964 22094 37992
rect 17736 37952 17742 37964
rect 16850 37924 16856 37936
rect 16316 37896 16856 37924
rect 15746 37856 15752 37868
rect 14766 37828 15752 37856
rect 15746 37816 15752 37828
rect 15804 37856 15810 37868
rect 16022 37856 16028 37868
rect 15804 37828 16028 37856
rect 15804 37816 15810 37828
rect 16022 37816 16028 37828
rect 16080 37816 16086 37868
rect 16117 37859 16175 37865
rect 16117 37825 16129 37859
rect 16163 37856 16175 37859
rect 16206 37856 16212 37868
rect 16163 37828 16212 37856
rect 16163 37825 16175 37828
rect 16117 37819 16175 37825
rect 16206 37816 16212 37828
rect 16264 37816 16270 37868
rect 13354 37748 13360 37800
rect 13412 37748 13418 37800
rect 13630 37748 13636 37800
rect 13688 37788 13694 37800
rect 16316 37797 16344 37896
rect 16850 37884 16856 37896
rect 16908 37924 16914 37936
rect 17310 37924 17316 37936
rect 16908 37896 17316 37924
rect 16908 37884 16914 37896
rect 17310 37884 17316 37896
rect 17368 37884 17374 37936
rect 17402 37884 17408 37936
rect 17460 37884 17466 37936
rect 17788 37933 17816 37964
rect 17773 37927 17831 37933
rect 17773 37893 17785 37927
rect 17819 37893 17831 37927
rect 17773 37887 17831 37893
rect 18414 37884 18420 37936
rect 18472 37884 18478 37936
rect 19058 37884 19064 37936
rect 19116 37884 19122 37936
rect 20622 37884 20628 37936
rect 20680 37924 20686 37936
rect 21545 37927 21603 37933
rect 21545 37924 21557 37927
rect 20680 37896 21557 37924
rect 20680 37884 20686 37896
rect 21545 37893 21557 37896
rect 21591 37924 21603 37927
rect 21910 37924 21916 37936
rect 21591 37896 21916 37924
rect 21591 37893 21603 37896
rect 21545 37887 21603 37893
rect 21910 37884 21916 37896
rect 21968 37884 21974 37936
rect 22066 37924 22094 37964
rect 28258 37952 28264 38004
rect 28316 37952 28322 38004
rect 29546 37952 29552 38004
rect 29604 37952 29610 38004
rect 35434 37952 35440 38004
rect 35492 37992 35498 38004
rect 35621 37995 35679 38001
rect 35621 37992 35633 37995
rect 35492 37964 35633 37992
rect 35492 37952 35498 37964
rect 35621 37961 35633 37964
rect 35667 37961 35679 37995
rect 35621 37955 35679 37961
rect 35989 37995 36047 38001
rect 35989 37961 36001 37995
rect 36035 37992 36047 37995
rect 37182 37992 37188 38004
rect 36035 37964 37188 37992
rect 36035 37961 36047 37964
rect 35989 37955 36047 37961
rect 37182 37952 37188 37964
rect 37240 37952 37246 38004
rect 39666 37952 39672 38004
rect 39724 37992 39730 38004
rect 39945 37995 40003 38001
rect 39945 37992 39957 37995
rect 39724 37964 39957 37992
rect 39724 37952 39730 37964
rect 39945 37961 39957 37964
rect 39991 37961 40003 37995
rect 39945 37955 40003 37961
rect 40310 37952 40316 38004
rect 40368 37952 40374 38004
rect 41141 37995 41199 38001
rect 41141 37961 41153 37995
rect 41187 37992 41199 37995
rect 41322 37992 41328 38004
rect 41187 37964 41328 37992
rect 41187 37961 41199 37964
rect 41141 37955 41199 37961
rect 41322 37952 41328 37964
rect 41380 37952 41386 38004
rect 26418 37924 26424 37936
rect 22066 37896 26424 37924
rect 26418 37884 26424 37896
rect 26476 37884 26482 37936
rect 34790 37924 34796 37936
rect 27540 37896 34796 37924
rect 18322 37816 18328 37868
rect 18380 37816 18386 37868
rect 16301 37791 16359 37797
rect 16301 37788 16313 37791
rect 13688 37760 16313 37788
rect 13688 37748 13694 37760
rect 16301 37757 16313 37760
rect 16347 37757 16359 37791
rect 16301 37751 16359 37757
rect 16574 37748 16580 37800
rect 16632 37788 16638 37800
rect 17221 37791 17279 37797
rect 17221 37788 17233 37791
rect 16632 37760 17233 37788
rect 16632 37748 16638 37760
rect 17221 37757 17233 37760
rect 17267 37757 17279 37791
rect 17221 37751 17279 37757
rect 18138 37748 18144 37800
rect 18196 37788 18202 37800
rect 18509 37791 18567 37797
rect 18509 37788 18521 37791
rect 18196 37760 18521 37788
rect 18196 37748 18202 37760
rect 18509 37757 18521 37760
rect 18555 37757 18567 37791
rect 18509 37751 18567 37757
rect 18785 37791 18843 37797
rect 18785 37757 18797 37791
rect 18831 37757 18843 37791
rect 18785 37751 18843 37757
rect 15105 37723 15163 37729
rect 15105 37689 15117 37723
rect 15151 37720 15163 37723
rect 18690 37720 18696 37732
rect 15151 37692 18696 37720
rect 15151 37689 15163 37692
rect 15105 37683 15163 37689
rect 18690 37680 18696 37692
rect 18748 37680 18754 37732
rect 17586 37612 17592 37664
rect 17644 37652 17650 37664
rect 17957 37655 18015 37661
rect 17957 37652 17969 37655
rect 17644 37624 17969 37652
rect 17644 37612 17650 37624
rect 17957 37621 17969 37624
rect 18003 37621 18015 37655
rect 18800 37652 18828 37751
rect 20070 37748 20076 37800
rect 20128 37788 20134 37800
rect 20180 37788 20208 37842
rect 20530 37816 20536 37868
rect 20588 37856 20594 37868
rect 20990 37856 20996 37868
rect 20588 37828 20996 37856
rect 20588 37816 20594 37828
rect 20990 37816 20996 37828
rect 21048 37816 21054 37868
rect 21174 37816 21180 37868
rect 21232 37816 21238 37868
rect 21266 37816 21272 37868
rect 21324 37816 21330 37868
rect 25409 37859 25467 37865
rect 25409 37825 25421 37859
rect 25455 37856 25467 37859
rect 25498 37856 25504 37868
rect 25455 37828 25504 37856
rect 25455 37825 25467 37828
rect 25409 37819 25467 37825
rect 25498 37816 25504 37828
rect 25556 37816 25562 37868
rect 27154 37816 27160 37868
rect 27212 37816 27218 37868
rect 27246 37816 27252 37868
rect 27304 37816 27310 37868
rect 21450 37788 21456 37800
rect 20128 37760 21456 37788
rect 20128 37748 20134 37760
rect 21450 37748 21456 37760
rect 21508 37748 21514 37800
rect 21637 37791 21695 37797
rect 21637 37757 21649 37791
rect 21683 37788 21695 37791
rect 22465 37791 22523 37797
rect 22465 37788 22477 37791
rect 21683 37760 22477 37788
rect 21683 37757 21695 37760
rect 21637 37751 21695 37757
rect 22465 37757 22477 37760
rect 22511 37757 22523 37791
rect 22465 37751 22523 37757
rect 23014 37748 23020 37800
rect 23072 37748 23078 37800
rect 27540 37797 27568 37896
rect 34790 37884 34796 37896
rect 34848 37884 34854 37936
rect 40681 37927 40739 37933
rect 40681 37893 40693 37927
rect 40727 37924 40739 37927
rect 40862 37924 40868 37936
rect 40727 37896 40868 37924
rect 40727 37893 40739 37896
rect 40681 37887 40739 37893
rect 40862 37884 40868 37896
rect 40920 37924 40926 37936
rect 41601 37927 41659 37933
rect 41601 37924 41613 37927
rect 40920 37896 41613 37924
rect 40920 37884 40926 37896
rect 41601 37893 41613 37896
rect 41647 37893 41659 37927
rect 41601 37887 41659 37893
rect 28077 37859 28135 37865
rect 28077 37825 28089 37859
rect 28123 37825 28135 37859
rect 28077 37819 28135 37825
rect 27525 37791 27583 37797
rect 27525 37757 27537 37791
rect 27571 37757 27583 37791
rect 27525 37751 27583 37757
rect 27617 37791 27675 37797
rect 27617 37757 27629 37791
rect 27663 37788 27675 37791
rect 27890 37788 27896 37800
rect 27663 37760 27896 37788
rect 27663 37757 27675 37760
rect 27617 37751 27675 37757
rect 20806 37680 20812 37732
rect 20864 37720 20870 37732
rect 27540 37720 27568 37751
rect 27890 37748 27896 37760
rect 27948 37748 27954 37800
rect 20864 37692 27568 37720
rect 20864 37680 20870 37692
rect 19426 37652 19432 37664
rect 18800 37624 19432 37652
rect 17957 37615 18015 37621
rect 19426 37612 19432 37624
rect 19484 37612 19490 37664
rect 20530 37612 20536 37664
rect 20588 37612 20594 37664
rect 20898 37612 20904 37664
rect 20956 37652 20962 37664
rect 20993 37655 21051 37661
rect 20993 37652 21005 37655
rect 20956 37624 21005 37652
rect 20956 37612 20962 37624
rect 20993 37621 21005 37624
rect 21039 37621 21051 37655
rect 20993 37615 21051 37621
rect 23658 37612 23664 37664
rect 23716 37652 23722 37664
rect 24762 37652 24768 37664
rect 23716 37624 24768 37652
rect 23716 37612 23722 37624
rect 24762 37612 24768 37624
rect 24820 37652 24826 37664
rect 25317 37655 25375 37661
rect 25317 37652 25329 37655
rect 24820 37624 25329 37652
rect 24820 37612 24826 37624
rect 25317 37621 25329 37624
rect 25363 37621 25375 37655
rect 25317 37615 25375 37621
rect 26510 37612 26516 37664
rect 26568 37652 26574 37664
rect 26973 37655 27031 37661
rect 26973 37652 26985 37655
rect 26568 37624 26985 37652
rect 26568 37612 26574 37624
rect 26973 37621 26985 37624
rect 27019 37621 27031 37655
rect 26973 37615 27031 37621
rect 27614 37612 27620 37664
rect 27672 37652 27678 37664
rect 27801 37655 27859 37661
rect 27801 37652 27813 37655
rect 27672 37624 27813 37652
rect 27672 37612 27678 37624
rect 27801 37621 27813 37624
rect 27847 37621 27859 37655
rect 28092 37652 28120 37819
rect 28534 37816 28540 37868
rect 28592 37816 28598 37868
rect 29457 37859 29515 37865
rect 29457 37825 29469 37859
rect 29503 37856 29515 37859
rect 29917 37859 29975 37865
rect 29917 37856 29929 37859
rect 29503 37828 29929 37856
rect 29503 37825 29515 37828
rect 29457 37819 29515 37825
rect 29917 37825 29929 37828
rect 29963 37825 29975 37859
rect 29917 37819 29975 37825
rect 33781 37859 33839 37865
rect 33781 37825 33793 37859
rect 33827 37856 33839 37859
rect 33962 37856 33968 37868
rect 33827 37828 33968 37856
rect 33827 37825 33839 37828
rect 33781 37819 33839 37825
rect 33962 37816 33968 37828
rect 34020 37816 34026 37868
rect 35986 37816 35992 37868
rect 36044 37856 36050 37868
rect 36081 37859 36139 37865
rect 36081 37856 36093 37859
rect 36044 37828 36093 37856
rect 36044 37816 36050 37828
rect 36081 37825 36093 37828
rect 36127 37825 36139 37859
rect 36081 37819 36139 37825
rect 37826 37816 37832 37868
rect 37884 37816 37890 37868
rect 39945 37859 40003 37865
rect 39945 37825 39957 37859
rect 39991 37856 40003 37859
rect 40034 37856 40040 37868
rect 39991 37828 40040 37856
rect 39991 37825 40003 37828
rect 39945 37819 40003 37825
rect 40034 37816 40040 37828
rect 40092 37816 40098 37868
rect 40126 37816 40132 37868
rect 40184 37816 40190 37868
rect 40773 37859 40831 37865
rect 40773 37825 40785 37859
rect 40819 37856 40831 37859
rect 41138 37856 41144 37868
rect 40819 37828 41144 37856
rect 40819 37825 40831 37828
rect 40773 37819 40831 37825
rect 41138 37816 41144 37828
rect 41196 37856 41202 37868
rect 41509 37859 41567 37865
rect 41509 37856 41521 37859
rect 41196 37828 41521 37856
rect 41196 37816 41202 37828
rect 41509 37825 41521 37828
rect 41555 37825 41567 37859
rect 41509 37819 41567 37825
rect 28261 37791 28319 37797
rect 28261 37757 28273 37791
rect 28307 37788 28319 37791
rect 28810 37788 28816 37800
rect 28307 37760 28816 37788
rect 28307 37757 28319 37760
rect 28261 37751 28319 37757
rect 28810 37748 28816 37760
rect 28868 37748 28874 37800
rect 28994 37748 29000 37800
rect 29052 37788 29058 37800
rect 29641 37791 29699 37797
rect 29641 37788 29653 37791
rect 29052 37760 29653 37788
rect 29052 37748 29058 37760
rect 29641 37757 29653 37760
rect 29687 37757 29699 37791
rect 29641 37751 29699 37757
rect 30466 37748 30472 37800
rect 30524 37748 30530 37800
rect 34146 37748 34152 37800
rect 34204 37788 34210 37800
rect 36173 37791 36231 37797
rect 36173 37788 36185 37791
rect 34204 37760 36185 37788
rect 34204 37748 34210 37760
rect 36173 37757 36185 37760
rect 36219 37757 36231 37791
rect 36173 37751 36231 37757
rect 37921 37791 37979 37797
rect 37921 37757 37933 37791
rect 37967 37788 37979 37791
rect 38105 37791 38163 37797
rect 38105 37788 38117 37791
rect 37967 37760 38117 37788
rect 37967 37757 37979 37760
rect 37921 37751 37979 37757
rect 38105 37757 38117 37760
rect 38151 37757 38163 37791
rect 38105 37751 38163 37757
rect 38562 37748 38568 37800
rect 38620 37748 38626 37800
rect 39850 37748 39856 37800
rect 39908 37788 39914 37800
rect 40865 37791 40923 37797
rect 40865 37788 40877 37791
rect 39908 37760 40877 37788
rect 39908 37748 39914 37760
rect 40865 37757 40877 37760
rect 40911 37788 40923 37791
rect 41690 37788 41696 37800
rect 40911 37760 41696 37788
rect 40911 37757 40923 37760
rect 40865 37751 40923 37757
rect 41690 37748 41696 37760
rect 41748 37748 41754 37800
rect 28445 37723 28503 37729
rect 28445 37689 28457 37723
rect 28491 37720 28503 37723
rect 28626 37720 28632 37732
rect 28491 37692 28632 37720
rect 28491 37689 28503 37692
rect 28445 37683 28503 37689
rect 28626 37680 28632 37692
rect 28684 37680 28690 37732
rect 30742 37720 30748 37732
rect 28736 37692 30748 37720
rect 28736 37652 28764 37692
rect 30742 37680 30748 37692
rect 30800 37680 30806 37732
rect 35066 37680 35072 37732
rect 35124 37720 35130 37732
rect 37461 37723 37519 37729
rect 37461 37720 37473 37723
rect 35124 37692 37473 37720
rect 35124 37680 35130 37692
rect 37461 37689 37473 37692
rect 37507 37689 37519 37723
rect 37461 37683 37519 37689
rect 38289 37723 38347 37729
rect 38289 37689 38301 37723
rect 38335 37720 38347 37723
rect 38654 37720 38660 37732
rect 38335 37692 38660 37720
rect 38335 37689 38347 37692
rect 38289 37683 38347 37689
rect 38654 37680 38660 37692
rect 38712 37680 38718 37732
rect 28092 37624 28764 37652
rect 27801 37615 27859 37621
rect 28810 37612 28816 37664
rect 28868 37652 28874 37664
rect 29089 37655 29147 37661
rect 29089 37652 29101 37655
rect 28868 37624 29101 37652
rect 28868 37612 28874 37624
rect 29089 37621 29101 37624
rect 29135 37621 29147 37655
rect 29089 37615 29147 37621
rect 33594 37612 33600 37664
rect 33652 37652 33658 37664
rect 35250 37652 35256 37664
rect 33652 37624 35256 37652
rect 33652 37612 33658 37624
rect 35250 37612 35256 37624
rect 35308 37612 35314 37664
rect 1104 37562 42504 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 42504 37562
rect 1104 37488 42504 37510
rect 16206 37408 16212 37460
rect 16264 37408 16270 37460
rect 17037 37451 17095 37457
rect 17037 37417 17049 37451
rect 17083 37448 17095 37451
rect 17126 37448 17132 37460
rect 17083 37420 17132 37448
rect 17083 37417 17095 37420
rect 17037 37411 17095 37417
rect 17126 37408 17132 37420
rect 17184 37408 17190 37460
rect 17402 37408 17408 37460
rect 17460 37408 17466 37460
rect 18322 37408 18328 37460
rect 18380 37448 18386 37460
rect 19245 37451 19303 37457
rect 19245 37448 19257 37451
rect 18380 37420 19257 37448
rect 18380 37408 18386 37420
rect 19245 37417 19257 37420
rect 19291 37417 19303 37451
rect 19245 37411 19303 37417
rect 22373 37451 22431 37457
rect 22373 37417 22385 37451
rect 22419 37448 22431 37451
rect 22462 37448 22468 37460
rect 22419 37420 22468 37448
rect 22419 37417 22431 37420
rect 22373 37411 22431 37417
rect 22462 37408 22468 37420
rect 22520 37448 22526 37460
rect 23014 37448 23020 37460
rect 22520 37420 23020 37448
rect 22520 37408 22526 37420
rect 23014 37408 23020 37420
rect 23072 37408 23078 37460
rect 27062 37448 27068 37460
rect 26252 37420 27068 37448
rect 15657 37315 15715 37321
rect 15657 37281 15669 37315
rect 15703 37312 15715 37315
rect 16485 37315 16543 37321
rect 16485 37312 16497 37315
rect 15703 37284 16497 37312
rect 15703 37281 15715 37284
rect 15657 37275 15715 37281
rect 16485 37281 16497 37284
rect 16531 37312 16543 37315
rect 17420 37312 17448 37408
rect 19518 37340 19524 37392
rect 19576 37380 19582 37392
rect 19978 37380 19984 37392
rect 19576 37352 19984 37380
rect 19576 37340 19582 37352
rect 19978 37340 19984 37352
rect 20036 37340 20042 37392
rect 16531 37284 17448 37312
rect 16531 37281 16543 37284
rect 16485 37275 16543 37281
rect 17586 37272 17592 37324
rect 17644 37272 17650 37324
rect 19426 37272 19432 37324
rect 19484 37312 19490 37324
rect 20625 37315 20683 37321
rect 20625 37312 20637 37315
rect 19484 37284 20637 37312
rect 19484 37272 19490 37284
rect 20625 37281 20637 37284
rect 20671 37281 20683 37315
rect 20625 37275 20683 37281
rect 20898 37272 20904 37324
rect 20956 37272 20962 37324
rect 23014 37272 23020 37324
rect 23072 37272 23078 37324
rect 24762 37272 24768 37324
rect 24820 37272 24826 37324
rect 24854 37272 24860 37324
rect 24912 37272 24918 37324
rect 26252 37321 26280 37420
rect 27062 37408 27068 37420
rect 27120 37408 27126 37460
rect 24949 37315 25007 37321
rect 24949 37281 24961 37315
rect 24995 37281 25007 37315
rect 24949 37275 25007 37281
rect 26237 37315 26295 37321
rect 26237 37281 26249 37315
rect 26283 37281 26295 37315
rect 26237 37275 26295 37281
rect 12894 37204 12900 37256
rect 12952 37244 12958 37256
rect 13265 37247 13323 37253
rect 13265 37244 13277 37247
rect 12952 37216 13277 37244
rect 12952 37204 12958 37216
rect 13265 37213 13277 37216
rect 13311 37244 13323 37247
rect 13354 37244 13360 37256
rect 13311 37216 13360 37244
rect 13311 37213 13323 37216
rect 13265 37207 13323 37213
rect 13354 37204 13360 37216
rect 13412 37244 13418 37256
rect 14826 37244 14832 37256
rect 13412 37216 14832 37244
rect 13412 37204 13418 37216
rect 14826 37204 14832 37216
rect 14884 37204 14890 37256
rect 16574 37204 16580 37256
rect 16632 37204 16638 37256
rect 17126 37204 17132 37256
rect 17184 37244 17190 37256
rect 17313 37247 17371 37253
rect 17313 37244 17325 37247
rect 17184 37216 17325 37244
rect 17184 37204 17190 37216
rect 17313 37213 17325 37216
rect 17359 37213 17371 37247
rect 17313 37207 17371 37213
rect 19518 37204 19524 37256
rect 19576 37244 19582 37256
rect 19797 37247 19855 37253
rect 19797 37244 19809 37247
rect 19576 37216 19809 37244
rect 19576 37204 19582 37216
rect 19797 37213 19809 37216
rect 19843 37244 19855 37247
rect 20162 37244 20168 37256
rect 19843 37216 20168 37244
rect 19843 37213 19855 37216
rect 19797 37207 19855 37213
rect 20162 37204 20168 37216
rect 20220 37204 20226 37256
rect 20257 37247 20315 37253
rect 20257 37213 20269 37247
rect 20303 37213 20315 37247
rect 24780 37244 24808 37272
rect 24964 37244 24992 37275
rect 26510 37272 26516 37324
rect 26568 37272 26574 37324
rect 32030 37272 32036 37324
rect 32088 37272 32094 37324
rect 33686 37272 33692 37324
rect 33744 37312 33750 37324
rect 33962 37312 33968 37324
rect 33744 37284 33968 37312
rect 33744 37272 33750 37284
rect 33962 37272 33968 37284
rect 34020 37272 34026 37324
rect 34146 37272 34152 37324
rect 34204 37272 34210 37324
rect 34790 37272 34796 37324
rect 34848 37312 34854 37324
rect 34848 37284 35296 37312
rect 34848 37272 34854 37284
rect 35268 37256 35296 37284
rect 24780 37216 24992 37244
rect 20257 37207 20315 37213
rect 14093 37179 14151 37185
rect 14093 37145 14105 37179
rect 14139 37176 14151 37179
rect 15102 37176 15108 37188
rect 14139 37148 15108 37176
rect 14139 37145 14151 37148
rect 14093 37139 14151 37145
rect 15102 37136 15108 37148
rect 15160 37136 15166 37188
rect 15749 37179 15807 37185
rect 15749 37145 15761 37179
rect 15795 37176 15807 37179
rect 16592 37176 16620 37204
rect 16669 37179 16727 37185
rect 16669 37176 16681 37179
rect 15795 37148 16681 37176
rect 15795 37145 15807 37148
rect 15749 37139 15807 37145
rect 16669 37145 16681 37148
rect 16715 37145 16727 37179
rect 20070 37176 20076 37188
rect 18814 37148 20076 37176
rect 16669 37139 16727 37145
rect 20070 37136 20076 37148
rect 20128 37136 20134 37188
rect 15841 37111 15899 37117
rect 15841 37077 15853 37111
rect 15887 37108 15899 37111
rect 16022 37108 16028 37120
rect 15887 37080 16028 37108
rect 15887 37077 15899 37080
rect 15841 37071 15899 37077
rect 16022 37068 16028 37080
rect 16080 37108 16086 37120
rect 16577 37111 16635 37117
rect 16577 37108 16589 37111
rect 16080 37080 16589 37108
rect 16080 37068 16086 37080
rect 16577 37077 16589 37080
rect 16623 37077 16635 37111
rect 16577 37071 16635 37077
rect 19061 37111 19119 37117
rect 19061 37077 19073 37111
rect 19107 37108 19119 37111
rect 19518 37108 19524 37120
rect 19107 37080 19524 37108
rect 19107 37077 19119 37080
rect 19061 37071 19119 37077
rect 19518 37068 19524 37080
rect 19576 37068 19582 37120
rect 19886 37068 19892 37120
rect 19944 37108 19950 37120
rect 20272 37108 20300 37207
rect 25038 37204 25044 37256
rect 25096 37244 25102 37256
rect 25682 37244 25688 37256
rect 25096 37216 25688 37244
rect 25096 37204 25102 37216
rect 25682 37204 25688 37216
rect 25740 37244 25746 37256
rect 25777 37247 25835 37253
rect 25777 37244 25789 37247
rect 25740 37216 25789 37244
rect 25740 37204 25746 37216
rect 25777 37213 25789 37216
rect 25823 37213 25835 37247
rect 25777 37207 25835 37213
rect 27614 37204 27620 37256
rect 27672 37204 27678 37256
rect 30650 37204 30656 37256
rect 30708 37244 30714 37256
rect 30837 37247 30895 37253
rect 30837 37244 30849 37247
rect 30708 37216 30849 37244
rect 30708 37204 30714 37216
rect 30837 37213 30849 37216
rect 30883 37213 30895 37247
rect 30837 37207 30895 37213
rect 31021 37247 31079 37253
rect 31021 37213 31033 37247
rect 31067 37244 31079 37247
rect 31110 37244 31116 37256
rect 31067 37216 31116 37244
rect 31067 37213 31079 37216
rect 31021 37207 31079 37213
rect 31110 37204 31116 37216
rect 31168 37204 31174 37256
rect 31202 37204 31208 37256
rect 31260 37244 31266 37256
rect 31297 37247 31355 37253
rect 31297 37244 31309 37247
rect 31260 37216 31309 37244
rect 31260 37204 31266 37216
rect 31297 37213 31309 37216
rect 31343 37213 31355 37247
rect 31297 37207 31355 37213
rect 31478 37204 31484 37256
rect 31536 37204 31542 37256
rect 32125 37247 32183 37253
rect 32125 37213 32137 37247
rect 32171 37244 32183 37247
rect 34974 37244 34980 37256
rect 32171 37216 34980 37244
rect 32171 37213 32183 37216
rect 32125 37207 32183 37213
rect 34974 37204 34980 37216
rect 35032 37204 35038 37256
rect 35069 37247 35127 37253
rect 35069 37213 35081 37247
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 20349 37179 20407 37185
rect 20349 37145 20361 37179
rect 20395 37176 20407 37179
rect 20806 37176 20812 37188
rect 20395 37148 20812 37176
rect 20395 37145 20407 37148
rect 20349 37139 20407 37145
rect 20806 37136 20812 37148
rect 20864 37136 20870 37188
rect 21450 37136 21456 37188
rect 21508 37136 21514 37188
rect 23109 37179 23167 37185
rect 23109 37145 23121 37179
rect 23155 37176 23167 37179
rect 30374 37176 30380 37188
rect 23155 37148 26924 37176
rect 23155 37145 23167 37148
rect 23109 37139 23167 37145
rect 20714 37108 20720 37120
rect 19944 37080 20720 37108
rect 19944 37068 19950 37080
rect 20714 37068 20720 37080
rect 20772 37108 20778 37120
rect 23014 37108 23020 37120
rect 20772 37080 23020 37108
rect 20772 37068 20778 37080
rect 23014 37068 23020 37080
rect 23072 37068 23078 37120
rect 23198 37068 23204 37120
rect 23256 37068 23262 37120
rect 23382 37068 23388 37120
rect 23440 37108 23446 37120
rect 23569 37111 23627 37117
rect 23569 37108 23581 37111
rect 23440 37080 23581 37108
rect 23440 37068 23446 37080
rect 23569 37077 23581 37080
rect 23615 37077 23627 37111
rect 23569 37071 23627 37077
rect 23658 37068 23664 37120
rect 23716 37108 23722 37120
rect 24397 37111 24455 37117
rect 24397 37108 24409 37111
rect 23716 37080 24409 37108
rect 23716 37068 23722 37080
rect 24397 37077 24409 37080
rect 24443 37077 24455 37111
rect 24397 37071 24455 37077
rect 24765 37111 24823 37117
rect 24765 37077 24777 37111
rect 24811 37108 24823 37111
rect 25225 37111 25283 37117
rect 25225 37108 25237 37111
rect 24811 37080 25237 37108
rect 24811 37077 24823 37080
rect 24765 37071 24823 37077
rect 25225 37077 25237 37080
rect 25271 37077 25283 37111
rect 26896 37108 26924 37148
rect 27816 37148 30380 37176
rect 27816 37108 27844 37148
rect 30374 37136 30380 37148
rect 30432 37136 30438 37188
rect 31754 37136 31760 37188
rect 31812 37176 31818 37188
rect 32766 37176 32772 37188
rect 31812 37148 32772 37176
rect 31812 37136 31818 37148
rect 32766 37136 32772 37148
rect 32824 37176 32830 37188
rect 32861 37179 32919 37185
rect 32861 37176 32873 37179
rect 32824 37148 32873 37176
rect 32824 37136 32830 37148
rect 32861 37145 32873 37148
rect 32907 37145 32919 37179
rect 32861 37139 32919 37145
rect 33962 37136 33968 37188
rect 34020 37136 34026 37188
rect 35084 37176 35112 37207
rect 35250 37204 35256 37256
rect 35308 37204 35314 37256
rect 37369 37247 37427 37253
rect 37369 37213 37381 37247
rect 37415 37244 37427 37247
rect 37458 37244 37464 37256
rect 37415 37216 37464 37244
rect 37415 37213 37427 37216
rect 37369 37207 37427 37213
rect 37458 37204 37464 37216
rect 37516 37204 37522 37256
rect 37553 37247 37611 37253
rect 37553 37213 37565 37247
rect 37599 37244 37611 37247
rect 37642 37244 37648 37256
rect 37599 37216 37648 37244
rect 37599 37213 37611 37216
rect 37553 37207 37611 37213
rect 37642 37204 37648 37216
rect 37700 37244 37706 37256
rect 37918 37244 37924 37256
rect 37700 37216 37924 37244
rect 37700 37204 37706 37216
rect 37918 37204 37924 37216
rect 37976 37204 37982 37256
rect 42150 37204 42156 37256
rect 42208 37204 42214 37256
rect 35342 37176 35348 37188
rect 35084 37148 35348 37176
rect 35342 37136 35348 37148
rect 35400 37136 35406 37188
rect 26896 37080 27844 37108
rect 25225 37071 25283 37077
rect 27890 37068 27896 37120
rect 27948 37108 27954 37120
rect 27985 37111 28043 37117
rect 27985 37108 27997 37111
rect 27948 37080 27997 37108
rect 27948 37068 27954 37080
rect 27985 37077 27997 37080
rect 28031 37077 28043 37111
rect 27985 37071 28043 37077
rect 30929 37111 30987 37117
rect 30929 37077 30941 37111
rect 30975 37108 30987 37111
rect 31294 37108 31300 37120
rect 30975 37080 31300 37108
rect 30975 37077 30987 37080
rect 30929 37071 30987 37077
rect 31294 37068 31300 37080
rect 31352 37068 31358 37120
rect 31389 37111 31447 37117
rect 31389 37077 31401 37111
rect 31435 37108 31447 37111
rect 31570 37108 31576 37120
rect 31435 37080 31576 37108
rect 31435 37077 31447 37080
rect 31389 37071 31447 37077
rect 31570 37068 31576 37080
rect 31628 37068 31634 37120
rect 32490 37068 32496 37120
rect 32548 37068 32554 37120
rect 35253 37111 35311 37117
rect 35253 37077 35265 37111
rect 35299 37108 35311 37111
rect 36354 37108 36360 37120
rect 35299 37080 36360 37108
rect 35299 37077 35311 37080
rect 35253 37071 35311 37077
rect 36354 37068 36360 37080
rect 36412 37068 36418 37120
rect 37274 37068 37280 37120
rect 37332 37108 37338 37120
rect 37461 37111 37519 37117
rect 37461 37108 37473 37111
rect 37332 37080 37473 37108
rect 37332 37068 37338 37080
rect 37461 37077 37473 37080
rect 37507 37077 37519 37111
rect 37461 37071 37519 37077
rect 41046 37068 41052 37120
rect 41104 37108 41110 37120
rect 41509 37111 41567 37117
rect 41509 37108 41521 37111
rect 41104 37080 41521 37108
rect 41104 37068 41110 37080
rect 41509 37077 41521 37080
rect 41555 37077 41567 37111
rect 41509 37071 41567 37077
rect 1104 37018 42504 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 42504 37018
rect 1104 36944 42504 36966
rect 3804 36876 7328 36904
rect 3234 36660 3240 36712
rect 3292 36700 3298 36712
rect 3804 36709 3832 36876
rect 7300 36848 7328 36876
rect 17788 36876 20209 36904
rect 5442 36836 5448 36848
rect 5290 36808 5448 36836
rect 5442 36796 5448 36808
rect 5500 36796 5506 36848
rect 7282 36796 7288 36848
rect 7340 36796 7346 36848
rect 8110 36728 8116 36780
rect 8168 36728 8174 36780
rect 15930 36728 15936 36780
rect 15988 36728 15994 36780
rect 16758 36728 16764 36780
rect 16816 36768 16822 36780
rect 17788 36777 17816 36876
rect 19153 36839 19211 36845
rect 19153 36805 19165 36839
rect 19199 36836 19211 36839
rect 20181 36836 20209 36876
rect 20254 36864 20260 36916
rect 20312 36904 20318 36916
rect 20349 36907 20407 36913
rect 20349 36904 20361 36907
rect 20312 36876 20361 36904
rect 20312 36864 20318 36876
rect 20349 36873 20361 36876
rect 20395 36873 20407 36907
rect 20349 36867 20407 36873
rect 23198 36864 23204 36916
rect 23256 36864 23262 36916
rect 23934 36864 23940 36916
rect 23992 36864 23998 36916
rect 25038 36864 25044 36916
rect 25096 36864 25102 36916
rect 25590 36864 25596 36916
rect 25648 36904 25654 36916
rect 25961 36907 26019 36913
rect 25961 36904 25973 36907
rect 25648 36876 25973 36904
rect 25648 36864 25654 36876
rect 25961 36873 25973 36876
rect 26007 36873 26019 36907
rect 28994 36904 29000 36916
rect 25961 36867 26019 36873
rect 27080 36876 29000 36904
rect 22830 36836 22836 36848
rect 19199 36808 19564 36836
rect 20181 36808 22836 36836
rect 19199 36805 19211 36808
rect 19153 36799 19211 36805
rect 17497 36771 17555 36777
rect 17497 36768 17509 36771
rect 16816 36740 17509 36768
rect 16816 36728 16822 36740
rect 17497 36737 17509 36740
rect 17543 36737 17555 36771
rect 17497 36731 17555 36737
rect 17681 36771 17739 36777
rect 17681 36737 17693 36771
rect 17727 36768 17739 36771
rect 17773 36771 17831 36777
rect 17773 36768 17785 36771
rect 17727 36740 17785 36768
rect 17727 36737 17739 36740
rect 17681 36731 17739 36737
rect 17773 36737 17785 36740
rect 17819 36737 17831 36771
rect 17773 36731 17831 36737
rect 18693 36771 18751 36777
rect 18693 36737 18705 36771
rect 18739 36737 18751 36771
rect 18693 36731 18751 36737
rect 3789 36703 3847 36709
rect 3789 36700 3801 36703
rect 3292 36672 3801 36700
rect 3292 36660 3298 36672
rect 3789 36669 3801 36672
rect 3835 36669 3847 36703
rect 3789 36663 3847 36669
rect 4062 36660 4068 36712
rect 4120 36660 4126 36712
rect 15562 36660 15568 36712
rect 15620 36660 15626 36712
rect 16209 36703 16267 36709
rect 16209 36669 16221 36703
rect 16255 36700 16267 36703
rect 16850 36700 16856 36712
rect 16255 36672 16856 36700
rect 16255 36669 16267 36672
rect 16209 36663 16267 36669
rect 16850 36660 16856 36672
rect 16908 36660 16914 36712
rect 17034 36660 17040 36712
rect 17092 36700 17098 36712
rect 17221 36703 17279 36709
rect 17221 36700 17233 36703
rect 17092 36672 17233 36700
rect 17092 36660 17098 36672
rect 17221 36669 17233 36672
rect 17267 36700 17279 36703
rect 18708 36700 18736 36731
rect 18782 36728 18788 36780
rect 18840 36728 18846 36780
rect 18969 36771 19027 36777
rect 18969 36737 18981 36771
rect 19015 36768 19027 36771
rect 19058 36768 19064 36780
rect 19015 36740 19064 36768
rect 19015 36737 19027 36740
rect 18969 36731 19027 36737
rect 19058 36728 19064 36740
rect 19116 36728 19122 36780
rect 19536 36777 19564 36808
rect 22830 36796 22836 36808
rect 22888 36796 22894 36848
rect 23474 36836 23480 36848
rect 23308 36808 23480 36836
rect 19429 36771 19487 36777
rect 19429 36737 19441 36771
rect 19475 36737 19487 36771
rect 19429 36731 19487 36737
rect 19521 36771 19579 36777
rect 19521 36737 19533 36771
rect 19567 36737 19579 36771
rect 19521 36731 19579 36737
rect 19797 36771 19855 36777
rect 19797 36737 19809 36771
rect 19843 36768 19855 36771
rect 19886 36768 19892 36780
rect 19843 36740 19892 36768
rect 19843 36737 19855 36740
rect 19797 36731 19855 36737
rect 17267 36672 18736 36700
rect 17267 36669 17279 36672
rect 17221 36663 17279 36669
rect 16117 36635 16175 36641
rect 16117 36601 16129 36635
rect 16163 36632 16175 36635
rect 16163 36604 17264 36632
rect 16163 36601 16175 36604
rect 16117 36595 16175 36601
rect 17236 36576 17264 36604
rect 18138 36592 18144 36644
rect 18196 36632 18202 36644
rect 19334 36632 19340 36644
rect 18196 36604 19340 36632
rect 18196 36592 18202 36604
rect 19334 36592 19340 36604
rect 19392 36592 19398 36644
rect 19444 36632 19472 36731
rect 19886 36728 19892 36740
rect 19944 36728 19950 36780
rect 20257 36771 20315 36777
rect 20257 36737 20269 36771
rect 20303 36737 20315 36771
rect 20257 36731 20315 36737
rect 20717 36771 20775 36777
rect 20717 36737 20729 36771
rect 20763 36768 20775 36771
rect 21358 36768 21364 36780
rect 20763 36740 21364 36768
rect 20763 36737 20775 36740
rect 20717 36731 20775 36737
rect 19610 36632 19616 36644
rect 19444 36604 19616 36632
rect 19610 36592 19616 36604
rect 19668 36592 19674 36644
rect 20272 36632 20300 36731
rect 21358 36728 21364 36740
rect 21416 36728 21422 36780
rect 23308 36777 23336 36808
rect 23474 36796 23480 36808
rect 23532 36796 23538 36848
rect 23569 36839 23627 36845
rect 23569 36805 23581 36839
rect 23615 36836 23627 36839
rect 23658 36836 23664 36848
rect 23615 36808 23664 36836
rect 23615 36805 23627 36808
rect 23569 36799 23627 36805
rect 23658 36796 23664 36808
rect 23716 36796 23722 36848
rect 23952 36836 23980 36864
rect 23952 36808 24058 36836
rect 23293 36771 23351 36777
rect 23293 36737 23305 36771
rect 23339 36737 23351 36771
rect 23293 36731 23351 36737
rect 25869 36771 25927 36777
rect 25869 36737 25881 36771
rect 25915 36768 25927 36771
rect 26973 36771 27031 36777
rect 26973 36768 26985 36771
rect 25915 36740 26985 36768
rect 25915 36737 25927 36740
rect 25869 36731 25927 36737
rect 26973 36737 26985 36740
rect 27019 36737 27031 36771
rect 26973 36731 27031 36737
rect 20806 36660 20812 36712
rect 20864 36660 20870 36712
rect 20993 36703 21051 36709
rect 20993 36669 21005 36703
rect 21039 36700 21051 36703
rect 21174 36700 21180 36712
rect 21039 36672 21180 36700
rect 21039 36669 21051 36672
rect 20993 36663 21051 36669
rect 21174 36660 21180 36672
rect 21232 36660 21238 36712
rect 22646 36660 22652 36712
rect 22704 36660 22710 36712
rect 23014 36660 23020 36712
rect 23072 36700 23078 36712
rect 26145 36703 26203 36709
rect 26145 36700 26157 36703
rect 23072 36672 26157 36700
rect 23072 36660 23078 36672
rect 26145 36669 26157 36672
rect 26191 36700 26203 36703
rect 27080 36700 27108 36876
rect 28994 36864 29000 36876
rect 29052 36864 29058 36916
rect 31297 36907 31355 36913
rect 31297 36873 31309 36907
rect 31343 36904 31355 36907
rect 31386 36904 31392 36916
rect 31343 36876 31392 36904
rect 31343 36873 31355 36876
rect 31297 36867 31355 36873
rect 31386 36864 31392 36876
rect 31444 36864 31450 36916
rect 31941 36907 31999 36913
rect 31941 36873 31953 36907
rect 31987 36904 31999 36907
rect 32030 36904 32036 36916
rect 31987 36876 32036 36904
rect 31987 36873 31999 36876
rect 31941 36867 31999 36873
rect 32030 36864 32036 36876
rect 32088 36864 32094 36916
rect 33686 36904 33692 36916
rect 32140 36876 33692 36904
rect 29086 36836 29092 36848
rect 28552 36808 29092 36836
rect 28552 36777 28580 36808
rect 29086 36796 29092 36808
rect 29144 36796 29150 36848
rect 30561 36839 30619 36845
rect 30561 36805 30573 36839
rect 30607 36836 30619 36839
rect 31478 36836 31484 36848
rect 30607 36808 30880 36836
rect 30607 36805 30619 36808
rect 30561 36799 30619 36805
rect 28537 36771 28595 36777
rect 28537 36737 28549 36771
rect 28583 36737 28595 36771
rect 30469 36771 30527 36777
rect 28537 36731 28595 36737
rect 26191 36672 27108 36700
rect 26191 36669 26203 36672
rect 26145 36663 26203 36669
rect 27338 36660 27344 36712
rect 27396 36700 27402 36712
rect 27525 36703 27583 36709
rect 27525 36700 27537 36703
rect 27396 36672 27537 36700
rect 27396 36660 27402 36672
rect 27525 36669 27537 36672
rect 27571 36669 27583 36703
rect 27525 36663 27583 36669
rect 28810 36660 28816 36712
rect 28868 36660 28874 36712
rect 28902 36660 28908 36712
rect 28960 36700 28966 36712
rect 29932 36700 29960 36754
rect 30469 36737 30481 36771
rect 30515 36737 30527 36771
rect 30469 36731 30527 36737
rect 28960 36672 29960 36700
rect 28960 36660 28966 36672
rect 21634 36632 21640 36644
rect 20272 36604 21640 36632
rect 21634 36592 21640 36604
rect 21692 36592 21698 36644
rect 24596 36604 25627 36632
rect 4798 36524 4804 36576
rect 4856 36564 4862 36576
rect 5537 36567 5595 36573
rect 5537 36564 5549 36567
rect 4856 36536 5549 36564
rect 4856 36524 4862 36536
rect 5537 36533 5549 36536
rect 5583 36533 5595 36567
rect 5537 36527 5595 36533
rect 15010 36524 15016 36576
rect 15068 36524 15074 36576
rect 15286 36524 15292 36576
rect 15344 36564 15350 36576
rect 15749 36567 15807 36573
rect 15749 36564 15761 36567
rect 15344 36536 15761 36564
rect 15344 36524 15350 36536
rect 15749 36533 15761 36536
rect 15795 36533 15807 36567
rect 15749 36527 15807 36533
rect 16666 36524 16672 36576
rect 16724 36524 16730 36576
rect 17218 36524 17224 36576
rect 17276 36564 17282 36576
rect 17957 36567 18015 36573
rect 17957 36564 17969 36567
rect 17276 36536 17969 36564
rect 17276 36524 17282 36536
rect 17957 36533 17969 36536
rect 18003 36533 18015 36567
rect 17957 36527 18015 36533
rect 18046 36524 18052 36576
rect 18104 36564 18110 36576
rect 19245 36567 19303 36573
rect 19245 36564 19257 36567
rect 18104 36536 19257 36564
rect 18104 36524 18110 36536
rect 19245 36533 19257 36536
rect 19291 36533 19303 36567
rect 19245 36527 19303 36533
rect 19705 36567 19763 36573
rect 19705 36533 19717 36567
rect 19751 36564 19763 36567
rect 19886 36564 19892 36576
rect 19751 36536 19892 36564
rect 19751 36533 19763 36536
rect 19705 36527 19763 36533
rect 19886 36524 19892 36536
rect 19944 36524 19950 36576
rect 20162 36524 20168 36576
rect 20220 36564 20226 36576
rect 24596 36564 24624 36604
rect 20220 36536 24624 36564
rect 20220 36524 20226 36536
rect 25314 36524 25320 36576
rect 25372 36564 25378 36576
rect 25501 36567 25559 36573
rect 25501 36564 25513 36567
rect 25372 36536 25513 36564
rect 25372 36524 25378 36536
rect 25501 36533 25513 36536
rect 25547 36533 25559 36567
rect 25599 36564 25627 36604
rect 25774 36592 25780 36644
rect 25832 36632 25838 36644
rect 27614 36632 27620 36644
rect 25832 36604 27620 36632
rect 25832 36592 25838 36604
rect 27614 36592 27620 36604
rect 27672 36592 27678 36644
rect 30484 36632 30512 36731
rect 30650 36728 30656 36780
rect 30708 36728 30714 36780
rect 30852 36777 30880 36808
rect 30944 36808 31484 36836
rect 30944 36777 30972 36808
rect 31478 36796 31484 36808
rect 31536 36796 31542 36848
rect 32140 36780 32168 36876
rect 33686 36864 33692 36876
rect 33744 36864 33750 36916
rect 34974 36864 34980 36916
rect 35032 36904 35038 36916
rect 35345 36907 35403 36913
rect 35345 36904 35357 36907
rect 35032 36876 35357 36904
rect 35032 36864 35038 36876
rect 35345 36873 35357 36876
rect 35391 36873 35403 36907
rect 35345 36867 35403 36873
rect 37277 36907 37335 36913
rect 37277 36873 37289 36907
rect 37323 36904 37335 36907
rect 37458 36904 37464 36916
rect 37323 36876 37464 36904
rect 37323 36873 37335 36876
rect 37277 36867 37335 36873
rect 37458 36864 37464 36876
rect 37516 36864 37522 36916
rect 38654 36864 38660 36916
rect 38712 36904 38718 36916
rect 40221 36907 40279 36913
rect 40221 36904 40233 36907
rect 38712 36876 40233 36904
rect 38712 36864 38718 36876
rect 40221 36873 40233 36876
rect 40267 36873 40279 36907
rect 40221 36867 40279 36873
rect 41046 36864 41052 36916
rect 41104 36864 41110 36916
rect 35250 36796 35256 36848
rect 35308 36836 35314 36848
rect 39577 36839 39635 36845
rect 35308 36808 35848 36836
rect 35308 36796 35314 36808
rect 30837 36771 30895 36777
rect 30837 36737 30849 36771
rect 30883 36737 30895 36771
rect 30837 36731 30895 36737
rect 30929 36771 30987 36777
rect 30929 36737 30941 36771
rect 30975 36737 30987 36771
rect 30929 36731 30987 36737
rect 31110 36728 31116 36780
rect 31168 36728 31174 36780
rect 31570 36728 31576 36780
rect 31628 36728 31634 36780
rect 32122 36728 32128 36780
rect 32180 36728 32186 36780
rect 33502 36728 33508 36780
rect 33560 36728 33566 36780
rect 34885 36771 34943 36777
rect 34885 36737 34897 36771
rect 34931 36737 34943 36771
rect 34885 36731 34943 36737
rect 31294 36660 31300 36712
rect 31352 36700 31358 36712
rect 31481 36703 31539 36709
rect 31481 36700 31493 36703
rect 31352 36672 31493 36700
rect 31352 36660 31358 36672
rect 31481 36669 31493 36672
rect 31527 36669 31539 36703
rect 31481 36663 31539 36669
rect 32398 36660 32404 36712
rect 32456 36660 32462 36712
rect 32858 36660 32864 36712
rect 32916 36700 32922 36712
rect 33873 36703 33931 36709
rect 33873 36700 33885 36703
rect 32916 36672 33885 36700
rect 32916 36660 32922 36672
rect 33873 36669 33885 36672
rect 33919 36700 33931 36703
rect 34517 36703 34575 36709
rect 34517 36700 34529 36703
rect 33919 36672 34529 36700
rect 33919 36669 33931 36672
rect 33873 36663 33931 36669
rect 34517 36669 34529 36672
rect 34563 36669 34575 36703
rect 34517 36663 34575 36669
rect 34790 36660 34796 36712
rect 34848 36660 34854 36712
rect 29840 36604 30512 36632
rect 31021 36635 31079 36641
rect 29840 36564 29868 36604
rect 31021 36601 31033 36635
rect 31067 36632 31079 36635
rect 31202 36632 31208 36644
rect 31067 36604 31208 36632
rect 31067 36601 31079 36604
rect 31021 36595 31079 36601
rect 31202 36592 31208 36604
rect 31260 36632 31266 36644
rect 31260 36604 31754 36632
rect 31260 36592 31266 36604
rect 25599 36536 29868 36564
rect 25501 36527 25559 36533
rect 29914 36524 29920 36576
rect 29972 36564 29978 36576
rect 30285 36567 30343 36573
rect 30285 36564 30297 36567
rect 29972 36536 30297 36564
rect 29972 36524 29978 36536
rect 30285 36533 30297 36536
rect 30331 36564 30343 36567
rect 30466 36564 30472 36576
rect 30331 36536 30472 36564
rect 30331 36533 30343 36536
rect 30285 36527 30343 36533
rect 30466 36524 30472 36536
rect 30524 36524 30530 36576
rect 31726 36564 31754 36604
rect 33778 36564 33784 36576
rect 31726 36536 33784 36564
rect 33778 36524 33784 36536
rect 33836 36524 33842 36576
rect 33962 36524 33968 36576
rect 34020 36524 34026 36576
rect 34900 36564 34928 36731
rect 35342 36728 35348 36780
rect 35400 36768 35406 36780
rect 35820 36777 35848 36808
rect 37476 36808 38056 36836
rect 35529 36771 35587 36777
rect 35529 36768 35541 36771
rect 35400 36740 35541 36768
rect 35400 36728 35406 36740
rect 35529 36737 35541 36740
rect 35575 36737 35587 36771
rect 35529 36731 35587 36737
rect 35805 36771 35863 36777
rect 35805 36737 35817 36771
rect 35851 36737 35863 36771
rect 35805 36731 35863 36737
rect 36354 36728 36360 36780
rect 36412 36728 36418 36780
rect 37366 36728 37372 36780
rect 37424 36768 37430 36780
rect 37476 36777 37504 36808
rect 37461 36771 37519 36777
rect 37461 36768 37473 36771
rect 37424 36740 37473 36768
rect 37424 36728 37430 36740
rect 37461 36737 37473 36740
rect 37507 36737 37519 36771
rect 37461 36731 37519 36737
rect 37642 36728 37648 36780
rect 37700 36728 37706 36780
rect 37737 36771 37795 36777
rect 37737 36737 37749 36771
rect 37783 36768 37795 36771
rect 37783 36740 37872 36768
rect 37783 36737 37795 36740
rect 37737 36731 37795 36737
rect 35621 36703 35679 36709
rect 35621 36669 35633 36703
rect 35667 36700 35679 36703
rect 36446 36700 36452 36712
rect 35667 36672 36452 36700
rect 35667 36669 35679 36672
rect 35621 36663 35679 36669
rect 36446 36660 36452 36672
rect 36504 36660 36510 36712
rect 37844 36700 37872 36740
rect 37918 36728 37924 36780
rect 37976 36728 37982 36780
rect 38028 36777 38056 36808
rect 39577 36805 39589 36839
rect 39623 36836 39635 36839
rect 40037 36839 40095 36845
rect 39623 36808 39988 36836
rect 39623 36805 39635 36808
rect 39577 36799 39635 36805
rect 38013 36771 38071 36777
rect 38013 36737 38025 36771
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 38102 36728 38108 36780
rect 38160 36774 38166 36780
rect 38160 36768 38240 36774
rect 39022 36768 39028 36780
rect 38160 36746 39028 36768
rect 38160 36728 38166 36746
rect 38212 36740 39028 36746
rect 39022 36728 39028 36740
rect 39080 36728 39086 36780
rect 39776 36777 39804 36808
rect 39485 36771 39543 36777
rect 39485 36737 39497 36771
rect 39531 36737 39543 36771
rect 39485 36731 39543 36737
rect 39669 36771 39727 36777
rect 39669 36737 39681 36771
rect 39715 36737 39727 36771
rect 39669 36731 39727 36737
rect 39761 36771 39819 36777
rect 39761 36737 39773 36771
rect 39807 36737 39819 36771
rect 39761 36731 39819 36737
rect 39853 36771 39911 36777
rect 39853 36737 39865 36771
rect 39899 36737 39911 36771
rect 39960 36768 39988 36808
rect 40037 36805 40049 36839
rect 40083 36836 40095 36839
rect 40083 36808 40448 36836
rect 40083 36805 40095 36808
rect 40037 36799 40095 36805
rect 40420 36777 40448 36808
rect 40129 36771 40187 36777
rect 40129 36768 40141 36771
rect 39960 36740 40141 36768
rect 39853 36731 39911 36737
rect 40129 36737 40141 36740
rect 40175 36737 40187 36771
rect 40129 36731 40187 36737
rect 40313 36771 40371 36777
rect 40313 36737 40325 36771
rect 40359 36737 40371 36771
rect 40313 36731 40371 36737
rect 40405 36771 40463 36777
rect 40405 36737 40417 36771
rect 40451 36768 40463 36771
rect 42150 36768 42156 36780
rect 40451 36740 42156 36768
rect 40451 36737 40463 36740
rect 40405 36731 40463 36737
rect 38120 36700 38148 36728
rect 37844 36672 38148 36700
rect 39500 36700 39528 36731
rect 39574 36700 39580 36712
rect 39500 36672 39580 36700
rect 39574 36660 39580 36672
rect 39632 36660 39638 36712
rect 35253 36635 35311 36641
rect 35253 36601 35265 36635
rect 35299 36632 35311 36635
rect 35710 36632 35716 36644
rect 35299 36604 35716 36632
rect 35299 36601 35311 36604
rect 35253 36595 35311 36601
rect 35710 36592 35716 36604
rect 35768 36592 35774 36644
rect 35986 36592 35992 36644
rect 36044 36592 36050 36644
rect 37550 36592 37556 36644
rect 37608 36632 37614 36644
rect 39684 36632 39712 36731
rect 39868 36700 39896 36731
rect 39942 36700 39948 36712
rect 39868 36672 39948 36700
rect 39942 36660 39948 36672
rect 40000 36700 40006 36712
rect 40328 36700 40356 36731
rect 42150 36728 42156 36740
rect 42208 36728 42214 36780
rect 40000 36672 40356 36700
rect 40000 36660 40006 36672
rect 41138 36660 41144 36712
rect 41196 36660 41202 36712
rect 41230 36660 41236 36712
rect 41288 36660 41294 36712
rect 42061 36703 42119 36709
rect 42061 36700 42073 36703
rect 41386 36672 42073 36700
rect 41386 36644 41414 36672
rect 42061 36669 42073 36672
rect 42107 36669 42119 36703
rect 42061 36663 42119 36669
rect 40310 36632 40316 36644
rect 37608 36604 38608 36632
rect 39684 36604 40316 36632
rect 37608 36592 37614 36604
rect 38580 36576 38608 36604
rect 40310 36592 40316 36604
rect 40368 36632 40374 36644
rect 41322 36632 41328 36644
rect 40368 36604 41328 36632
rect 40368 36592 40374 36604
rect 41322 36592 41328 36604
rect 41380 36604 41414 36644
rect 41380 36592 41386 36604
rect 37182 36564 37188 36576
rect 34900 36536 37188 36564
rect 37182 36524 37188 36536
rect 37240 36524 37246 36576
rect 37458 36524 37464 36576
rect 37516 36564 37522 36576
rect 38197 36567 38255 36573
rect 38197 36564 38209 36567
rect 37516 36536 38209 36564
rect 37516 36524 37522 36536
rect 38197 36533 38209 36536
rect 38243 36533 38255 36567
rect 38197 36527 38255 36533
rect 38562 36524 38568 36576
rect 38620 36564 38626 36576
rect 40037 36567 40095 36573
rect 40037 36564 40049 36567
rect 38620 36536 40049 36564
rect 38620 36524 38626 36536
rect 40037 36533 40049 36536
rect 40083 36533 40095 36567
rect 40037 36527 40095 36533
rect 40678 36524 40684 36576
rect 40736 36524 40742 36576
rect 40770 36524 40776 36576
rect 40828 36564 40834 36576
rect 41509 36567 41567 36573
rect 41509 36564 41521 36567
rect 40828 36536 41521 36564
rect 40828 36524 40834 36536
rect 41509 36533 41521 36536
rect 41555 36533 41567 36567
rect 41509 36527 41567 36533
rect 1104 36474 42504 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 42504 36474
rect 1104 36400 42504 36422
rect 3881 36363 3939 36369
rect 3881 36329 3893 36363
rect 3927 36360 3939 36363
rect 4062 36360 4068 36372
rect 3927 36332 4068 36360
rect 3927 36329 3939 36332
rect 3881 36323 3939 36329
rect 4062 36320 4068 36332
rect 4120 36320 4126 36372
rect 13817 36363 13875 36369
rect 13817 36329 13829 36363
rect 13863 36360 13875 36363
rect 13906 36360 13912 36372
rect 13863 36332 13912 36360
rect 13863 36329 13875 36332
rect 13817 36323 13875 36329
rect 13906 36320 13912 36332
rect 13964 36360 13970 36372
rect 13964 36332 16620 36360
rect 13964 36320 13970 36332
rect 4525 36295 4583 36301
rect 4525 36261 4537 36295
rect 4571 36261 4583 36295
rect 4525 36255 4583 36261
rect 3970 36184 3976 36236
rect 4028 36224 4034 36236
rect 4028 36196 4384 36224
rect 4028 36184 4034 36196
rect 3878 36116 3884 36168
rect 3936 36156 3942 36168
rect 4065 36159 4123 36165
rect 4065 36156 4077 36159
rect 3936 36128 4077 36156
rect 3936 36116 3942 36128
rect 4065 36125 4077 36128
rect 4111 36125 4123 36159
rect 4065 36119 4123 36125
rect 4157 36091 4215 36097
rect 4157 36057 4169 36091
rect 4203 36057 4215 36091
rect 4157 36051 4215 36057
rect 4172 36020 4200 36051
rect 4246 36048 4252 36100
rect 4304 36048 4310 36100
rect 4356 36088 4384 36196
rect 4433 36159 4491 36165
rect 4433 36125 4445 36159
rect 4479 36156 4491 36159
rect 4540 36156 4568 36255
rect 4614 36252 4620 36304
rect 4672 36292 4678 36304
rect 5442 36292 5448 36304
rect 4672 36264 5448 36292
rect 4672 36252 4678 36264
rect 5442 36252 5448 36264
rect 5500 36252 5506 36304
rect 7282 36252 7288 36304
rect 7340 36252 7346 36304
rect 16482 36252 16488 36304
rect 16540 36252 16546 36304
rect 16592 36292 16620 36332
rect 16758 36320 16764 36372
rect 16816 36320 16822 36372
rect 16868 36332 18644 36360
rect 16868 36292 16896 36332
rect 16592 36264 16896 36292
rect 18616 36292 18644 36332
rect 19886 36320 19892 36372
rect 19944 36320 19950 36372
rect 20438 36320 20444 36372
rect 20496 36360 20502 36372
rect 20533 36363 20591 36369
rect 20533 36360 20545 36363
rect 20496 36332 20545 36360
rect 20496 36320 20502 36332
rect 20533 36329 20545 36332
rect 20579 36329 20591 36363
rect 25498 36360 25504 36372
rect 20533 36323 20591 36329
rect 22066 36332 25504 36360
rect 22066 36292 22094 36332
rect 25498 36320 25504 36332
rect 25556 36360 25562 36372
rect 30466 36360 30472 36372
rect 25556 36332 28764 36360
rect 25556 36320 25562 36332
rect 18616 36264 22094 36292
rect 7300 36224 7328 36252
rect 10689 36227 10747 36233
rect 10689 36224 10701 36227
rect 4479 36128 4568 36156
rect 4632 36196 4936 36224
rect 4479 36125 4491 36128
rect 4433 36119 4491 36125
rect 4525 36091 4583 36097
rect 4525 36088 4537 36091
rect 4356 36060 4537 36088
rect 4525 36057 4537 36060
rect 4571 36088 4583 36091
rect 4632 36088 4660 36196
rect 4706 36116 4712 36168
rect 4764 36156 4770 36168
rect 4908 36165 4936 36196
rect 6012 36196 6868 36224
rect 7300 36196 10701 36224
rect 6012 36165 6040 36196
rect 4801 36159 4859 36165
rect 4801 36156 4813 36159
rect 4764 36128 4813 36156
rect 4764 36116 4770 36128
rect 4801 36125 4813 36128
rect 4847 36125 4859 36159
rect 4801 36119 4859 36125
rect 4893 36159 4951 36165
rect 4893 36125 4905 36159
rect 4939 36125 4951 36159
rect 4893 36119 4951 36125
rect 5077 36159 5135 36165
rect 5077 36125 5089 36159
rect 5123 36156 5135 36159
rect 5813 36159 5871 36165
rect 5813 36156 5825 36159
rect 5123 36128 5825 36156
rect 5123 36125 5135 36128
rect 5077 36119 5135 36125
rect 5813 36125 5825 36128
rect 5859 36125 5871 36159
rect 5813 36119 5871 36125
rect 5997 36159 6055 36165
rect 5997 36125 6009 36159
rect 6043 36125 6055 36159
rect 5997 36119 6055 36125
rect 6181 36159 6239 36165
rect 6181 36125 6193 36159
rect 6227 36156 6239 36159
rect 6549 36159 6607 36165
rect 6549 36156 6561 36159
rect 6227 36128 6561 36156
rect 6227 36125 6239 36128
rect 6181 36119 6239 36125
rect 6549 36125 6561 36128
rect 6595 36156 6607 36159
rect 6730 36156 6736 36168
rect 6595 36128 6736 36156
rect 6595 36125 6607 36128
rect 6549 36119 6607 36125
rect 4571 36060 4660 36088
rect 4816 36088 4844 36119
rect 5092 36088 5120 36119
rect 6730 36116 6736 36128
rect 6788 36116 6794 36168
rect 6840 36165 6868 36196
rect 10689 36193 10701 36196
rect 10735 36224 10747 36227
rect 11054 36224 11060 36236
rect 10735 36196 11060 36224
rect 10735 36193 10747 36196
rect 10689 36187 10747 36193
rect 11054 36184 11060 36196
rect 11112 36184 11118 36236
rect 12069 36227 12127 36233
rect 12069 36193 12081 36227
rect 12115 36224 12127 36227
rect 12894 36224 12900 36236
rect 12115 36196 12900 36224
rect 12115 36193 12127 36196
rect 12069 36187 12127 36193
rect 12894 36184 12900 36196
rect 12952 36184 12958 36236
rect 6825 36159 6883 36165
rect 6825 36125 6837 36159
rect 6871 36156 6883 36159
rect 7006 36156 7012 36168
rect 6871 36128 7012 36156
rect 6871 36125 6883 36128
rect 6825 36119 6883 36125
rect 7006 36116 7012 36128
rect 7064 36116 7070 36168
rect 8662 36116 8668 36168
rect 8720 36116 8726 36168
rect 4816 36060 5120 36088
rect 4571 36057 4583 36060
rect 4525 36051 4583 36057
rect 5534 36048 5540 36100
rect 5592 36088 5598 36100
rect 6365 36091 6423 36097
rect 6365 36088 6377 36091
rect 5592 36060 6377 36088
rect 5592 36048 5598 36060
rect 6365 36057 6377 36060
rect 6411 36057 6423 36091
rect 7958 36060 8156 36088
rect 6365 36051 6423 36057
rect 4709 36023 4767 36029
rect 4709 36020 4721 36023
rect 4172 35992 4721 36020
rect 4709 35989 4721 35992
rect 4755 36020 4767 36023
rect 4798 36020 4804 36032
rect 4755 35992 4804 36020
rect 4755 35989 4767 35992
rect 4709 35983 4767 35989
rect 4798 35980 4804 35992
rect 4856 35980 4862 36032
rect 4985 36023 5043 36029
rect 4985 35989 4997 36023
rect 5031 36020 5043 36023
rect 5350 36020 5356 36032
rect 5031 35992 5356 36020
rect 5031 35989 5043 35992
rect 4985 35983 5043 35989
rect 5350 35980 5356 35992
rect 5408 35980 5414 36032
rect 6733 36023 6791 36029
rect 6733 35989 6745 36023
rect 6779 36020 6791 36023
rect 6822 36020 6828 36032
rect 6779 35992 6828 36020
rect 6779 35989 6791 35992
rect 6733 35983 6791 35989
rect 6822 35980 6828 35992
rect 6880 35980 6886 36032
rect 6914 35980 6920 36032
rect 6972 35980 6978 36032
rect 7098 35980 7104 36032
rect 7156 36020 7162 36032
rect 8128 36020 8156 36060
rect 8386 36048 8392 36100
rect 8444 36048 8450 36100
rect 9232 36094 9352 36122
rect 13446 36116 13452 36168
rect 13504 36122 13510 36168
rect 13504 36116 13768 36122
rect 14090 36116 14096 36168
rect 14148 36116 14154 36168
rect 14458 36116 14464 36168
rect 14516 36156 14522 36168
rect 15013 36159 15071 36165
rect 15013 36156 15025 36159
rect 14516 36128 15025 36156
rect 14516 36116 14522 36128
rect 15013 36125 15025 36128
rect 15059 36125 15071 36159
rect 16500 36156 16528 36252
rect 17589 36227 17647 36233
rect 17589 36193 17601 36227
rect 17635 36224 17647 36227
rect 18046 36224 18052 36236
rect 17635 36196 18052 36224
rect 17635 36193 17647 36196
rect 17589 36187 17647 36193
rect 18046 36184 18052 36196
rect 18104 36184 18110 36236
rect 18708 36196 20300 36224
rect 16853 36159 16911 36165
rect 16853 36156 16865 36159
rect 16500 36128 16865 36156
rect 15013 36119 15071 36125
rect 16853 36125 16865 36128
rect 16899 36125 16911 36159
rect 16853 36119 16911 36125
rect 16942 36116 16948 36168
rect 17000 36156 17006 36168
rect 17000 36128 17045 36156
rect 17000 36116 17006 36128
rect 17126 36116 17132 36168
rect 17184 36156 17190 36168
rect 17313 36159 17371 36165
rect 17313 36156 17325 36159
rect 17184 36128 17325 36156
rect 17184 36116 17190 36128
rect 17313 36125 17325 36128
rect 17359 36125 17371 36159
rect 18708 36142 18736 36196
rect 19245 36159 19303 36165
rect 19245 36156 19257 36159
rect 17313 36119 17371 36125
rect 19076 36128 19257 36156
rect 9232 36088 9260 36094
rect 8496 36074 9260 36088
rect 8496 36060 9246 36074
rect 8496 36020 8524 36060
rect 7156 35992 8524 36020
rect 7156 35980 7162 35992
rect 8938 35980 8944 36032
rect 8996 35980 9002 36032
rect 9324 36020 9352 36094
rect 10318 36088 10324 36100
rect 9982 36060 10324 36088
rect 10060 36020 10088 36060
rect 10318 36048 10324 36060
rect 10376 36048 10382 36100
rect 10410 36048 10416 36100
rect 10468 36048 10474 36100
rect 12345 36091 12403 36097
rect 13464 36094 13768 36116
rect 12345 36057 12357 36091
rect 12391 36057 12403 36091
rect 13740 36088 13768 36094
rect 13740 36060 14872 36088
rect 12345 36051 12403 36057
rect 9324 35992 10088 36020
rect 12360 36020 12388 36051
rect 13722 36020 13728 36032
rect 12360 35992 13728 36020
rect 13722 35980 13728 35992
rect 13780 35980 13786 36032
rect 14182 35980 14188 36032
rect 14240 36020 14246 36032
rect 14737 36023 14795 36029
rect 14737 36020 14749 36023
rect 14240 35992 14749 36020
rect 14240 35980 14246 35992
rect 14737 35989 14749 35992
rect 14783 35989 14795 36023
rect 14844 36020 14872 36060
rect 15286 36048 15292 36100
rect 15344 36048 15350 36100
rect 15746 36088 15752 36100
rect 15396 36060 15752 36088
rect 15396 36020 15424 36060
rect 15746 36048 15752 36060
rect 15804 36048 15810 36100
rect 14844 35992 15424 36020
rect 14737 35983 14795 35989
rect 15930 35980 15936 36032
rect 15988 36020 15994 36032
rect 17221 36023 17279 36029
rect 17221 36020 17233 36023
rect 15988 35992 17233 36020
rect 15988 35980 15994 35992
rect 17221 35989 17233 35992
rect 17267 35989 17279 36023
rect 17221 35983 17279 35989
rect 18506 35980 18512 36032
rect 18564 36020 18570 36032
rect 19076 36029 19104 36128
rect 19245 36125 19257 36128
rect 19291 36125 19303 36159
rect 20272 36156 20300 36196
rect 21174 36184 21180 36236
rect 21232 36224 21238 36236
rect 21634 36224 21640 36236
rect 21232 36196 21640 36224
rect 21232 36184 21238 36196
rect 21634 36184 21640 36196
rect 21692 36184 21698 36236
rect 21913 36227 21971 36233
rect 21913 36193 21925 36227
rect 21959 36224 21971 36227
rect 22646 36224 22652 36236
rect 21959 36196 22652 36224
rect 21959 36193 21971 36196
rect 21913 36187 21971 36193
rect 22646 36184 22652 36196
rect 22704 36224 22710 36236
rect 23014 36224 23020 36236
rect 22704 36196 23020 36224
rect 22704 36184 22710 36196
rect 23014 36184 23020 36196
rect 23072 36184 23078 36236
rect 23382 36184 23388 36236
rect 23440 36184 23446 36236
rect 21450 36156 21456 36168
rect 20272 36128 21456 36156
rect 19245 36119 19303 36125
rect 21450 36116 21456 36128
rect 21508 36116 21514 36168
rect 23661 36159 23719 36165
rect 23661 36125 23673 36159
rect 23707 36125 23719 36159
rect 23661 36119 23719 36125
rect 22954 36060 23428 36088
rect 19061 36023 19119 36029
rect 19061 36020 19073 36023
rect 18564 35992 19073 36020
rect 18564 35980 18570 35992
rect 19061 35989 19073 35992
rect 19107 35989 19119 36023
rect 19061 35983 19119 35989
rect 20898 35980 20904 36032
rect 20956 35980 20962 36032
rect 20993 36023 21051 36029
rect 20993 35989 21005 36023
rect 21039 36020 21051 36023
rect 21358 36020 21364 36032
rect 21039 35992 21364 36020
rect 21039 35989 21051 35992
rect 20993 35983 21051 35989
rect 21358 35980 21364 35992
rect 21416 35980 21422 36032
rect 23400 36020 23428 36060
rect 23474 36048 23480 36100
rect 23532 36088 23538 36100
rect 23676 36088 23704 36119
rect 24394 36116 24400 36168
rect 24452 36156 24458 36168
rect 25041 36159 25099 36165
rect 25041 36156 25053 36159
rect 24452 36128 25053 36156
rect 24452 36116 24458 36128
rect 25041 36125 25053 36128
rect 25087 36125 25099 36159
rect 25041 36119 25099 36125
rect 27062 36116 27068 36168
rect 27120 36156 27126 36168
rect 27249 36159 27307 36165
rect 27249 36156 27261 36159
rect 27120 36128 27261 36156
rect 27120 36116 27126 36128
rect 27249 36125 27261 36128
rect 27295 36125 27307 36159
rect 28736 36156 28764 36332
rect 28920 36332 30472 36360
rect 28920 36224 28948 36332
rect 30466 36320 30472 36332
rect 30524 36320 30530 36372
rect 30650 36320 30656 36372
rect 30708 36360 30714 36372
rect 30745 36363 30803 36369
rect 30745 36360 30757 36363
rect 30708 36332 30757 36360
rect 30708 36320 30714 36332
rect 30745 36329 30757 36332
rect 30791 36329 30803 36363
rect 30745 36323 30803 36329
rect 30929 36363 30987 36369
rect 30929 36329 30941 36363
rect 30975 36329 30987 36363
rect 30929 36323 30987 36329
rect 28997 36295 29055 36301
rect 28997 36261 29009 36295
rect 29043 36292 29055 36295
rect 30098 36292 30104 36304
rect 29043 36264 30104 36292
rect 29043 36261 29055 36264
rect 28997 36255 29055 36261
rect 30098 36252 30104 36264
rect 30156 36252 30162 36304
rect 30944 36292 30972 36323
rect 31110 36320 31116 36372
rect 31168 36360 31174 36372
rect 31481 36363 31539 36369
rect 31481 36360 31493 36363
rect 31168 36332 31493 36360
rect 31168 36320 31174 36332
rect 31481 36329 31493 36332
rect 31527 36329 31539 36363
rect 31481 36323 31539 36329
rect 32217 36363 32275 36369
rect 32217 36329 32229 36363
rect 32263 36360 32275 36363
rect 32398 36360 32404 36372
rect 32263 36332 32404 36360
rect 32263 36329 32275 36332
rect 32217 36323 32275 36329
rect 32398 36320 32404 36332
rect 32456 36320 32462 36372
rect 34146 36360 34152 36372
rect 32876 36332 34152 36360
rect 30668 36264 30972 36292
rect 30668 36233 30696 36264
rect 30653 36227 30711 36233
rect 28920 36196 29224 36224
rect 29086 36156 29092 36168
rect 28736 36128 29092 36156
rect 27249 36119 27307 36125
rect 29086 36116 29092 36128
rect 29144 36116 29150 36168
rect 29196 36165 29224 36196
rect 29380 36196 30328 36224
rect 29380 36165 29408 36196
rect 29181 36159 29239 36165
rect 29181 36125 29193 36159
rect 29227 36125 29239 36159
rect 29181 36119 29239 36125
rect 29365 36159 29423 36165
rect 29365 36125 29377 36159
rect 29411 36125 29423 36159
rect 29365 36119 29423 36125
rect 30098 36116 30104 36168
rect 30156 36116 30162 36168
rect 30300 36165 30328 36196
rect 30653 36193 30665 36227
rect 30699 36193 30711 36227
rect 30944 36224 30972 36264
rect 30944 36196 31340 36224
rect 30653 36187 30711 36193
rect 30285 36159 30343 36165
rect 30285 36125 30297 36159
rect 30331 36156 30343 36159
rect 31018 36156 31024 36168
rect 30331 36128 31024 36156
rect 30331 36125 30343 36128
rect 30285 36119 30343 36125
rect 31018 36116 31024 36128
rect 31076 36116 31082 36168
rect 31202 36116 31208 36168
rect 31260 36116 31266 36168
rect 31312 36165 31340 36196
rect 32490 36184 32496 36236
rect 32548 36224 32554 36236
rect 32876 36233 32904 36332
rect 34146 36320 34152 36332
rect 34204 36320 34210 36372
rect 34425 36363 34483 36369
rect 34425 36329 34437 36363
rect 34471 36360 34483 36363
rect 34790 36360 34796 36372
rect 34471 36332 34796 36360
rect 34471 36329 34483 36332
rect 34425 36323 34483 36329
rect 34790 36320 34796 36332
rect 34848 36320 34854 36372
rect 35161 36363 35219 36369
rect 35161 36329 35173 36363
rect 35207 36360 35219 36363
rect 36446 36360 36452 36372
rect 35207 36332 36452 36360
rect 35207 36329 35219 36332
rect 35161 36323 35219 36329
rect 36446 36320 36452 36332
rect 36504 36360 36510 36372
rect 36633 36363 36691 36369
rect 36633 36360 36645 36363
rect 36504 36332 36645 36360
rect 36504 36320 36510 36332
rect 36633 36329 36645 36332
rect 36679 36329 36691 36363
rect 36633 36323 36691 36329
rect 37182 36320 37188 36372
rect 37240 36320 37246 36372
rect 37918 36360 37924 36372
rect 37292 36332 37924 36360
rect 33962 36292 33968 36304
rect 32968 36264 33968 36292
rect 32677 36227 32735 36233
rect 32677 36224 32689 36227
rect 32548 36196 32689 36224
rect 32548 36184 32554 36196
rect 32677 36193 32689 36196
rect 32723 36193 32735 36227
rect 32677 36187 32735 36193
rect 32861 36227 32919 36233
rect 32861 36193 32873 36227
rect 32907 36193 32919 36227
rect 32861 36187 32919 36193
rect 31297 36159 31355 36165
rect 31297 36125 31309 36159
rect 31343 36125 31355 36159
rect 31297 36119 31355 36125
rect 32585 36159 32643 36165
rect 32585 36125 32597 36159
rect 32631 36156 32643 36159
rect 32968 36156 32996 36264
rect 33962 36252 33968 36264
rect 34020 36252 34026 36304
rect 34333 36295 34391 36301
rect 34333 36261 34345 36295
rect 34379 36292 34391 36295
rect 34882 36292 34888 36304
rect 34379 36264 34888 36292
rect 34379 36261 34391 36264
rect 34333 36255 34391 36261
rect 34882 36252 34888 36264
rect 34940 36292 34946 36304
rect 37292 36292 37320 36332
rect 37918 36320 37924 36332
rect 37976 36320 37982 36372
rect 39022 36320 39028 36372
rect 39080 36320 39086 36372
rect 39942 36320 39948 36372
rect 40000 36320 40006 36372
rect 40218 36320 40224 36372
rect 40276 36360 40282 36372
rect 41230 36360 41236 36372
rect 40276 36332 41236 36360
rect 40276 36320 40282 36332
rect 41230 36320 41236 36332
rect 41288 36320 41294 36372
rect 42150 36320 42156 36372
rect 42208 36320 42214 36372
rect 34940 36264 37320 36292
rect 34940 36252 34946 36264
rect 37458 36252 37464 36304
rect 37516 36252 37522 36304
rect 37553 36295 37611 36301
rect 37553 36261 37565 36295
rect 37599 36292 37611 36295
rect 37642 36292 37648 36304
rect 37599 36264 37648 36292
rect 37599 36261 37611 36264
rect 37553 36255 37611 36261
rect 37642 36252 37648 36264
rect 37700 36252 37706 36304
rect 38930 36292 38936 36304
rect 37844 36264 38936 36292
rect 33060 36196 33548 36224
rect 33060 36165 33088 36196
rect 33520 36165 33548 36196
rect 33778 36184 33784 36236
rect 33836 36224 33842 36236
rect 34773 36227 34831 36233
rect 34773 36224 34785 36227
rect 33836 36196 34785 36224
rect 33836 36184 33842 36196
rect 34773 36193 34785 36196
rect 34819 36193 34831 36227
rect 34773 36187 34831 36193
rect 35345 36227 35403 36233
rect 35345 36193 35357 36227
rect 35391 36224 35403 36227
rect 36170 36224 36176 36236
rect 35391 36196 36176 36224
rect 35391 36193 35403 36196
rect 35345 36187 35403 36193
rect 36170 36184 36176 36196
rect 36228 36184 36234 36236
rect 37001 36227 37059 36233
rect 37001 36193 37013 36227
rect 37047 36224 37059 36227
rect 37476 36224 37504 36252
rect 37047 36196 37504 36224
rect 37047 36193 37059 36196
rect 37001 36187 37059 36193
rect 32631 36128 32996 36156
rect 33045 36159 33103 36165
rect 32631 36125 32643 36128
rect 32585 36119 32643 36125
rect 33045 36125 33057 36159
rect 33091 36125 33103 36159
rect 33045 36119 33103 36125
rect 33229 36159 33287 36165
rect 33229 36125 33241 36159
rect 33275 36125 33287 36159
rect 33229 36119 33287 36125
rect 33505 36159 33563 36165
rect 33505 36125 33517 36159
rect 33551 36125 33563 36159
rect 34977 36159 35035 36165
rect 34977 36156 34989 36159
rect 33505 36119 33563 36125
rect 33612 36128 34989 36156
rect 23532 36060 23704 36088
rect 23532 36048 23538 36060
rect 25314 36048 25320 36100
rect 25372 36048 25378 36100
rect 25774 36088 25780 36100
rect 25424 36060 25780 36088
rect 23934 36020 23940 36032
rect 23400 35992 23940 36020
rect 23934 35980 23940 35992
rect 23992 36020 23998 36032
rect 25130 36020 25136 36032
rect 23992 35992 25136 36020
rect 23992 35980 23998 35992
rect 25130 35980 25136 35992
rect 25188 36020 25194 36032
rect 25424 36020 25452 36060
rect 25774 36048 25780 36060
rect 25832 36048 25838 36100
rect 27525 36091 27583 36097
rect 27525 36057 27537 36091
rect 27571 36088 27583 36091
rect 27798 36088 27804 36100
rect 27571 36060 27804 36088
rect 27571 36057 27583 36060
rect 27525 36051 27583 36057
rect 27798 36048 27804 36060
rect 27856 36048 27862 36100
rect 28902 36088 28908 36100
rect 28750 36060 28908 36088
rect 28902 36048 28908 36060
rect 28960 36048 28966 36100
rect 29273 36091 29331 36097
rect 29273 36057 29285 36091
rect 29319 36088 29331 36091
rect 29319 36060 30420 36088
rect 29319 36057 29331 36060
rect 29273 36051 29331 36057
rect 25188 35992 25452 36020
rect 26789 36023 26847 36029
rect 25188 35980 25194 35992
rect 26789 35989 26801 36023
rect 26835 36020 26847 36023
rect 27338 36020 27344 36032
rect 26835 35992 27344 36020
rect 26835 35989 26847 35992
rect 26789 35983 26847 35989
rect 27338 35980 27344 35992
rect 27396 35980 27402 36032
rect 29546 35980 29552 36032
rect 29604 35980 29610 36032
rect 30392 36020 30420 36060
rect 30466 36048 30472 36100
rect 30524 36048 30530 36100
rect 31113 36091 31171 36097
rect 31113 36057 31125 36091
rect 31159 36088 31171 36091
rect 31478 36088 31484 36100
rect 31159 36060 31484 36088
rect 31159 36057 31171 36060
rect 31113 36051 31171 36057
rect 31478 36048 31484 36060
rect 31536 36048 31542 36100
rect 31662 36048 31668 36100
rect 31720 36088 31726 36100
rect 33060 36088 33088 36119
rect 31720 36060 33088 36088
rect 33244 36088 33272 36119
rect 33321 36091 33379 36097
rect 33321 36088 33333 36091
rect 33244 36060 33333 36088
rect 31720 36048 31726 36060
rect 33321 36057 33333 36060
rect 33367 36088 33379 36091
rect 33410 36088 33416 36100
rect 33367 36060 33416 36088
rect 33367 36057 33379 36060
rect 33321 36051 33379 36057
rect 33410 36048 33416 36060
rect 33468 36048 33474 36100
rect 30903 36023 30961 36029
rect 30903 36020 30915 36023
rect 30392 35992 30915 36020
rect 30903 35989 30915 35992
rect 30949 36020 30961 36023
rect 31202 36020 31208 36032
rect 30949 35992 31208 36020
rect 30949 35989 30961 35992
rect 30903 35983 30961 35989
rect 31202 35980 31208 35992
rect 31260 35980 31266 36032
rect 33137 36023 33195 36029
rect 33137 35989 33149 36023
rect 33183 36020 33195 36023
rect 33612 36020 33640 36128
rect 34808 36100 34836 36128
rect 34977 36125 34989 36128
rect 35023 36125 35035 36159
rect 34977 36119 35035 36125
rect 35069 36159 35127 36165
rect 35069 36125 35081 36159
rect 35115 36156 35127 36159
rect 35250 36156 35256 36168
rect 35115 36128 35256 36156
rect 35115 36125 35127 36128
rect 35069 36119 35127 36125
rect 35250 36116 35256 36128
rect 35308 36116 35314 36168
rect 36909 36159 36967 36165
rect 36909 36125 36921 36159
rect 36955 36156 36967 36159
rect 37274 36156 37280 36168
rect 36955 36128 37280 36156
rect 36955 36125 36967 36128
rect 36909 36119 36967 36125
rect 37274 36116 37280 36128
rect 37332 36116 37338 36168
rect 37366 36116 37372 36168
rect 37424 36116 37430 36168
rect 37461 36159 37519 36165
rect 37461 36125 37473 36159
rect 37507 36156 37519 36159
rect 37550 36156 37556 36168
rect 37507 36128 37556 36156
rect 37507 36125 37519 36128
rect 37461 36119 37519 36125
rect 37550 36116 37556 36128
rect 37608 36116 37614 36168
rect 37844 36165 37872 36264
rect 38930 36252 38936 36264
rect 38988 36252 38994 36304
rect 39574 36252 39580 36304
rect 39632 36292 39638 36304
rect 39669 36295 39727 36301
rect 39669 36292 39681 36295
rect 39632 36264 39681 36292
rect 39632 36252 39638 36264
rect 39669 36261 39681 36264
rect 39715 36292 39727 36295
rect 40034 36292 40040 36304
rect 39715 36264 40040 36292
rect 39715 36261 39727 36264
rect 39669 36255 39727 36261
rect 40034 36252 40040 36264
rect 40092 36252 40098 36304
rect 38580 36196 39344 36224
rect 37645 36159 37703 36165
rect 37645 36125 37657 36159
rect 37691 36125 37703 36159
rect 37645 36119 37703 36125
rect 37829 36159 37887 36165
rect 37829 36125 37841 36159
rect 37875 36125 37887 36159
rect 37829 36119 37887 36125
rect 33778 36048 33784 36100
rect 33836 36088 33842 36100
rect 33965 36091 34023 36097
rect 33965 36088 33977 36091
rect 33836 36060 33977 36088
rect 33836 36048 33842 36060
rect 33965 36057 33977 36060
rect 34011 36057 34023 36091
rect 33965 36051 34023 36057
rect 34606 36048 34612 36100
rect 34664 36088 34670 36100
rect 34701 36091 34759 36097
rect 34701 36088 34713 36091
rect 34664 36060 34713 36088
rect 34664 36048 34670 36060
rect 34701 36057 34713 36060
rect 34747 36057 34759 36091
rect 34701 36051 34759 36057
rect 34790 36048 34796 36100
rect 34848 36048 34854 36100
rect 33183 35992 33640 36020
rect 33689 36023 33747 36029
rect 33183 35989 33195 35992
rect 33137 35983 33195 35989
rect 33689 35989 33701 36023
rect 33735 36020 33747 36023
rect 34514 36020 34520 36032
rect 33735 35992 34520 36020
rect 33735 35989 33747 35992
rect 33689 35983 33747 35989
rect 34514 35980 34520 35992
rect 34572 36020 34578 36032
rect 34885 36023 34943 36029
rect 34885 36020 34897 36023
rect 34572 35992 34897 36020
rect 34572 35980 34578 35992
rect 34885 35989 34897 35992
rect 34931 35989 34943 36023
rect 34885 35983 34943 35989
rect 35345 36023 35403 36029
rect 35345 35989 35357 36023
rect 35391 36020 35403 36023
rect 36078 36020 36084 36032
rect 35391 35992 36084 36020
rect 35391 35989 35403 35992
rect 35345 35983 35403 35989
rect 36078 35980 36084 35992
rect 36136 35980 36142 36032
rect 37384 36020 37412 36116
rect 37660 36088 37688 36119
rect 38010 36116 38016 36168
rect 38068 36116 38074 36168
rect 38105 36159 38163 36165
rect 38105 36125 38117 36159
rect 38151 36156 38163 36159
rect 38580 36156 38608 36196
rect 39316 36168 39344 36196
rect 40678 36184 40684 36236
rect 40736 36184 40742 36236
rect 38151 36128 38608 36156
rect 38151 36125 38163 36128
rect 38105 36119 38163 36125
rect 38654 36116 38660 36168
rect 38712 36116 38718 36168
rect 38930 36116 38936 36168
rect 38988 36156 38994 36168
rect 39025 36159 39083 36165
rect 39025 36156 39037 36159
rect 38988 36128 39037 36156
rect 38988 36116 38994 36128
rect 39025 36125 39037 36128
rect 39071 36125 39083 36159
rect 39025 36119 39083 36125
rect 39298 36116 39304 36168
rect 39356 36116 39362 36168
rect 39574 36116 39580 36168
rect 39632 36156 39638 36168
rect 40405 36159 40463 36165
rect 40405 36156 40417 36159
rect 39632 36128 40417 36156
rect 39632 36116 39638 36128
rect 40405 36125 40417 36128
rect 40451 36125 40463 36159
rect 40405 36119 40463 36125
rect 38028 36088 38056 36116
rect 37660 36060 38056 36088
rect 38381 36091 38439 36097
rect 38381 36057 38393 36091
rect 38427 36088 38439 36091
rect 38470 36088 38476 36100
rect 38427 36060 38476 36088
rect 38427 36057 38439 36060
rect 38381 36051 38439 36057
rect 38470 36048 38476 36060
rect 38528 36048 38534 36100
rect 38562 36048 38568 36100
rect 38620 36048 38626 36100
rect 39117 36091 39175 36097
rect 39117 36088 39129 36091
rect 38672 36060 39129 36088
rect 37927 36023 37985 36029
rect 37927 36020 37939 36023
rect 37384 35992 37939 36020
rect 37927 35989 37939 35992
rect 37973 35989 37985 36023
rect 37927 35983 37985 35989
rect 38013 36023 38071 36029
rect 38013 35989 38025 36023
rect 38059 36020 38071 36023
rect 38197 36023 38255 36029
rect 38197 36020 38209 36023
rect 38059 35992 38209 36020
rect 38059 35989 38071 35992
rect 38013 35983 38071 35989
rect 38197 35989 38209 35992
rect 38243 36020 38255 36023
rect 38672 36020 38700 36060
rect 39117 36057 39129 36060
rect 39163 36057 39175 36091
rect 39117 36051 39175 36057
rect 39206 36048 39212 36100
rect 39264 36088 39270 36100
rect 39485 36091 39543 36097
rect 39485 36088 39497 36091
rect 39264 36060 39497 36088
rect 39264 36048 39270 36060
rect 39485 36057 39497 36060
rect 39531 36057 39543 36091
rect 39485 36051 39543 36057
rect 40034 36048 40040 36100
rect 40092 36088 40098 36100
rect 40129 36091 40187 36097
rect 40129 36088 40141 36091
rect 40092 36060 40141 36088
rect 40092 36048 40098 36060
rect 40129 36057 40141 36060
rect 40175 36057 40187 36091
rect 40129 36051 40187 36057
rect 40310 36048 40316 36100
rect 40368 36048 40374 36100
rect 41414 36048 41420 36100
rect 41472 36048 41478 36100
rect 38243 35992 38700 36020
rect 38243 35989 38255 35992
rect 38197 35983 38255 35989
rect 38746 35980 38752 36032
rect 38804 36020 38810 36032
rect 38841 36023 38899 36029
rect 38841 36020 38853 36023
rect 38804 35992 38853 36020
rect 38804 35980 38810 35992
rect 38841 35989 38853 35992
rect 38887 36020 38899 36023
rect 40218 36020 40224 36032
rect 38887 35992 40224 36020
rect 38887 35989 38899 35992
rect 38841 35983 38899 35989
rect 40218 35980 40224 35992
rect 40276 35980 40282 36032
rect 1104 35930 42504 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 42504 35930
rect 1104 35856 42504 35878
rect 3878 35776 3884 35828
rect 3936 35816 3942 35828
rect 3936 35788 5488 35816
rect 3936 35776 3942 35788
rect 3234 35748 3240 35760
rect 2700 35720 3240 35748
rect 2700 35689 2728 35720
rect 3234 35708 3240 35720
rect 3292 35708 3298 35760
rect 4614 35748 4620 35760
rect 4186 35720 4620 35748
rect 4614 35708 4620 35720
rect 4672 35708 4678 35760
rect 4798 35708 4804 35760
rect 4856 35748 4862 35760
rect 4856 35720 4936 35748
rect 4856 35708 4862 35720
rect 2685 35683 2743 35689
rect 2685 35649 2697 35683
rect 2731 35649 2743 35683
rect 2685 35643 2743 35649
rect 4706 35640 4712 35692
rect 4764 35640 4770 35692
rect 4908 35689 4936 35720
rect 4893 35683 4951 35689
rect 4893 35649 4905 35683
rect 4939 35649 4951 35683
rect 4893 35643 4951 35649
rect 4982 35640 4988 35692
rect 5040 35640 5046 35692
rect 5350 35640 5356 35692
rect 5408 35640 5414 35692
rect 5460 35680 5488 35788
rect 8386 35776 8392 35828
rect 8444 35776 8450 35828
rect 9953 35819 10011 35825
rect 9953 35785 9965 35819
rect 9999 35816 10011 35819
rect 10410 35816 10416 35828
rect 9999 35788 10416 35816
rect 9999 35785 10011 35788
rect 9953 35779 10011 35785
rect 10410 35776 10416 35788
rect 10468 35776 10474 35828
rect 13311 35819 13369 35825
rect 13311 35785 13323 35819
rect 13357 35816 13369 35819
rect 14090 35816 14096 35828
rect 13357 35788 14096 35816
rect 13357 35785 13369 35788
rect 13311 35779 13369 35785
rect 14090 35776 14096 35788
rect 14148 35776 14154 35828
rect 14458 35776 14464 35828
rect 14516 35816 14522 35828
rect 16209 35819 16267 35825
rect 14516 35788 16160 35816
rect 14516 35776 14522 35788
rect 5534 35708 5540 35760
rect 5592 35708 5598 35760
rect 5629 35751 5687 35757
rect 5629 35717 5641 35751
rect 5675 35748 5687 35751
rect 6365 35751 6423 35757
rect 6365 35748 6377 35751
rect 5675 35720 6377 35748
rect 5675 35717 5687 35720
rect 5629 35711 5687 35717
rect 6365 35717 6377 35720
rect 6411 35717 6423 35751
rect 6365 35711 6423 35717
rect 6822 35708 6828 35760
rect 6880 35748 6886 35760
rect 8754 35748 8760 35760
rect 6880 35720 8760 35748
rect 6880 35708 6886 35720
rect 8754 35708 8760 35720
rect 8812 35708 8818 35760
rect 8895 35751 8953 35757
rect 8895 35717 8907 35751
rect 8941 35748 8953 35751
rect 9861 35751 9919 35757
rect 8941 35720 9628 35748
rect 8941 35717 8953 35720
rect 8895 35711 8953 35717
rect 5721 35683 5779 35689
rect 5721 35680 5733 35683
rect 5460 35652 5733 35680
rect 5721 35649 5733 35652
rect 5767 35649 5779 35683
rect 6840 35680 6868 35708
rect 5721 35643 5779 35649
rect 5828 35652 6868 35680
rect 2958 35572 2964 35624
rect 3016 35572 3022 35624
rect 4614 35572 4620 35624
rect 4672 35612 4678 35624
rect 4801 35615 4859 35621
rect 4801 35612 4813 35615
rect 4672 35584 4813 35612
rect 4672 35572 4678 35584
rect 4801 35581 4813 35584
rect 4847 35612 4859 35615
rect 5828 35612 5856 35652
rect 7282 35640 7288 35692
rect 7340 35640 7346 35692
rect 7374 35640 7380 35692
rect 7432 35680 7438 35692
rect 8573 35683 8631 35689
rect 8573 35680 8585 35683
rect 7432 35652 8585 35680
rect 7432 35640 7438 35652
rect 8573 35649 8585 35652
rect 8619 35649 8631 35683
rect 8573 35643 8631 35649
rect 8665 35683 8723 35689
rect 8665 35649 8677 35683
rect 8711 35680 8723 35683
rect 8711 35652 8892 35680
rect 8711 35649 8723 35652
rect 8665 35643 8723 35649
rect 4847 35584 5856 35612
rect 4847 35581 4859 35584
rect 4801 35575 4859 35581
rect 5368 35556 5396 35584
rect 6822 35572 6828 35624
rect 6880 35612 6886 35624
rect 6917 35615 6975 35621
rect 6917 35612 6929 35615
rect 6880 35584 6929 35612
rect 6880 35572 6886 35584
rect 6917 35581 6929 35584
rect 6963 35581 6975 35615
rect 6917 35575 6975 35581
rect 4525 35547 4583 35553
rect 4525 35544 4537 35547
rect 3988 35516 4537 35544
rect 3326 35436 3332 35488
rect 3384 35476 3390 35488
rect 3988 35476 4016 35516
rect 4525 35513 4537 35516
rect 4571 35513 4583 35547
rect 4525 35507 4583 35513
rect 5350 35504 5356 35556
rect 5408 35504 5414 35556
rect 5442 35504 5448 35556
rect 5500 35544 5506 35556
rect 7098 35544 7104 35556
rect 5500 35516 7104 35544
rect 5500 35504 5506 35516
rect 7098 35504 7104 35516
rect 7156 35504 7162 35556
rect 8864 35544 8892 35652
rect 9030 35640 9036 35692
rect 9088 35640 9094 35692
rect 9600 35680 9628 35720
rect 9861 35717 9873 35751
rect 9907 35748 9919 35751
rect 10229 35751 10287 35757
rect 10229 35748 10241 35751
rect 9907 35720 10241 35748
rect 9907 35717 9919 35720
rect 9861 35711 9919 35717
rect 10229 35717 10241 35720
rect 10275 35717 10287 35751
rect 10229 35711 10287 35717
rect 10796 35720 11008 35748
rect 10796 35692 10824 35720
rect 9950 35680 9956 35692
rect 9600 35652 9956 35680
rect 9950 35640 9956 35652
rect 10008 35680 10014 35692
rect 10137 35683 10195 35689
rect 10137 35680 10149 35683
rect 10008 35652 10149 35680
rect 10008 35640 10014 35652
rect 10137 35649 10149 35652
rect 10183 35649 10195 35683
rect 10137 35643 10195 35649
rect 10321 35683 10379 35689
rect 10321 35649 10333 35683
rect 10367 35680 10379 35683
rect 10410 35680 10416 35692
rect 10367 35652 10416 35680
rect 10367 35649 10379 35652
rect 10321 35643 10379 35649
rect 10410 35640 10416 35652
rect 10468 35640 10474 35692
rect 10502 35640 10508 35692
rect 10560 35640 10566 35692
rect 10597 35683 10655 35689
rect 10597 35649 10609 35683
rect 10643 35649 10655 35683
rect 10597 35643 10655 35649
rect 8938 35572 8944 35624
rect 8996 35612 9002 35624
rect 9309 35615 9367 35621
rect 9309 35612 9321 35615
rect 8996 35584 9321 35612
rect 8996 35572 9002 35584
rect 9309 35581 9321 35584
rect 9355 35612 9367 35615
rect 10612 35612 10640 35643
rect 10778 35640 10784 35692
rect 10836 35640 10842 35692
rect 10870 35640 10876 35692
rect 10928 35640 10934 35692
rect 10980 35689 11008 35720
rect 11054 35708 11060 35760
rect 11112 35748 11118 35760
rect 13446 35748 13452 35760
rect 11112 35720 11560 35748
rect 12926 35720 13452 35748
rect 11112 35708 11118 35720
rect 11532 35689 11560 35720
rect 13446 35708 13452 35720
rect 13504 35708 13510 35760
rect 13722 35708 13728 35760
rect 13780 35748 13786 35760
rect 14001 35751 14059 35757
rect 14001 35748 14013 35751
rect 13780 35720 14013 35748
rect 13780 35708 13786 35720
rect 14001 35717 14013 35720
rect 14047 35717 14059 35751
rect 14001 35711 14059 35717
rect 14737 35751 14795 35757
rect 14737 35717 14749 35751
rect 14783 35748 14795 35751
rect 15010 35748 15016 35760
rect 14783 35720 15016 35748
rect 14783 35717 14795 35720
rect 14737 35711 14795 35717
rect 15010 35708 15016 35720
rect 15068 35708 15074 35760
rect 15746 35708 15752 35760
rect 15804 35708 15810 35760
rect 16132 35748 16160 35788
rect 16209 35785 16221 35819
rect 16255 35816 16267 35819
rect 17034 35816 17040 35828
rect 16255 35788 17040 35816
rect 16255 35785 16267 35788
rect 16209 35779 16267 35785
rect 17034 35776 17040 35788
rect 17092 35776 17098 35828
rect 17221 35819 17279 35825
rect 17221 35785 17233 35819
rect 17267 35816 17279 35819
rect 18785 35819 18843 35825
rect 18785 35816 18797 35819
rect 17267 35788 18797 35816
rect 17267 35785 17279 35788
rect 17221 35779 17279 35785
rect 18785 35785 18797 35788
rect 18831 35785 18843 35819
rect 18785 35779 18843 35785
rect 22738 35776 22744 35828
rect 22796 35816 22802 35828
rect 22833 35819 22891 35825
rect 22833 35816 22845 35819
rect 22796 35788 22845 35816
rect 22796 35776 22802 35788
rect 22833 35785 22845 35788
rect 22879 35785 22891 35819
rect 22833 35779 22891 35785
rect 22922 35776 22928 35828
rect 22980 35776 22986 35828
rect 23385 35819 23443 35825
rect 23385 35785 23397 35819
rect 23431 35816 23443 35819
rect 26234 35816 26240 35828
rect 23431 35788 26240 35816
rect 23431 35785 23443 35788
rect 23385 35779 23443 35785
rect 17126 35748 17132 35760
rect 16132 35720 17132 35748
rect 17126 35708 17132 35720
rect 17184 35748 17190 35760
rect 18509 35751 18567 35757
rect 18509 35748 18521 35751
rect 17184 35720 18521 35748
rect 17184 35708 17190 35720
rect 18509 35717 18521 35720
rect 18555 35748 18567 35751
rect 18598 35748 18604 35760
rect 18555 35720 18604 35748
rect 18555 35717 18567 35720
rect 18509 35711 18567 35717
rect 18598 35708 18604 35720
rect 18656 35708 18662 35760
rect 20901 35751 20959 35757
rect 20901 35717 20913 35751
rect 20947 35748 20959 35751
rect 21174 35748 21180 35760
rect 20947 35720 21180 35748
rect 20947 35717 20959 35720
rect 20901 35711 20959 35717
rect 21174 35708 21180 35720
rect 21232 35708 21238 35760
rect 22465 35751 22523 35757
rect 22465 35717 22477 35751
rect 22511 35748 22523 35751
rect 22554 35748 22560 35760
rect 22511 35720 22560 35748
rect 22511 35717 22523 35720
rect 22465 35711 22523 35717
rect 22554 35708 22560 35720
rect 22612 35748 22618 35760
rect 23400 35748 23428 35779
rect 26234 35776 26240 35788
rect 26292 35776 26298 35828
rect 27798 35776 27804 35828
rect 27856 35816 27862 35828
rect 27985 35819 28043 35825
rect 27985 35816 27997 35819
rect 27856 35788 27997 35816
rect 27856 35776 27862 35788
rect 27985 35785 27997 35788
rect 28031 35785 28043 35819
rect 27985 35779 28043 35785
rect 28442 35776 28448 35828
rect 28500 35776 28506 35828
rect 30466 35776 30472 35828
rect 30524 35816 30530 35828
rect 31662 35816 31668 35828
rect 30524 35788 31668 35816
rect 30524 35776 30530 35788
rect 31662 35776 31668 35788
rect 31720 35776 31726 35828
rect 34609 35819 34667 35825
rect 34609 35785 34621 35819
rect 34655 35816 34667 35819
rect 34882 35816 34888 35828
rect 34655 35788 34888 35816
rect 34655 35785 34667 35788
rect 34609 35779 34667 35785
rect 34882 35776 34888 35788
rect 34940 35776 34946 35828
rect 35434 35776 35440 35828
rect 35492 35816 35498 35828
rect 35492 35788 35756 35816
rect 35492 35776 35498 35788
rect 22612 35720 23428 35748
rect 22612 35708 22618 35720
rect 23474 35708 23480 35760
rect 23532 35748 23538 35760
rect 23532 35720 24440 35748
rect 23532 35708 23538 35720
rect 10965 35683 11023 35689
rect 10965 35649 10977 35683
rect 11011 35649 11023 35683
rect 10965 35643 11023 35649
rect 11149 35683 11207 35689
rect 11149 35649 11161 35683
rect 11195 35649 11207 35683
rect 11149 35643 11207 35649
rect 11517 35683 11575 35689
rect 11517 35649 11529 35683
rect 11563 35649 11575 35683
rect 11517 35643 11575 35649
rect 9355 35584 10640 35612
rect 10888 35612 10916 35640
rect 11164 35612 11192 35643
rect 13354 35640 13360 35692
rect 13412 35680 13418 35692
rect 13633 35683 13691 35689
rect 13633 35680 13645 35683
rect 13412 35652 13645 35680
rect 13412 35640 13418 35652
rect 13633 35649 13645 35652
rect 13679 35649 13691 35683
rect 13633 35643 13691 35649
rect 13817 35683 13875 35689
rect 13817 35649 13829 35683
rect 13863 35649 13875 35683
rect 13817 35643 13875 35649
rect 13909 35683 13967 35689
rect 13909 35649 13921 35683
rect 13955 35680 13967 35683
rect 14090 35680 14096 35692
rect 13955 35652 14096 35680
rect 13955 35649 13967 35652
rect 13909 35643 13967 35649
rect 10888 35584 11192 35612
rect 11885 35615 11943 35621
rect 9355 35581 9367 35584
rect 9309 35575 9367 35581
rect 11885 35581 11897 35615
rect 11931 35612 11943 35615
rect 12250 35612 12256 35624
rect 11931 35584 12256 35612
rect 11931 35581 11943 35584
rect 11885 35575 11943 35581
rect 12250 35572 12256 35584
rect 12308 35572 12314 35624
rect 12434 35572 12440 35624
rect 12492 35612 12498 35624
rect 13832 35612 13860 35643
rect 14090 35640 14096 35652
rect 14148 35640 14154 35692
rect 14182 35640 14188 35692
rect 14240 35640 14246 35692
rect 14458 35640 14464 35692
rect 14516 35640 14522 35692
rect 17313 35683 17371 35689
rect 17313 35649 17325 35683
rect 17359 35680 17371 35683
rect 17586 35680 17592 35692
rect 17359 35652 17592 35680
rect 17359 35649 17371 35652
rect 17313 35643 17371 35649
rect 17586 35640 17592 35652
rect 17644 35640 17650 35692
rect 17773 35683 17831 35689
rect 17773 35649 17785 35683
rect 17819 35680 17831 35683
rect 19978 35680 19984 35692
rect 17819 35652 19984 35680
rect 17819 35649 17831 35652
rect 17773 35643 17831 35649
rect 14369 35615 14427 35621
rect 14369 35612 14381 35615
rect 12492 35584 14381 35612
rect 12492 35572 12498 35584
rect 14369 35581 14381 35584
rect 14415 35581 14427 35615
rect 14369 35575 14427 35581
rect 15102 35572 15108 35624
rect 15160 35612 15166 35624
rect 15160 35584 16620 35612
rect 15160 35572 15166 35584
rect 11057 35547 11115 35553
rect 11057 35544 11069 35547
rect 8864 35516 11069 35544
rect 11057 35513 11069 35516
rect 11103 35513 11115 35547
rect 11057 35507 11115 35513
rect 13354 35504 13360 35556
rect 13412 35544 13418 35556
rect 16592 35544 16620 35584
rect 17034 35572 17040 35624
rect 17092 35572 17098 35624
rect 16850 35544 16856 35556
rect 13412 35516 14596 35544
rect 16592 35516 16856 35544
rect 13412 35504 13418 35516
rect 3384 35448 4016 35476
rect 4433 35479 4491 35485
rect 3384 35436 3390 35448
rect 4433 35445 4445 35479
rect 4479 35476 4491 35479
rect 4982 35476 4988 35488
rect 4479 35448 4988 35476
rect 4479 35445 4491 35448
rect 4433 35439 4491 35445
rect 4982 35436 4988 35448
rect 5040 35436 5046 35488
rect 5534 35436 5540 35488
rect 5592 35476 5598 35488
rect 5905 35479 5963 35485
rect 5905 35476 5917 35479
rect 5592 35448 5917 35476
rect 5592 35436 5598 35448
rect 5905 35445 5917 35448
rect 5951 35445 5963 35479
rect 5905 35439 5963 35445
rect 8754 35436 8760 35488
rect 8812 35476 8818 35488
rect 10226 35476 10232 35488
rect 8812 35448 10232 35476
rect 8812 35436 8818 35448
rect 10226 35436 10232 35448
rect 10284 35476 10290 35488
rect 10410 35476 10416 35488
rect 10284 35448 10416 35476
rect 10284 35436 10290 35448
rect 10410 35436 10416 35448
rect 10468 35436 10474 35488
rect 10594 35436 10600 35488
rect 10652 35436 10658 35488
rect 12618 35436 12624 35488
rect 12676 35476 12682 35488
rect 13449 35479 13507 35485
rect 13449 35476 13461 35479
rect 12676 35448 13461 35476
rect 12676 35436 12682 35448
rect 13449 35445 13461 35448
rect 13495 35445 13507 35479
rect 14568 35476 14596 35516
rect 16850 35504 16856 35516
rect 16908 35544 16914 35556
rect 18064 35544 18092 35652
rect 19978 35640 19984 35652
rect 20036 35640 20042 35692
rect 21542 35640 21548 35692
rect 21600 35640 21606 35692
rect 24412 35689 24440 35720
rect 25130 35708 25136 35760
rect 25188 35708 25194 35760
rect 28353 35751 28411 35757
rect 28353 35717 28365 35751
rect 28399 35748 28411 35751
rect 29546 35748 29552 35760
rect 28399 35720 29552 35748
rect 28399 35717 28411 35720
rect 28353 35711 28411 35717
rect 29546 35708 29552 35720
rect 29604 35708 29610 35760
rect 30193 35751 30251 35757
rect 30193 35717 30205 35751
rect 30239 35748 30251 35751
rect 30837 35751 30895 35757
rect 30837 35748 30849 35751
rect 30239 35720 30849 35748
rect 30239 35717 30251 35720
rect 30193 35711 30251 35717
rect 30837 35717 30849 35720
rect 30883 35717 30895 35751
rect 30837 35711 30895 35717
rect 31754 35708 31760 35760
rect 31812 35708 31818 35760
rect 34514 35708 34520 35760
rect 34572 35708 34578 35760
rect 34701 35751 34759 35757
rect 34701 35717 34713 35751
rect 34747 35748 34759 35751
rect 34790 35748 34796 35760
rect 34747 35720 34796 35748
rect 34747 35717 34759 35720
rect 34701 35711 34759 35717
rect 34790 35708 34796 35720
rect 34848 35708 34854 35760
rect 35529 35751 35587 35757
rect 35529 35748 35541 35751
rect 35084 35720 35541 35748
rect 35084 35689 35112 35720
rect 35529 35717 35541 35720
rect 35575 35717 35587 35751
rect 35529 35711 35587 35717
rect 35728 35748 35756 35788
rect 39298 35776 39304 35828
rect 39356 35776 39362 35828
rect 40236 35788 41184 35816
rect 35728 35720 36400 35748
rect 23293 35683 23351 35689
rect 23293 35649 23305 35683
rect 23339 35649 23351 35683
rect 23293 35643 23351 35649
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35649 24455 35683
rect 24397 35643 24455 35649
rect 33229 35683 33287 35689
rect 33229 35649 33241 35683
rect 33275 35680 33287 35683
rect 33689 35683 33747 35689
rect 33689 35680 33701 35683
rect 33275 35652 33701 35680
rect 33275 35649 33287 35652
rect 33229 35643 33287 35649
rect 33689 35649 33701 35652
rect 33735 35649 33747 35683
rect 33689 35643 33747 35649
rect 34425 35683 34483 35689
rect 34425 35649 34437 35683
rect 34471 35680 34483 35683
rect 35069 35683 35127 35689
rect 34471 35652 34505 35680
rect 34471 35649 34483 35652
rect 34425 35643 34483 35649
rect 35069 35649 35081 35683
rect 35115 35649 35127 35683
rect 35069 35643 35127 35649
rect 18230 35572 18236 35624
rect 18288 35612 18294 35624
rect 19337 35615 19395 35621
rect 19337 35612 19349 35615
rect 18288 35584 19349 35612
rect 18288 35572 18294 35584
rect 19337 35581 19349 35584
rect 19383 35581 19395 35615
rect 19337 35575 19395 35581
rect 19889 35615 19947 35621
rect 19889 35581 19901 35615
rect 19935 35581 19947 35615
rect 19889 35575 19947 35581
rect 20441 35615 20499 35621
rect 20441 35581 20453 35615
rect 20487 35612 20499 35615
rect 20993 35615 21051 35621
rect 20993 35612 21005 35615
rect 20487 35584 21005 35612
rect 20487 35581 20499 35584
rect 20441 35575 20499 35581
rect 20993 35581 21005 35584
rect 21039 35581 21051 35615
rect 20993 35575 21051 35581
rect 21177 35615 21235 35621
rect 21177 35581 21189 35615
rect 21223 35612 21235 35615
rect 21223 35584 21496 35612
rect 21223 35581 21235 35584
rect 21177 35575 21235 35581
rect 16908 35516 18092 35544
rect 19904 35544 19932 35575
rect 20898 35544 20904 35556
rect 19904 35516 20904 35544
rect 16908 35504 16914 35516
rect 20898 35504 20904 35516
rect 20956 35504 20962 35556
rect 17310 35476 17316 35488
rect 14568 35448 17316 35476
rect 13449 35439 13507 35445
rect 17310 35436 17316 35448
rect 17368 35436 17374 35488
rect 17678 35436 17684 35488
rect 17736 35436 17742 35488
rect 20530 35436 20536 35488
rect 20588 35436 20594 35488
rect 21468 35485 21496 35584
rect 21634 35572 21640 35624
rect 21692 35612 21698 35624
rect 22281 35615 22339 35621
rect 22281 35612 22293 35615
rect 21692 35584 22293 35612
rect 21692 35572 21698 35584
rect 22281 35581 22293 35584
rect 22327 35581 22339 35615
rect 22281 35575 22339 35581
rect 22296 35544 22324 35575
rect 22370 35572 22376 35624
rect 22428 35612 22434 35624
rect 23308 35612 23336 35643
rect 22428 35584 23336 35612
rect 23569 35615 23627 35621
rect 22428 35572 22434 35584
rect 23569 35581 23581 35615
rect 23615 35581 23627 35615
rect 23569 35575 23627 35581
rect 23584 35544 23612 35575
rect 24670 35572 24676 35624
rect 24728 35572 24734 35624
rect 25406 35572 25412 35624
rect 25464 35612 25470 35624
rect 26145 35615 26203 35621
rect 26145 35612 26157 35615
rect 25464 35584 26157 35612
rect 25464 35572 25470 35584
rect 26145 35581 26157 35584
rect 26191 35612 26203 35615
rect 27525 35615 27583 35621
rect 27525 35612 27537 35615
rect 26191 35584 27537 35612
rect 26191 35581 26203 35584
rect 26145 35575 26203 35581
rect 27525 35581 27537 35584
rect 27571 35581 27583 35615
rect 27525 35575 27583 35581
rect 28629 35615 28687 35621
rect 28629 35581 28641 35615
rect 28675 35612 28687 35615
rect 28902 35612 28908 35624
rect 28675 35584 28908 35612
rect 28675 35581 28687 35584
rect 28629 35575 28687 35581
rect 28902 35572 28908 35584
rect 28960 35572 28966 35624
rect 30285 35615 30343 35621
rect 30285 35612 30297 35615
rect 30208 35584 30297 35612
rect 30208 35556 30236 35584
rect 30285 35581 30297 35584
rect 30331 35581 30343 35615
rect 30285 35575 30343 35581
rect 30469 35615 30527 35621
rect 30469 35581 30481 35615
rect 30515 35581 30527 35615
rect 30469 35575 30527 35581
rect 22296 35516 23612 35544
rect 21453 35479 21511 35485
rect 21453 35445 21465 35479
rect 21499 35476 21511 35479
rect 22094 35476 22100 35488
rect 21499 35448 22100 35476
rect 21499 35445 21511 35448
rect 21453 35439 21511 35445
rect 22094 35436 22100 35448
rect 22152 35436 22158 35488
rect 23584 35476 23612 35516
rect 30190 35504 30196 35556
rect 30248 35504 30254 35556
rect 30484 35544 30512 35575
rect 31018 35572 31024 35624
rect 31076 35612 31082 35624
rect 31389 35615 31447 35621
rect 31389 35612 31401 35615
rect 31076 35584 31401 35612
rect 31076 35572 31082 35584
rect 31389 35581 31401 35584
rect 31435 35581 31447 35615
rect 31389 35575 31447 35581
rect 31726 35584 33272 35612
rect 31726 35544 31754 35584
rect 33244 35556 33272 35584
rect 33318 35572 33324 35624
rect 33376 35572 33382 35624
rect 33505 35615 33563 35621
rect 33505 35581 33517 35615
rect 33551 35581 33563 35615
rect 33505 35575 33563 35581
rect 34333 35615 34391 35621
rect 34333 35581 34345 35615
rect 34379 35612 34391 35615
rect 34440 35612 34468 35643
rect 35158 35640 35164 35692
rect 35216 35640 35222 35692
rect 35728 35689 35756 35720
rect 35437 35683 35495 35689
rect 35437 35680 35449 35683
rect 35360 35652 35449 35680
rect 34514 35612 34520 35624
rect 34379 35584 34520 35612
rect 34379 35581 34391 35584
rect 34333 35575 34391 35581
rect 30484 35516 31754 35544
rect 33226 35504 33232 35556
rect 33284 35544 33290 35556
rect 33520 35544 33548 35575
rect 34514 35572 34520 35584
rect 34572 35572 34578 35624
rect 35360 35612 35388 35652
rect 35437 35649 35449 35652
rect 35483 35649 35495 35683
rect 35437 35643 35495 35649
rect 35713 35683 35771 35689
rect 35713 35649 35725 35683
rect 35759 35649 35771 35683
rect 35713 35643 35771 35649
rect 35897 35683 35955 35689
rect 35897 35649 35909 35683
rect 35943 35680 35955 35683
rect 36078 35680 36084 35692
rect 35943 35652 36084 35680
rect 35943 35649 35955 35652
rect 35897 35643 35955 35649
rect 36078 35640 36084 35652
rect 36136 35680 36142 35692
rect 36265 35683 36323 35689
rect 36265 35680 36277 35683
rect 36136 35652 36277 35680
rect 36136 35640 36142 35652
rect 36265 35649 36277 35652
rect 36311 35649 36323 35683
rect 36265 35643 36323 35649
rect 35802 35612 35808 35624
rect 35360 35584 35808 35612
rect 33284 35516 33548 35544
rect 33284 35504 33290 35516
rect 25406 35476 25412 35488
rect 23584 35448 25412 35476
rect 25406 35436 25412 35448
rect 25464 35436 25470 35488
rect 26326 35436 26332 35488
rect 26384 35476 26390 35488
rect 26973 35479 27031 35485
rect 26973 35476 26985 35479
rect 26384 35448 26985 35476
rect 26384 35436 26390 35448
rect 26973 35445 26985 35448
rect 27019 35445 27031 35479
rect 26973 35439 27031 35445
rect 29822 35436 29828 35488
rect 29880 35436 29886 35488
rect 32398 35436 32404 35488
rect 32456 35476 32462 35488
rect 32861 35479 32919 35485
rect 32861 35476 32873 35479
rect 32456 35448 32873 35476
rect 32456 35436 32462 35448
rect 32861 35445 32873 35448
rect 32907 35445 32919 35479
rect 33520 35476 33548 35516
rect 34146 35504 34152 35556
rect 34204 35544 34210 35556
rect 35360 35544 35388 35584
rect 35802 35572 35808 35584
rect 35860 35612 35866 35624
rect 35989 35615 36047 35621
rect 35989 35612 36001 35615
rect 35860 35584 36001 35612
rect 35860 35572 35866 35584
rect 35989 35581 36001 35584
rect 36035 35581 36047 35615
rect 35989 35575 36047 35581
rect 36173 35615 36231 35621
rect 36173 35581 36185 35615
rect 36219 35612 36231 35615
rect 36372 35612 36400 35720
rect 38654 35708 38660 35760
rect 38712 35748 38718 35760
rect 39206 35748 39212 35760
rect 38712 35720 39212 35748
rect 38712 35708 38718 35720
rect 39206 35708 39212 35720
rect 39264 35748 39270 35760
rect 39264 35720 39528 35748
rect 39264 35708 39270 35720
rect 38013 35683 38071 35689
rect 38013 35649 38025 35683
rect 38059 35680 38071 35683
rect 38565 35683 38623 35689
rect 38565 35680 38577 35683
rect 38059 35652 38577 35680
rect 38059 35649 38071 35652
rect 38013 35643 38071 35649
rect 38565 35649 38577 35652
rect 38611 35649 38623 35683
rect 38565 35643 38623 35649
rect 38930 35640 38936 35692
rect 38988 35680 38994 35692
rect 39500 35689 39528 35720
rect 39758 35708 39764 35760
rect 39816 35748 39822 35760
rect 40236 35748 40264 35788
rect 41156 35748 41184 35788
rect 41322 35776 41328 35828
rect 41380 35776 41386 35828
rect 41414 35748 41420 35760
rect 39816 35720 40342 35748
rect 41156 35720 41420 35748
rect 39816 35708 39822 35720
rect 41414 35708 41420 35720
rect 41472 35708 41478 35760
rect 39117 35683 39175 35689
rect 39117 35680 39129 35683
rect 38988 35652 39129 35680
rect 38988 35640 38994 35652
rect 39117 35649 39129 35652
rect 39163 35649 39175 35683
rect 39117 35643 39175 35649
rect 39301 35683 39359 35689
rect 39301 35649 39313 35683
rect 39347 35649 39359 35683
rect 39301 35643 39359 35649
rect 39485 35683 39543 35689
rect 39485 35649 39497 35683
rect 39531 35649 39543 35683
rect 39485 35643 39543 35649
rect 36219 35584 36400 35612
rect 36219 35581 36231 35584
rect 36173 35575 36231 35581
rect 38102 35572 38108 35624
rect 38160 35572 38166 35624
rect 38289 35615 38347 35621
rect 38289 35581 38301 35615
rect 38335 35581 38347 35615
rect 38289 35575 38347 35581
rect 34204 35516 35388 35544
rect 34204 35504 34210 35516
rect 35434 35504 35440 35556
rect 35492 35544 35498 35556
rect 36081 35547 36139 35553
rect 36081 35544 36093 35547
rect 35492 35516 36093 35544
rect 35492 35504 35498 35516
rect 36081 35513 36093 35516
rect 36127 35513 36139 35547
rect 38304 35544 38332 35575
rect 38470 35572 38476 35624
rect 38528 35612 38534 35624
rect 39316 35612 39344 35643
rect 39574 35640 39580 35692
rect 39632 35640 39638 35692
rect 38528 35584 39344 35612
rect 38528 35572 38534 35584
rect 38746 35544 38752 35556
rect 38304 35516 38752 35544
rect 36081 35507 36139 35513
rect 38746 35504 38752 35516
rect 38804 35504 38810 35556
rect 34422 35476 34428 35488
rect 33520 35448 34428 35476
rect 32861 35439 32919 35445
rect 34422 35436 34428 35448
rect 34480 35436 34486 35488
rect 34790 35436 34796 35488
rect 34848 35476 34854 35488
rect 34885 35479 34943 35485
rect 34885 35476 34897 35479
rect 34848 35448 34897 35476
rect 34848 35436 34854 35448
rect 34885 35445 34897 35448
rect 34931 35445 34943 35479
rect 34885 35439 34943 35445
rect 35342 35436 35348 35488
rect 35400 35436 35406 35488
rect 37642 35436 37648 35488
rect 37700 35436 37706 35488
rect 39316 35476 39344 35584
rect 39850 35572 39856 35624
rect 39908 35572 39914 35624
rect 41230 35572 41236 35624
rect 41288 35612 41294 35624
rect 41509 35615 41567 35621
rect 41509 35612 41521 35615
rect 41288 35584 41521 35612
rect 41288 35572 41294 35584
rect 41509 35581 41521 35584
rect 41555 35581 41567 35615
rect 41509 35575 41567 35581
rect 40034 35476 40040 35488
rect 39316 35448 40040 35476
rect 40034 35436 40040 35448
rect 40092 35436 40098 35488
rect 42150 35436 42156 35488
rect 42208 35436 42214 35488
rect 1104 35386 42504 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 42504 35386
rect 1104 35312 42504 35334
rect 2958 35232 2964 35284
rect 3016 35272 3022 35284
rect 3145 35275 3203 35281
rect 3145 35272 3157 35275
rect 3016 35244 3157 35272
rect 3016 35232 3022 35244
rect 3145 35241 3157 35244
rect 3191 35241 3203 35275
rect 3145 35235 3203 35241
rect 3973 35275 4031 35281
rect 3973 35241 3985 35275
rect 4019 35272 4031 35275
rect 4062 35272 4068 35284
rect 4019 35244 4068 35272
rect 4019 35241 4031 35244
rect 3973 35235 4031 35241
rect 4062 35232 4068 35244
rect 4120 35232 4126 35284
rect 4709 35275 4767 35281
rect 4709 35241 4721 35275
rect 4755 35272 4767 35275
rect 4890 35272 4896 35284
rect 4755 35244 4896 35272
rect 4755 35241 4767 35244
rect 4709 35235 4767 35241
rect 4724 35136 4752 35235
rect 4890 35232 4896 35244
rect 4948 35272 4954 35284
rect 5350 35272 5356 35284
rect 4948 35244 5356 35272
rect 4948 35232 4954 35244
rect 5350 35232 5356 35244
rect 5408 35232 5414 35284
rect 7101 35275 7159 35281
rect 7101 35241 7113 35275
rect 7147 35272 7159 35275
rect 7374 35272 7380 35284
rect 7147 35244 7380 35272
rect 7147 35241 7159 35244
rect 7101 35235 7159 35241
rect 7374 35232 7380 35244
rect 7432 35232 7438 35284
rect 8205 35275 8263 35281
rect 8205 35241 8217 35275
rect 8251 35241 8263 35275
rect 8205 35235 8263 35241
rect 8665 35275 8723 35281
rect 8665 35241 8677 35275
rect 8711 35272 8723 35275
rect 10502 35272 10508 35284
rect 8711 35244 10508 35272
rect 8711 35241 8723 35244
rect 8665 35235 8723 35241
rect 7006 35164 7012 35216
rect 7064 35204 7070 35216
rect 8021 35207 8079 35213
rect 8021 35204 8033 35207
rect 7064 35176 8033 35204
rect 7064 35164 7070 35176
rect 8021 35173 8033 35176
rect 8067 35173 8079 35207
rect 8220 35204 8248 35235
rect 10502 35232 10508 35244
rect 10560 35232 10566 35284
rect 12250 35232 12256 35284
rect 12308 35232 12314 35284
rect 13170 35232 13176 35284
rect 13228 35272 13234 35284
rect 13630 35272 13636 35284
rect 13228 35244 13636 35272
rect 13228 35232 13234 35244
rect 13630 35232 13636 35244
rect 13688 35272 13694 35284
rect 13725 35275 13783 35281
rect 13725 35272 13737 35275
rect 13688 35244 13737 35272
rect 13688 35232 13694 35244
rect 13725 35241 13737 35244
rect 13771 35241 13783 35275
rect 13725 35235 13783 35241
rect 15197 35275 15255 35281
rect 15197 35241 15209 35275
rect 15243 35272 15255 35275
rect 15562 35272 15568 35284
rect 15243 35244 15568 35272
rect 15243 35241 15255 35244
rect 15197 35235 15255 35241
rect 15562 35232 15568 35244
rect 15620 35232 15626 35284
rect 17310 35232 17316 35284
rect 17368 35272 17374 35284
rect 18138 35272 18144 35284
rect 17368 35244 18144 35272
rect 17368 35232 17374 35244
rect 18138 35232 18144 35244
rect 18196 35232 18202 35284
rect 18230 35232 18236 35284
rect 18288 35272 18294 35284
rect 18509 35275 18567 35281
rect 18509 35272 18521 35275
rect 18288 35244 18521 35272
rect 18288 35232 18294 35244
rect 18509 35241 18521 35244
rect 18555 35241 18567 35275
rect 18509 35235 18567 35241
rect 24670 35232 24676 35284
rect 24728 35272 24734 35284
rect 24857 35275 24915 35281
rect 24857 35272 24869 35275
rect 24728 35244 24869 35272
rect 24728 35232 24734 35244
rect 24857 35241 24869 35244
rect 24903 35241 24915 35275
rect 24857 35235 24915 35241
rect 28629 35275 28687 35281
rect 28629 35241 28641 35275
rect 28675 35272 28687 35275
rect 29270 35272 29276 35284
rect 28675 35244 29276 35272
rect 28675 35241 28687 35244
rect 28629 35235 28687 35241
rect 29270 35232 29276 35244
rect 29328 35232 29334 35284
rect 31018 35232 31024 35284
rect 31076 35272 31082 35284
rect 31297 35275 31355 35281
rect 31297 35272 31309 35275
rect 31076 35244 31309 35272
rect 31076 35232 31082 35244
rect 31297 35241 31309 35244
rect 31343 35241 31355 35275
rect 31297 35235 31355 35241
rect 33873 35275 33931 35281
rect 33873 35241 33885 35275
rect 33919 35272 33931 35275
rect 34514 35272 34520 35284
rect 33919 35244 34520 35272
rect 33919 35241 33931 35244
rect 33873 35235 33931 35241
rect 34514 35232 34520 35244
rect 34572 35232 34578 35284
rect 35342 35232 35348 35284
rect 35400 35272 35406 35284
rect 36357 35275 36415 35281
rect 36357 35272 36369 35275
rect 35400 35244 36369 35272
rect 35400 35232 35406 35244
rect 36357 35241 36369 35244
rect 36403 35241 36415 35275
rect 36357 35235 36415 35241
rect 38654 35232 38660 35284
rect 38712 35272 38718 35284
rect 39758 35272 39764 35284
rect 38712 35244 39764 35272
rect 38712 35232 38718 35244
rect 39758 35232 39764 35244
rect 39816 35232 39822 35284
rect 39850 35232 39856 35284
rect 39908 35272 39914 35284
rect 40129 35275 40187 35281
rect 40129 35272 40141 35275
rect 39908 35244 40141 35272
rect 39908 35232 39914 35244
rect 40129 35241 40141 35244
rect 40175 35241 40187 35275
rect 40129 35235 40187 35241
rect 41414 35232 41420 35284
rect 41472 35272 41478 35284
rect 41969 35275 42027 35281
rect 41969 35272 41981 35275
rect 41472 35244 41981 35272
rect 41472 35232 41478 35244
rect 41969 35241 41981 35244
rect 42015 35241 42027 35275
rect 41969 35235 42027 35241
rect 8938 35204 8944 35216
rect 8220 35176 8944 35204
rect 8021 35167 8079 35173
rect 4172 35108 4752 35136
rect 3326 35028 3332 35080
rect 3384 35028 3390 35080
rect 3510 35028 3516 35080
rect 3568 35028 3574 35080
rect 3605 35071 3663 35077
rect 3605 35037 3617 35071
rect 3651 35068 3663 35071
rect 3878 35068 3884 35080
rect 3651 35040 3884 35068
rect 3651 35037 3663 35040
rect 3605 35031 3663 35037
rect 3878 35028 3884 35040
rect 3936 35068 3942 35080
rect 4062 35068 4068 35080
rect 3936 35040 4068 35068
rect 3936 35028 3942 35040
rect 4062 35028 4068 35040
rect 4120 35028 4126 35080
rect 4172 35077 4200 35108
rect 5534 35096 5540 35148
rect 5592 35096 5598 35148
rect 4157 35071 4215 35077
rect 4157 35037 4169 35071
rect 4203 35037 4215 35071
rect 4157 35031 4215 35037
rect 4433 35071 4491 35077
rect 4433 35037 4445 35071
rect 4479 35037 4491 35071
rect 4433 35031 4491 35037
rect 4448 35000 4476 35031
rect 5258 35028 5264 35080
rect 5316 35028 5322 35080
rect 6914 35028 6920 35080
rect 6972 35068 6978 35080
rect 7285 35071 7343 35077
rect 7285 35068 7297 35071
rect 6972 35040 7297 35068
rect 6972 35028 6978 35040
rect 7285 35037 7297 35040
rect 7331 35068 7343 35071
rect 8036 35068 8064 35167
rect 8938 35164 8944 35176
rect 8996 35164 9002 35216
rect 9030 35164 9036 35216
rect 9088 35204 9094 35216
rect 10778 35204 10784 35216
rect 9088 35176 10784 35204
rect 9088 35164 9094 35176
rect 10778 35164 10784 35176
rect 10836 35164 10842 35216
rect 14182 35204 14188 35216
rect 12728 35176 14188 35204
rect 8481 35071 8539 35077
rect 8481 35068 8493 35071
rect 7331 35040 7972 35068
rect 8036 35040 8493 35068
rect 7331 35037 7343 35040
rect 7285 35031 7343 35037
rect 4706 35009 4712 35012
rect 4693 35003 4712 35009
rect 4693 35000 4705 35003
rect 4448 34972 4705 35000
rect 4693 34969 4705 34972
rect 4693 34963 4712 34969
rect 4706 34960 4712 34963
rect 4764 34960 4770 35012
rect 4798 34960 4804 35012
rect 4856 35000 4862 35012
rect 4893 35003 4951 35009
rect 4893 35000 4905 35003
rect 4856 34972 4905 35000
rect 4856 34960 4862 34972
rect 4893 34969 4905 34972
rect 4939 35000 4951 35003
rect 4982 35000 4988 35012
rect 4939 34972 4988 35000
rect 4939 34969 4951 34972
rect 4893 34963 4951 34969
rect 4982 34960 4988 34972
rect 5040 34960 5046 35012
rect 7098 35000 7104 35012
rect 6762 34972 7104 35000
rect 7098 34960 7104 34972
rect 7156 34960 7162 35012
rect 7469 35003 7527 35009
rect 7469 34969 7481 35003
rect 7515 35000 7527 35003
rect 7742 35000 7748 35012
rect 7515 34972 7748 35000
rect 7515 34969 7527 34972
rect 7469 34963 7527 34969
rect 7742 34960 7748 34972
rect 7800 34960 7806 35012
rect 7944 35000 7972 35040
rect 8481 35037 8493 35040
rect 8527 35037 8539 35071
rect 8481 35031 8539 35037
rect 8665 35071 8723 35077
rect 8665 35037 8677 35071
rect 8711 35068 8723 35071
rect 10594 35068 10600 35080
rect 8711 35040 10600 35068
rect 8711 35037 8723 35040
rect 8665 35031 8723 35037
rect 10594 35028 10600 35040
rect 10652 35028 10658 35080
rect 12434 35028 12440 35080
rect 12492 35028 12498 35080
rect 12728 35077 12756 35176
rect 14182 35164 14188 35176
rect 14240 35164 14246 35216
rect 16666 35204 16672 35216
rect 15672 35176 16672 35204
rect 13814 35096 13820 35148
rect 13872 35136 13878 35148
rect 15672 35145 15700 35176
rect 16666 35164 16672 35176
rect 16724 35164 16730 35216
rect 14093 35139 14151 35145
rect 14093 35136 14105 35139
rect 13872 35108 14105 35136
rect 13872 35096 13878 35108
rect 14093 35105 14105 35108
rect 14139 35105 14151 35139
rect 14093 35099 14151 35105
rect 15657 35139 15715 35145
rect 15657 35105 15669 35139
rect 15703 35105 15715 35139
rect 15657 35099 15715 35105
rect 15841 35139 15899 35145
rect 15841 35105 15853 35139
rect 15887 35136 15899 35139
rect 15930 35136 15936 35148
rect 15887 35108 15936 35136
rect 15887 35105 15899 35108
rect 15841 35099 15899 35105
rect 15930 35096 15936 35108
rect 15988 35096 15994 35148
rect 17126 35096 17132 35148
rect 17184 35096 17190 35148
rect 19981 35139 20039 35145
rect 19981 35136 19993 35139
rect 18708 35108 19993 35136
rect 12713 35071 12771 35077
rect 12713 35037 12725 35071
rect 12759 35037 12771 35071
rect 12713 35031 12771 35037
rect 12897 35071 12955 35077
rect 12897 35037 12909 35071
rect 12943 35037 12955 35071
rect 12897 35031 12955 35037
rect 12989 35071 13047 35077
rect 12989 35037 13001 35071
rect 13035 35068 13047 35071
rect 14642 35068 14648 35080
rect 13035 35040 14648 35068
rect 13035 35037 13047 35040
rect 12989 35031 13047 35037
rect 8389 35003 8447 35009
rect 8389 35000 8401 35003
rect 7944 34972 8401 35000
rect 8389 34969 8401 34972
rect 8435 35000 8447 35003
rect 9030 35000 9036 35012
rect 8435 34972 9036 35000
rect 8435 34969 8447 34972
rect 8389 34963 8447 34969
rect 9030 34960 9036 34972
rect 9088 34960 9094 35012
rect 4341 34935 4399 34941
rect 4341 34901 4353 34935
rect 4387 34932 4399 34935
rect 4430 34932 4436 34944
rect 4387 34904 4436 34932
rect 4387 34901 4399 34904
rect 4341 34895 4399 34901
rect 4430 34892 4436 34904
rect 4488 34892 4494 34944
rect 4522 34892 4528 34944
rect 4580 34892 4586 34944
rect 6822 34892 6828 34944
rect 6880 34932 6886 34944
rect 7009 34935 7067 34941
rect 7009 34932 7021 34935
rect 6880 34904 7021 34932
rect 6880 34892 6886 34904
rect 7009 34901 7021 34904
rect 7055 34901 7067 34935
rect 7760 34932 7788 34960
rect 8179 34935 8237 34941
rect 8179 34932 8191 34935
rect 7760 34904 8191 34932
rect 7009 34895 7067 34901
rect 8179 34901 8191 34904
rect 8225 34932 8237 34935
rect 9306 34932 9312 34944
rect 8225 34904 9312 34932
rect 8225 34901 8237 34904
rect 8179 34895 8237 34901
rect 9306 34892 9312 34904
rect 9364 34932 9370 34944
rect 10870 34932 10876 34944
rect 9364 34904 10876 34932
rect 9364 34892 9370 34904
rect 10870 34892 10876 34904
rect 10928 34892 10934 34944
rect 12912 34932 12940 35031
rect 14642 35028 14648 35040
rect 14700 35028 14706 35080
rect 16022 35028 16028 35080
rect 16080 35028 16086 35080
rect 17396 35071 17454 35077
rect 17396 35037 17408 35071
rect 17442 35068 17454 35071
rect 17678 35068 17684 35080
rect 17442 35040 17684 35068
rect 17442 35037 17454 35040
rect 17396 35031 17454 35037
rect 17678 35028 17684 35040
rect 17736 35028 17742 35080
rect 18598 35028 18604 35080
rect 18656 35068 18662 35080
rect 18708 35077 18736 35108
rect 19981 35105 19993 35108
rect 20027 35105 20039 35139
rect 19981 35099 20039 35105
rect 22005 35139 22063 35145
rect 22005 35105 22017 35139
rect 22051 35136 22063 35139
rect 22094 35136 22100 35148
rect 22051 35108 22100 35136
rect 22051 35105 22063 35108
rect 22005 35099 22063 35105
rect 22094 35096 22100 35108
rect 22152 35136 22158 35148
rect 23014 35136 23020 35148
rect 22152 35108 23020 35136
rect 22152 35096 22158 35108
rect 23014 35096 23020 35108
rect 23072 35096 23078 35148
rect 23382 35096 23388 35148
rect 23440 35096 23446 35148
rect 24762 35096 24768 35148
rect 24820 35136 24826 35148
rect 25409 35139 25467 35145
rect 25409 35136 25421 35139
rect 24820 35108 25421 35136
rect 24820 35096 24826 35108
rect 25409 35105 25421 35108
rect 25455 35105 25467 35139
rect 26326 35136 26332 35148
rect 25409 35099 25467 35105
rect 26151 35108 26332 35136
rect 18693 35071 18751 35077
rect 18693 35068 18705 35071
rect 18656 35040 18705 35068
rect 18656 35028 18662 35040
rect 18693 35037 18705 35040
rect 18739 35037 18751 35071
rect 18693 35031 18751 35037
rect 19797 35071 19855 35077
rect 19797 35037 19809 35071
rect 19843 35037 19855 35071
rect 19797 35031 19855 35037
rect 25225 35071 25283 35077
rect 25225 35037 25237 35071
rect 25271 35068 25283 35071
rect 26151 35068 26179 35108
rect 26326 35096 26332 35108
rect 26384 35096 26390 35148
rect 29288 35145 29316 35232
rect 35802 35164 35808 35216
rect 35860 35204 35866 35216
rect 35860 35176 36124 35204
rect 35860 35164 35866 35176
rect 29273 35139 29331 35145
rect 29273 35105 29285 35139
rect 29319 35105 29331 35139
rect 29273 35099 29331 35105
rect 29822 35096 29828 35148
rect 29880 35096 29886 35148
rect 31478 35096 31484 35148
rect 31536 35136 31542 35148
rect 31941 35139 31999 35145
rect 31941 35136 31953 35139
rect 31536 35108 31953 35136
rect 31536 35096 31542 35108
rect 31941 35105 31953 35108
rect 31987 35105 31999 35139
rect 31941 35099 31999 35105
rect 32122 35096 32128 35148
rect 32180 35096 32186 35148
rect 32398 35096 32404 35148
rect 32456 35096 32462 35148
rect 33410 35096 33416 35148
rect 33468 35136 33474 35148
rect 33468 35108 33824 35136
rect 33468 35096 33474 35108
rect 33796 35080 33824 35108
rect 35986 35096 35992 35148
rect 36044 35096 36050 35148
rect 36096 35145 36124 35176
rect 37090 35164 37096 35216
rect 37148 35204 37154 35216
rect 37148 35176 40264 35204
rect 37148 35164 37154 35176
rect 36081 35139 36139 35145
rect 36081 35105 36093 35139
rect 36127 35105 36139 35139
rect 39117 35139 39175 35145
rect 39117 35136 39129 35139
rect 36081 35099 36139 35105
rect 36188 35108 39129 35136
rect 25271 35040 26179 35068
rect 25271 35037 25283 35040
rect 25225 35031 25283 35037
rect 13170 34960 13176 35012
rect 13228 34960 13234 35012
rect 13354 34960 13360 35012
rect 13412 34960 13418 35012
rect 13817 35003 13875 35009
rect 13817 34969 13829 35003
rect 13863 35000 13875 35003
rect 13906 35000 13912 35012
rect 13863 34972 13912 35000
rect 13863 34969 13875 34972
rect 13817 34963 13875 34969
rect 13906 34960 13912 34972
rect 13964 34960 13970 35012
rect 17218 34960 17224 35012
rect 17276 35000 17282 35012
rect 17770 35000 17776 35012
rect 17276 34972 17776 35000
rect 17276 34960 17282 34972
rect 17770 34960 17776 34972
rect 17828 35000 17834 35012
rect 19812 35000 19840 35031
rect 26234 35028 26240 35080
rect 26292 35028 26298 35080
rect 26881 35071 26939 35077
rect 26881 35037 26893 35071
rect 26927 35037 26939 35071
rect 26881 35031 26939 35037
rect 29549 35071 29607 35077
rect 29549 35037 29561 35071
rect 29595 35037 29607 35071
rect 29549 35031 29607 35037
rect 17828 34972 19840 35000
rect 20248 35003 20306 35009
rect 17828 34960 17834 34972
rect 20248 34969 20260 35003
rect 20294 35000 20306 35003
rect 21821 35003 21879 35009
rect 20294 34972 21496 35000
rect 20294 34969 20306 34972
rect 20248 34963 20306 34969
rect 14090 34932 14096 34944
rect 12912 34904 14096 34932
rect 14090 34892 14096 34904
rect 14148 34932 14154 34944
rect 14458 34932 14464 34944
rect 14148 34904 14464 34932
rect 14148 34892 14154 34904
rect 14458 34892 14464 34904
rect 14516 34932 14522 34944
rect 14737 34935 14795 34941
rect 14737 34932 14749 34935
rect 14516 34904 14749 34932
rect 14516 34892 14522 34904
rect 14737 34901 14749 34904
rect 14783 34901 14795 34935
rect 14737 34895 14795 34901
rect 15565 34935 15623 34941
rect 15565 34901 15577 34935
rect 15611 34932 15623 34935
rect 15838 34932 15844 34944
rect 15611 34904 15844 34932
rect 15611 34901 15623 34904
rect 15565 34895 15623 34901
rect 15838 34892 15844 34904
rect 15896 34892 15902 34944
rect 16666 34892 16672 34944
rect 16724 34892 16730 34944
rect 19150 34892 19156 34944
rect 19208 34932 19214 34944
rect 19245 34935 19303 34941
rect 19245 34932 19257 34935
rect 19208 34904 19257 34932
rect 19208 34892 19214 34904
rect 19245 34901 19257 34904
rect 19291 34901 19303 34935
rect 19245 34895 19303 34901
rect 21358 34892 21364 34944
rect 21416 34892 21422 34944
rect 21468 34941 21496 34972
rect 21821 34969 21833 35003
rect 21867 35000 21879 35003
rect 22186 35000 22192 35012
rect 21867 34972 22192 35000
rect 21867 34969 21879 34972
rect 21821 34963 21879 34969
rect 22186 34960 22192 34972
rect 22244 34960 22250 35012
rect 23293 35003 23351 35009
rect 23293 34969 23305 35003
rect 23339 35000 23351 35003
rect 25685 35003 25743 35009
rect 25685 35000 25697 35003
rect 23339 34972 25697 35000
rect 23339 34969 23351 34972
rect 23293 34963 23351 34969
rect 25685 34969 25697 34972
rect 25731 34969 25743 35003
rect 26896 35000 26924 35031
rect 27062 35000 27068 35012
rect 26896 34972 27068 35000
rect 25685 34963 25743 34969
rect 27062 34960 27068 34972
rect 27120 34960 27126 35012
rect 27154 34960 27160 35012
rect 27212 34960 27218 35012
rect 28810 35000 28816 35012
rect 28382 34972 28816 35000
rect 28810 34960 28816 34972
rect 28868 34960 28874 35012
rect 29564 35000 29592 35031
rect 33502 35028 33508 35080
rect 33560 35028 33566 35080
rect 33778 35028 33784 35080
rect 33836 35068 33842 35080
rect 35253 35071 35311 35077
rect 35253 35068 35265 35071
rect 33836 35040 35265 35068
rect 33836 35028 33842 35040
rect 35253 35037 35265 35040
rect 35299 35037 35311 35071
rect 35253 35031 35311 35037
rect 29730 35000 29736 35012
rect 29564 34972 29736 35000
rect 29730 34960 29736 34972
rect 29788 34960 29794 35012
rect 30282 35000 30288 35012
rect 29840 34972 30288 35000
rect 21453 34935 21511 34941
rect 21453 34901 21465 34935
rect 21499 34901 21511 34935
rect 21453 34895 21511 34901
rect 21910 34892 21916 34944
rect 21968 34892 21974 34944
rect 22830 34892 22836 34944
rect 22888 34892 22894 34944
rect 23198 34892 23204 34944
rect 23256 34892 23262 34944
rect 25314 34892 25320 34944
rect 25372 34892 25378 34944
rect 28718 34892 28724 34944
rect 28776 34892 28782 34944
rect 28828 34932 28856 34960
rect 29840 34932 29868 34972
rect 30282 34960 30288 34972
rect 30340 34960 30346 35012
rect 34422 34960 34428 35012
rect 34480 35000 34486 35012
rect 36188 35000 36216 35108
rect 39117 35105 39129 35108
rect 39163 35105 39175 35139
rect 39117 35099 39175 35105
rect 36998 35028 37004 35080
rect 37056 35028 37062 35080
rect 38289 35071 38347 35077
rect 38289 35037 38301 35071
rect 38335 35068 38347 35071
rect 39574 35068 39580 35080
rect 38335 35040 39580 35068
rect 38335 35037 38347 35040
rect 38289 35031 38347 35037
rect 39574 35028 39580 35040
rect 39632 35028 39638 35080
rect 34480 34972 36216 35000
rect 38933 35003 38991 35009
rect 34480 34960 34486 34972
rect 38933 34969 38945 35003
rect 38979 35000 38991 35003
rect 40126 35000 40132 35012
rect 38979 34972 40132 35000
rect 38979 34969 38991 34972
rect 38933 34963 38991 34969
rect 40126 34960 40132 34972
rect 40184 34960 40190 35012
rect 40236 35000 40264 35176
rect 40310 35096 40316 35148
rect 40368 35136 40374 35148
rect 40681 35139 40739 35145
rect 40681 35136 40693 35139
rect 40368 35108 40693 35136
rect 40368 35096 40374 35108
rect 40681 35105 40693 35108
rect 40727 35105 40739 35139
rect 40681 35099 40739 35105
rect 40497 35071 40555 35077
rect 40497 35037 40509 35071
rect 40543 35068 40555 35071
rect 40770 35068 40776 35080
rect 40543 35040 40776 35068
rect 40543 35037 40555 35040
rect 40497 35031 40555 35037
rect 40770 35028 40776 35040
rect 40828 35028 40834 35080
rect 41322 35028 41328 35080
rect 41380 35068 41386 35080
rect 41509 35071 41567 35077
rect 41509 35068 41521 35071
rect 41380 35040 41521 35068
rect 41380 35028 41386 35040
rect 41509 35037 41521 35040
rect 41555 35037 41567 35071
rect 41509 35031 41567 35037
rect 41782 35028 41788 35080
rect 41840 35028 41846 35080
rect 41800 35000 41828 35028
rect 40236 34972 41828 35000
rect 28828 34904 29868 34932
rect 31386 34892 31392 34944
rect 31444 34892 31450 34944
rect 34330 34892 34336 34944
rect 34388 34932 34394 34944
rect 34701 34935 34759 34941
rect 34701 34932 34713 34935
rect 34388 34904 34713 34932
rect 34388 34892 34394 34904
rect 34701 34901 34713 34904
rect 34747 34901 34759 34935
rect 34701 34895 34759 34901
rect 35342 34892 35348 34944
rect 35400 34932 35406 34944
rect 35529 34935 35587 34941
rect 35529 34932 35541 34935
rect 35400 34904 35541 34932
rect 35400 34892 35406 34904
rect 35529 34901 35541 34904
rect 35575 34901 35587 34935
rect 35529 34895 35587 34901
rect 35897 34935 35955 34941
rect 35897 34901 35909 34935
rect 35943 34932 35955 34935
rect 36262 34932 36268 34944
rect 35943 34904 36268 34932
rect 35943 34901 35955 34904
rect 35897 34895 35955 34901
rect 36262 34892 36268 34904
rect 36320 34892 36326 34944
rect 37550 34892 37556 34944
rect 37608 34932 37614 34944
rect 38565 34935 38623 34941
rect 38565 34932 38577 34935
rect 37608 34904 38577 34932
rect 37608 34892 37614 34904
rect 38565 34901 38577 34904
rect 38611 34901 38623 34935
rect 38565 34895 38623 34901
rect 39022 34892 39028 34944
rect 39080 34892 39086 34944
rect 40586 34892 40592 34944
rect 40644 34892 40650 34944
rect 40954 34892 40960 34944
rect 41012 34892 41018 34944
rect 1104 34842 42504 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 42504 34842
rect 1104 34768 42504 34790
rect 3510 34688 3516 34740
rect 3568 34728 3574 34740
rect 3973 34731 4031 34737
rect 3973 34728 3985 34731
rect 3568 34700 3985 34728
rect 3568 34688 3574 34700
rect 3973 34697 3985 34700
rect 4019 34697 4031 34731
rect 11333 34731 11391 34737
rect 11333 34728 11345 34731
rect 3973 34691 4031 34697
rect 8496 34700 11345 34728
rect 4522 34660 4528 34672
rect 3896 34632 4528 34660
rect 3896 34601 3924 34632
rect 4522 34620 4528 34632
rect 4580 34620 4586 34672
rect 3881 34595 3939 34601
rect 3881 34561 3893 34595
rect 3927 34561 3939 34595
rect 3881 34555 3939 34561
rect 4065 34595 4123 34601
rect 4065 34561 4077 34595
rect 4111 34561 4123 34595
rect 4065 34555 4123 34561
rect 5169 34595 5227 34601
rect 5169 34561 5181 34595
rect 5215 34561 5227 34595
rect 5169 34555 5227 34561
rect 3234 34484 3240 34536
rect 3292 34524 3298 34536
rect 3970 34524 3976 34536
rect 3292 34496 3976 34524
rect 3292 34484 3298 34496
rect 3970 34484 3976 34496
rect 4028 34524 4034 34536
rect 4080 34524 4108 34555
rect 4028 34496 4108 34524
rect 4028 34484 4034 34496
rect 5184 34456 5212 34555
rect 5350 34552 5356 34604
rect 5408 34552 5414 34604
rect 5445 34595 5503 34601
rect 5445 34561 5457 34595
rect 5491 34592 5503 34595
rect 6822 34592 6828 34604
rect 5491 34564 6828 34592
rect 5491 34561 5503 34564
rect 5445 34555 5503 34561
rect 6822 34552 6828 34564
rect 6880 34552 6886 34604
rect 8113 34595 8171 34601
rect 8113 34561 8125 34595
rect 8159 34592 8171 34595
rect 8294 34592 8300 34604
rect 8159 34564 8300 34592
rect 8159 34561 8171 34564
rect 8113 34555 8171 34561
rect 8294 34552 8300 34564
rect 8352 34552 8358 34604
rect 8496 34601 8524 34700
rect 11333 34697 11345 34700
rect 11379 34728 11391 34731
rect 11422 34728 11428 34740
rect 11379 34700 11428 34728
rect 11379 34697 11391 34700
rect 11333 34691 11391 34697
rect 11422 34688 11428 34700
rect 11480 34688 11486 34740
rect 15105 34731 15163 34737
rect 15105 34697 15117 34731
rect 15151 34728 15163 34731
rect 16022 34728 16028 34740
rect 15151 34700 16028 34728
rect 15151 34697 15163 34700
rect 15105 34691 15163 34697
rect 16022 34688 16028 34700
rect 16080 34688 16086 34740
rect 17218 34688 17224 34740
rect 17276 34688 17282 34740
rect 18693 34731 18751 34737
rect 18693 34728 18705 34731
rect 18524 34700 18705 34728
rect 8938 34660 8944 34672
rect 8772 34632 8944 34660
rect 8772 34601 8800 34632
rect 8938 34620 8944 34632
rect 8996 34620 9002 34672
rect 10594 34620 10600 34672
rect 10652 34620 10658 34672
rect 13446 34620 13452 34672
rect 13504 34660 13510 34672
rect 13504 34632 13662 34660
rect 13504 34620 13510 34632
rect 15746 34620 15752 34672
rect 15804 34660 15810 34672
rect 16669 34663 16727 34669
rect 16669 34660 16681 34663
rect 15804 34632 16681 34660
rect 15804 34620 15810 34632
rect 16669 34629 16681 34632
rect 16715 34629 16727 34663
rect 16669 34623 16727 34629
rect 18356 34663 18414 34669
rect 18356 34629 18368 34663
rect 18402 34660 18414 34663
rect 18524 34660 18552 34700
rect 18693 34697 18705 34700
rect 18739 34697 18751 34731
rect 18693 34691 18751 34697
rect 19150 34688 19156 34740
rect 19208 34688 19214 34740
rect 19242 34688 19248 34740
rect 19300 34728 19306 34740
rect 19300 34700 20668 34728
rect 19300 34688 19306 34700
rect 20156 34663 20214 34669
rect 18402 34632 18552 34660
rect 18616 34632 19932 34660
rect 18402 34629 18414 34632
rect 18356 34623 18414 34629
rect 18616 34604 18644 34632
rect 8481 34595 8539 34601
rect 8481 34561 8493 34595
rect 8527 34561 8539 34595
rect 8481 34555 8539 34561
rect 8757 34595 8815 34601
rect 8757 34561 8769 34595
rect 8803 34561 8815 34595
rect 8757 34555 8815 34561
rect 9122 34552 9128 34604
rect 9180 34552 9186 34604
rect 9306 34552 9312 34604
rect 9364 34552 9370 34604
rect 16229 34595 16287 34601
rect 16229 34561 16241 34595
rect 16275 34592 16287 34595
rect 16390 34592 16396 34604
rect 16275 34564 16396 34592
rect 16275 34561 16287 34564
rect 16229 34555 16287 34561
rect 16390 34552 16396 34564
rect 16448 34552 16454 34604
rect 17037 34595 17095 34601
rect 17037 34561 17049 34595
rect 17083 34592 17095 34595
rect 17083 34564 18552 34592
rect 17083 34561 17095 34564
rect 17037 34555 17095 34561
rect 8941 34527 8999 34533
rect 8941 34524 8953 34527
rect 8588 34496 8953 34524
rect 8588 34468 8616 34496
rect 8941 34493 8953 34496
rect 8987 34493 8999 34527
rect 8941 34487 8999 34493
rect 9030 34484 9036 34536
rect 9088 34484 9094 34536
rect 9582 34484 9588 34536
rect 9640 34484 9646 34536
rect 11422 34484 11428 34536
rect 11480 34524 11486 34536
rect 12069 34527 12127 34533
rect 12069 34524 12081 34527
rect 11480 34496 12081 34524
rect 11480 34484 11486 34496
rect 12069 34493 12081 34496
rect 12115 34493 12127 34527
rect 12069 34487 12127 34493
rect 12894 34484 12900 34536
rect 12952 34484 12958 34536
rect 14550 34484 14556 34536
rect 14608 34524 14614 34536
rect 14645 34527 14703 34533
rect 14645 34524 14657 34527
rect 14608 34496 14657 34524
rect 14608 34484 14614 34496
rect 14645 34493 14657 34496
rect 14691 34493 14703 34527
rect 14645 34487 14703 34493
rect 16485 34527 16543 34533
rect 16485 34493 16497 34527
rect 16531 34524 16543 34527
rect 17126 34524 17132 34536
rect 16531 34496 17132 34524
rect 16531 34493 16543 34496
rect 16485 34487 16543 34493
rect 17126 34484 17132 34496
rect 17184 34484 17190 34536
rect 18524 34524 18552 34564
rect 18598 34552 18604 34604
rect 18656 34552 18662 34604
rect 19061 34595 19119 34601
rect 19061 34561 19073 34595
rect 19107 34592 19119 34595
rect 19334 34592 19340 34604
rect 19107 34564 19340 34592
rect 19107 34561 19119 34564
rect 19061 34555 19119 34561
rect 19334 34552 19340 34564
rect 19392 34552 19398 34604
rect 19904 34601 19932 34632
rect 20156 34629 20168 34663
rect 20202 34660 20214 34663
rect 20530 34660 20536 34672
rect 20202 34632 20536 34660
rect 20202 34629 20214 34632
rect 20156 34623 20214 34629
rect 20530 34620 20536 34632
rect 20588 34620 20594 34672
rect 20640 34660 20668 34700
rect 20898 34688 20904 34740
rect 20956 34728 20962 34740
rect 21269 34731 21327 34737
rect 21269 34728 21281 34731
rect 20956 34700 21281 34728
rect 20956 34688 20962 34700
rect 21269 34697 21281 34700
rect 21315 34697 21327 34731
rect 21269 34691 21327 34697
rect 22281 34731 22339 34737
rect 22281 34697 22293 34731
rect 22327 34728 22339 34731
rect 22554 34728 22560 34740
rect 22327 34700 22560 34728
rect 22327 34697 22339 34700
rect 22281 34691 22339 34697
rect 22554 34688 22560 34700
rect 22612 34688 22618 34740
rect 23474 34728 23480 34740
rect 22756 34700 23480 34728
rect 22756 34660 22784 34700
rect 23474 34688 23480 34700
rect 23532 34688 23538 34740
rect 24854 34688 24860 34740
rect 24912 34688 24918 34740
rect 25314 34688 25320 34740
rect 25372 34728 25378 34740
rect 25685 34731 25743 34737
rect 25685 34728 25697 34731
rect 25372 34700 25697 34728
rect 25372 34688 25378 34700
rect 25685 34697 25697 34700
rect 25731 34697 25743 34731
rect 25685 34691 25743 34697
rect 27154 34688 27160 34740
rect 27212 34728 27218 34740
rect 27525 34731 27583 34737
rect 27525 34728 27537 34731
rect 27212 34700 27537 34728
rect 27212 34688 27218 34700
rect 27525 34697 27537 34700
rect 27571 34697 27583 34731
rect 27525 34691 27583 34697
rect 27893 34731 27951 34737
rect 27893 34697 27905 34731
rect 27939 34728 27951 34731
rect 28718 34728 28724 34740
rect 27939 34700 28724 34728
rect 27939 34697 27951 34700
rect 27893 34691 27951 34697
rect 28718 34688 28724 34700
rect 28776 34688 28782 34740
rect 30392 34700 31340 34728
rect 20640 34632 22784 34660
rect 22830 34620 22836 34672
rect 22888 34660 22894 34672
rect 23394 34663 23452 34669
rect 23394 34660 23406 34663
rect 22888 34632 23406 34660
rect 22888 34620 22894 34632
rect 23394 34629 23406 34632
rect 23440 34629 23452 34663
rect 23394 34623 23452 34629
rect 25225 34663 25283 34669
rect 25225 34629 25237 34663
rect 25271 34660 25283 34663
rect 25590 34660 25596 34672
rect 25271 34632 25596 34660
rect 25271 34629 25283 34632
rect 25225 34623 25283 34629
rect 25590 34620 25596 34632
rect 25648 34660 25654 34672
rect 26145 34663 26203 34669
rect 26145 34660 26157 34663
rect 25648 34632 26157 34660
rect 25648 34620 25654 34632
rect 26145 34629 26157 34632
rect 26191 34629 26203 34663
rect 26145 34623 26203 34629
rect 29086 34620 29092 34672
rect 29144 34620 29150 34672
rect 30282 34620 30288 34672
rect 30340 34660 30346 34672
rect 30392 34660 30420 34700
rect 31312 34660 31340 34700
rect 31478 34688 31484 34740
rect 31536 34688 31542 34740
rect 31665 34731 31723 34737
rect 31665 34697 31677 34731
rect 31711 34697 31723 34731
rect 38286 34728 38292 34740
rect 31665 34691 31723 34697
rect 33888 34700 38292 34728
rect 31680 34660 31708 34691
rect 33888 34669 33916 34700
rect 38286 34688 38292 34700
rect 38344 34728 38350 34740
rect 38344 34700 39160 34728
rect 38344 34688 38350 34700
rect 30340 34632 30498 34660
rect 31312 34632 31708 34660
rect 33873 34663 33931 34669
rect 30340 34620 30346 34632
rect 33873 34629 33885 34663
rect 33919 34629 33931 34663
rect 33873 34623 33931 34629
rect 19889 34595 19947 34601
rect 19889 34561 19901 34595
rect 19935 34561 19947 34595
rect 19889 34555 19947 34561
rect 19996 34564 21956 34592
rect 18524 34496 19196 34524
rect 5350 34456 5356 34468
rect 5184 34428 5356 34456
rect 5350 34416 5356 34428
rect 5408 34416 5414 34468
rect 8570 34416 8576 34468
rect 8628 34416 8634 34468
rect 8665 34459 8723 34465
rect 8665 34425 8677 34459
rect 8711 34456 8723 34459
rect 9048 34456 9076 34484
rect 8711 34428 9076 34456
rect 19168 34456 19196 34496
rect 19242 34484 19248 34536
rect 19300 34484 19306 34536
rect 19996 34524 20024 34564
rect 19352 34496 20024 34524
rect 21928 34524 21956 34564
rect 24118 34552 24124 34604
rect 24176 34552 24182 34604
rect 26053 34595 26111 34601
rect 26053 34592 26065 34595
rect 25332 34564 26065 34592
rect 22002 34524 22008 34536
rect 21928 34496 22008 34524
rect 19352 34456 19380 34496
rect 22002 34484 22008 34496
rect 22060 34484 22066 34536
rect 23658 34484 23664 34536
rect 23716 34484 23722 34536
rect 23842 34484 23848 34536
rect 23900 34524 23906 34536
rect 24213 34527 24271 34533
rect 24213 34524 24225 34527
rect 23900 34496 24225 34524
rect 23900 34484 23906 34496
rect 24213 34493 24225 34496
rect 24259 34493 24271 34527
rect 24213 34487 24271 34493
rect 24397 34527 24455 34533
rect 24397 34493 24409 34527
rect 24443 34493 24455 34527
rect 24397 34487 24455 34493
rect 24412 34456 24440 34487
rect 25130 34484 25136 34536
rect 25188 34524 25194 34536
rect 25332 34533 25360 34564
rect 26053 34561 26065 34564
rect 26099 34561 26111 34595
rect 31294 34592 31300 34604
rect 26053 34555 26111 34561
rect 31220 34564 31300 34592
rect 25317 34527 25375 34533
rect 25317 34524 25329 34527
rect 25188 34496 25329 34524
rect 25188 34484 25194 34496
rect 25317 34493 25329 34496
rect 25363 34493 25375 34527
rect 25317 34487 25375 34493
rect 25406 34484 25412 34536
rect 25464 34524 25470 34536
rect 25501 34527 25559 34533
rect 25501 34524 25513 34527
rect 25464 34496 25513 34524
rect 25464 34484 25470 34496
rect 25501 34493 25513 34496
rect 25547 34524 25559 34527
rect 26237 34527 26295 34533
rect 26237 34524 26249 34527
rect 25547 34496 26249 34524
rect 25547 34493 25559 34496
rect 25501 34487 25559 34493
rect 26237 34493 26249 34496
rect 26283 34493 26295 34527
rect 26237 34487 26295 34493
rect 27982 34484 27988 34536
rect 28040 34484 28046 34536
rect 28166 34484 28172 34536
rect 28224 34524 28230 34536
rect 28813 34527 28871 34533
rect 28813 34524 28825 34527
rect 28224 34496 28825 34524
rect 28224 34484 28230 34496
rect 28813 34493 28825 34496
rect 28859 34524 28871 34527
rect 28902 34524 28908 34536
rect 28859 34496 28908 34524
rect 28859 34493 28871 34496
rect 28813 34487 28871 34493
rect 28902 34484 28908 34496
rect 28960 34484 28966 34536
rect 29730 34484 29736 34536
rect 29788 34484 29794 34536
rect 30006 34484 30012 34536
rect 30064 34484 30070 34536
rect 30742 34484 30748 34536
rect 30800 34524 30806 34536
rect 31220 34524 31248 34564
rect 31294 34552 31300 34564
rect 31352 34592 31358 34604
rect 31849 34595 31907 34601
rect 31849 34592 31861 34595
rect 31352 34564 31861 34592
rect 31352 34552 31358 34564
rect 31849 34561 31861 34564
rect 31895 34561 31907 34595
rect 31849 34555 31907 34561
rect 32122 34552 32128 34604
rect 32180 34552 32186 34604
rect 32766 34524 32772 34536
rect 30800 34496 31248 34524
rect 31726 34496 32772 34524
rect 30800 34484 30806 34496
rect 19168 34428 19380 34456
rect 23676 34428 25360 34456
rect 8711 34425 8723 34428
rect 8665 34419 8723 34425
rect 4798 34348 4804 34400
rect 4856 34388 4862 34400
rect 5169 34391 5227 34397
rect 5169 34388 5181 34391
rect 4856 34360 5181 34388
rect 4856 34348 4862 34360
rect 5169 34357 5181 34360
rect 5215 34357 5227 34391
rect 5169 34351 5227 34357
rect 5626 34348 5632 34400
rect 5684 34348 5690 34400
rect 6914 34348 6920 34400
rect 6972 34388 6978 34400
rect 8297 34391 8355 34397
rect 8297 34388 8309 34391
rect 6972 34360 8309 34388
rect 6972 34348 6978 34360
rect 8297 34357 8309 34360
rect 8343 34357 8355 34391
rect 8297 34351 8355 34357
rect 9674 34348 9680 34400
rect 9732 34388 9738 34400
rect 9842 34391 9900 34397
rect 9842 34388 9854 34391
rect 9732 34360 9854 34388
rect 9732 34348 9738 34360
rect 9842 34357 9854 34360
rect 9888 34357 9900 34391
rect 9842 34351 9900 34357
rect 10042 34348 10048 34400
rect 10100 34388 10106 34400
rect 11517 34391 11575 34397
rect 11517 34388 11529 34391
rect 10100 34360 11529 34388
rect 10100 34348 10106 34360
rect 11517 34357 11529 34360
rect 11563 34357 11575 34391
rect 11517 34351 11575 34357
rect 13160 34391 13218 34397
rect 13160 34357 13172 34391
rect 13206 34388 13218 34391
rect 13906 34388 13912 34400
rect 13206 34360 13912 34388
rect 13206 34357 13218 34360
rect 13160 34351 13218 34357
rect 13906 34348 13912 34360
rect 13964 34348 13970 34400
rect 23014 34348 23020 34400
rect 23072 34388 23078 34400
rect 23676 34388 23704 34428
rect 25332 34400 25360 34428
rect 31110 34416 31116 34468
rect 31168 34456 31174 34468
rect 31726 34456 31754 34496
rect 32766 34484 32772 34496
rect 32824 34524 32830 34536
rect 33888 34524 33916 34623
rect 34330 34620 34336 34672
rect 34388 34620 34394 34672
rect 34422 34620 34428 34672
rect 34480 34620 34486 34672
rect 34790 34620 34796 34672
rect 34848 34660 34854 34672
rect 35069 34663 35127 34669
rect 35069 34660 35081 34663
rect 34848 34632 35081 34660
rect 34848 34620 34854 34632
rect 35069 34629 35081 34632
rect 35115 34629 35127 34663
rect 35069 34623 35127 34629
rect 35526 34620 35532 34672
rect 35584 34620 35590 34672
rect 37001 34663 37059 34669
rect 37001 34629 37013 34663
rect 37047 34660 37059 34663
rect 37090 34660 37096 34672
rect 37047 34632 37096 34660
rect 37047 34629 37059 34632
rect 37001 34623 37059 34629
rect 37090 34620 37096 34632
rect 37148 34620 37154 34672
rect 37553 34663 37611 34669
rect 37553 34629 37565 34663
rect 37599 34660 37611 34663
rect 37642 34660 37648 34672
rect 37599 34632 37648 34660
rect 37599 34629 37611 34632
rect 37553 34623 37611 34629
rect 37642 34620 37648 34632
rect 37700 34620 37706 34672
rect 34440 34592 34468 34620
rect 39132 34604 39160 34700
rect 40126 34688 40132 34740
rect 40184 34688 40190 34740
rect 40865 34731 40923 34737
rect 40865 34697 40877 34731
rect 40911 34728 40923 34731
rect 41138 34728 41144 34740
rect 40911 34700 41144 34728
rect 40911 34697 40923 34700
rect 40865 34691 40923 34697
rect 41138 34688 41144 34700
rect 41196 34688 41202 34740
rect 41230 34688 41236 34740
rect 41288 34688 41294 34740
rect 41322 34688 41328 34740
rect 41380 34688 41386 34740
rect 39574 34620 39580 34672
rect 39632 34660 39638 34672
rect 39853 34663 39911 34669
rect 39853 34660 39865 34663
rect 39632 34632 39865 34660
rect 39632 34620 39638 34632
rect 39853 34629 39865 34632
rect 39899 34629 39911 34663
rect 39853 34623 39911 34629
rect 41690 34620 41696 34672
rect 41748 34620 41754 34672
rect 34440 34564 34560 34592
rect 32824 34496 33916 34524
rect 32824 34484 32830 34496
rect 34422 34484 34428 34536
rect 34480 34484 34486 34536
rect 34532 34533 34560 34564
rect 38654 34552 38660 34604
rect 38712 34552 38718 34604
rect 39114 34552 39120 34604
rect 39172 34552 39178 34604
rect 39206 34552 39212 34604
rect 39264 34592 39270 34604
rect 40681 34595 40739 34601
rect 40681 34592 40693 34595
rect 39264 34564 40693 34592
rect 39264 34552 39270 34564
rect 40681 34561 40693 34564
rect 40727 34561 40739 34595
rect 40681 34555 40739 34561
rect 34517 34527 34575 34533
rect 34517 34493 34529 34527
rect 34563 34493 34575 34527
rect 34517 34487 34575 34493
rect 34790 34484 34796 34536
rect 34848 34484 34854 34536
rect 35526 34524 35532 34536
rect 34900 34496 35532 34524
rect 31168 34428 31754 34456
rect 31168 34416 31174 34428
rect 33502 34416 33508 34468
rect 33560 34456 33566 34468
rect 34900 34456 34928 34496
rect 35526 34484 35532 34496
rect 35584 34484 35590 34536
rect 35618 34484 35624 34536
rect 35676 34524 35682 34536
rect 37274 34524 37280 34536
rect 35676 34496 37280 34524
rect 35676 34484 35682 34496
rect 37274 34484 37280 34496
rect 37332 34484 37338 34536
rect 38930 34484 38936 34536
rect 38988 34524 38994 34536
rect 39025 34527 39083 34533
rect 39025 34524 39037 34527
rect 38988 34496 39037 34524
rect 38988 34484 38994 34496
rect 39025 34493 39037 34496
rect 39071 34493 39083 34527
rect 39025 34487 39083 34493
rect 41509 34527 41567 34533
rect 41509 34493 41521 34527
rect 41555 34524 41567 34527
rect 41708 34524 41736 34620
rect 41874 34552 41880 34604
rect 41932 34552 41938 34604
rect 41555 34496 41736 34524
rect 41555 34493 41567 34496
rect 41509 34487 41567 34493
rect 33560 34428 34928 34456
rect 36541 34459 36599 34465
rect 33560 34416 33566 34428
rect 36541 34425 36553 34459
rect 36587 34456 36599 34459
rect 36998 34456 37004 34468
rect 36587 34428 37004 34456
rect 36587 34425 36599 34428
rect 36541 34419 36599 34425
rect 36998 34416 37004 34428
rect 37056 34416 37062 34468
rect 23072 34360 23704 34388
rect 23072 34348 23078 34360
rect 23750 34348 23756 34400
rect 23808 34348 23814 34400
rect 25314 34348 25320 34400
rect 25372 34348 25378 34400
rect 33962 34348 33968 34400
rect 34020 34348 34026 34400
rect 35526 34348 35532 34400
rect 35584 34388 35590 34400
rect 36725 34391 36783 34397
rect 36725 34388 36737 34391
rect 35584 34360 36737 34388
rect 35584 34348 35590 34360
rect 36725 34357 36737 34360
rect 36771 34357 36783 34391
rect 36725 34351 36783 34357
rect 1104 34298 42504 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 42504 34298
rect 1104 34224 42504 34246
rect 5626 34144 5632 34196
rect 5684 34184 5690 34196
rect 6089 34187 6147 34193
rect 6089 34184 6101 34187
rect 5684 34156 6101 34184
rect 5684 34144 5690 34156
rect 6089 34153 6101 34156
rect 6135 34153 6147 34187
rect 6089 34147 6147 34153
rect 8481 34187 8539 34193
rect 8481 34153 8493 34187
rect 8527 34184 8539 34187
rect 8570 34184 8576 34196
rect 8527 34156 8576 34184
rect 8527 34153 8539 34156
rect 8481 34147 8539 34153
rect 8570 34144 8576 34156
rect 8628 34144 8634 34196
rect 9674 34144 9680 34196
rect 9732 34144 9738 34196
rect 9766 34144 9772 34196
rect 9824 34184 9830 34196
rect 10594 34184 10600 34196
rect 9824 34156 10600 34184
rect 9824 34144 9830 34156
rect 10594 34144 10600 34156
rect 10652 34144 10658 34196
rect 11146 34144 11152 34196
rect 11204 34184 11210 34196
rect 11422 34184 11428 34196
rect 11204 34156 11428 34184
rect 11204 34144 11210 34156
rect 11422 34144 11428 34156
rect 11480 34184 11486 34196
rect 11517 34187 11575 34193
rect 11517 34184 11529 34187
rect 11480 34156 11529 34184
rect 11480 34144 11486 34156
rect 11517 34153 11529 34156
rect 11563 34153 11575 34187
rect 11517 34147 11575 34153
rect 13725 34187 13783 34193
rect 13725 34153 13737 34187
rect 13771 34184 13783 34187
rect 13814 34184 13820 34196
rect 13771 34156 13820 34184
rect 13771 34153 13783 34156
rect 13725 34147 13783 34153
rect 13814 34144 13820 34156
rect 13872 34144 13878 34196
rect 13906 34144 13912 34196
rect 13964 34184 13970 34196
rect 14093 34187 14151 34193
rect 14093 34184 14105 34187
rect 13964 34156 14105 34184
rect 13964 34144 13970 34156
rect 14093 34153 14105 34156
rect 14139 34153 14151 34187
rect 14093 34147 14151 34153
rect 16390 34144 16396 34196
rect 16448 34144 16454 34196
rect 19242 34144 19248 34196
rect 19300 34144 19306 34196
rect 20990 34144 20996 34196
rect 21048 34144 21054 34196
rect 25866 34144 25872 34196
rect 25924 34144 25930 34196
rect 27706 34144 27712 34196
rect 27764 34184 27770 34196
rect 27893 34187 27951 34193
rect 27893 34184 27905 34187
rect 27764 34156 27905 34184
rect 27764 34144 27770 34156
rect 27893 34153 27905 34156
rect 27939 34153 27951 34187
rect 27893 34147 27951 34153
rect 30190 34144 30196 34196
rect 30248 34144 30254 34196
rect 33042 34144 33048 34196
rect 33100 34184 33106 34196
rect 33100 34156 33364 34184
rect 33100 34144 33106 34156
rect 9122 34076 9128 34128
rect 9180 34116 9186 34128
rect 11333 34119 11391 34125
rect 11333 34116 11345 34119
rect 9180 34088 11345 34116
rect 9180 34076 9186 34088
rect 5258 34008 5264 34060
rect 5316 34048 5322 34060
rect 6733 34051 6791 34057
rect 6733 34048 6745 34051
rect 5316 34020 6745 34048
rect 5316 34008 5322 34020
rect 6733 34017 6745 34020
rect 6779 34048 6791 34051
rect 8294 34048 8300 34060
rect 6779 34020 8300 34048
rect 6779 34017 6791 34020
rect 6733 34011 6791 34017
rect 8294 34008 8300 34020
rect 8352 34008 8358 34060
rect 8570 34008 8576 34060
rect 8628 34048 8634 34060
rect 9493 34051 9551 34057
rect 9493 34048 9505 34051
rect 8628 34020 9505 34048
rect 8628 34008 8634 34020
rect 9493 34017 9505 34020
rect 9539 34017 9551 34051
rect 9493 34011 9551 34017
rect 10042 34008 10048 34060
rect 10100 34008 10106 34060
rect 5902 33940 5908 33992
rect 5960 33940 5966 33992
rect 6181 33983 6239 33989
rect 6181 33949 6193 33983
rect 6227 33949 6239 33983
rect 9766 33980 9772 33992
rect 8142 33952 9772 33980
rect 6181 33943 6239 33949
rect 6196 33912 6224 33943
rect 9766 33940 9772 33952
rect 9824 33940 9830 33992
rect 9858 33940 9864 33992
rect 9916 33940 9922 33992
rect 9953 33983 10011 33989
rect 9953 33949 9965 33983
rect 9999 33980 10011 33983
rect 10060 33980 10088 34008
rect 10336 33989 10364 34088
rect 11333 34085 11345 34088
rect 11379 34085 11391 34119
rect 11333 34079 11391 34085
rect 15749 34119 15807 34125
rect 15749 34085 15761 34119
rect 15795 34116 15807 34119
rect 17494 34116 17500 34128
rect 15795 34088 17500 34116
rect 15795 34085 15807 34088
rect 15749 34079 15807 34085
rect 17494 34076 17500 34088
rect 17552 34076 17558 34128
rect 19260 34116 19288 34144
rect 18064 34088 19288 34116
rect 10962 34008 10968 34060
rect 11020 34048 11026 34060
rect 11149 34051 11207 34057
rect 11149 34048 11161 34051
rect 11020 34020 11161 34048
rect 11020 34008 11026 34020
rect 11149 34017 11161 34020
rect 11195 34017 11207 34051
rect 11149 34011 11207 34017
rect 11977 34051 12035 34057
rect 11977 34017 11989 34051
rect 12023 34048 12035 34051
rect 12894 34048 12900 34060
rect 12023 34020 12900 34048
rect 12023 34017 12035 34020
rect 11977 34011 12035 34017
rect 9999 33952 10088 33980
rect 10229 33983 10287 33989
rect 9999 33949 10011 33952
rect 9953 33943 10011 33949
rect 10229 33949 10241 33983
rect 10275 33949 10287 33983
rect 10229 33943 10287 33949
rect 10321 33983 10379 33989
rect 10321 33949 10333 33983
rect 10367 33949 10379 33983
rect 10321 33943 10379 33949
rect 10505 33983 10563 33989
rect 10505 33949 10517 33983
rect 10551 33980 10563 33983
rect 11054 33980 11060 33992
rect 10551 33952 11060 33980
rect 10551 33949 10563 33952
rect 10505 33943 10563 33949
rect 6914 33912 6920 33924
rect 6196 33884 6920 33912
rect 6914 33872 6920 33884
rect 6972 33872 6978 33924
rect 7006 33872 7012 33924
rect 7064 33872 7070 33924
rect 8662 33872 8668 33924
rect 8720 33912 8726 33924
rect 10045 33915 10103 33921
rect 10045 33912 10057 33915
rect 8720 33884 10057 33912
rect 8720 33872 8726 33884
rect 10045 33881 10057 33884
rect 10091 33881 10103 33915
rect 10244 33912 10272 33943
rect 11054 33940 11060 33952
rect 11112 33940 11118 33992
rect 10413 33915 10471 33921
rect 10413 33912 10425 33915
rect 10244 33884 10425 33912
rect 10045 33875 10103 33881
rect 10413 33881 10425 33884
rect 10459 33881 10471 33915
rect 11164 33912 11192 34011
rect 12894 34008 12900 34020
rect 12952 34008 12958 34060
rect 13446 34008 13452 34060
rect 13504 34008 13510 34060
rect 14642 34008 14648 34060
rect 14700 34008 14706 34060
rect 16482 34048 16488 34060
rect 15672 34020 16488 34048
rect 13464 33980 13492 34008
rect 15672 33992 15700 34020
rect 16482 34008 16488 34020
rect 16540 34008 16546 34060
rect 16666 34008 16672 34060
rect 16724 34048 16730 34060
rect 16853 34051 16911 34057
rect 16853 34048 16865 34051
rect 16724 34020 16865 34048
rect 16724 34008 16730 34020
rect 16853 34017 16865 34020
rect 16899 34017 16911 34051
rect 16853 34011 16911 34017
rect 17034 34008 17040 34060
rect 17092 34048 17098 34060
rect 18064 34048 18092 34088
rect 17092 34020 18092 34048
rect 17092 34008 17098 34020
rect 18598 34008 18604 34060
rect 18656 34048 18662 34060
rect 19245 34051 19303 34057
rect 19245 34048 19257 34051
rect 18656 34020 19257 34048
rect 18656 34008 18662 34020
rect 19245 34017 19257 34020
rect 19291 34017 19303 34051
rect 21008 34048 21036 34144
rect 33336 34116 33364 34156
rect 33778 34144 33784 34196
rect 33836 34144 33842 34196
rect 39025 34187 39083 34193
rect 33888 34156 38608 34184
rect 33888 34116 33916 34156
rect 33336 34088 33916 34116
rect 38580 34116 38608 34156
rect 39025 34153 39037 34187
rect 39071 34184 39083 34187
rect 39206 34184 39212 34196
rect 39071 34156 39212 34184
rect 39071 34153 39083 34156
rect 39025 34147 39083 34153
rect 39206 34144 39212 34156
rect 39264 34144 39270 34196
rect 40586 34144 40592 34196
rect 40644 34184 40650 34196
rect 40957 34187 41015 34193
rect 40957 34184 40969 34187
rect 40644 34156 40969 34184
rect 40644 34144 40650 34156
rect 40957 34153 40969 34156
rect 41003 34153 41015 34187
rect 40957 34147 41015 34153
rect 41966 34116 41972 34128
rect 38580 34088 41972 34116
rect 41966 34076 41972 34088
rect 42024 34076 42030 34128
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 21008 34020 21649 34048
rect 19245 34011 19303 34017
rect 21637 34017 21649 34020
rect 21683 34017 21695 34051
rect 21637 34011 21695 34017
rect 26418 34008 26424 34060
rect 26476 34048 26482 34060
rect 28445 34051 28503 34057
rect 28445 34048 28457 34051
rect 26476 34020 28457 34048
rect 26476 34008 26482 34020
rect 28445 34017 28457 34020
rect 28491 34017 28503 34051
rect 28445 34011 28503 34017
rect 30834 34008 30840 34060
rect 30892 34048 30898 34060
rect 31662 34048 31668 34060
rect 30892 34020 31668 34048
rect 30892 34008 30898 34020
rect 31662 34008 31668 34020
rect 31720 34008 31726 34060
rect 32030 34008 32036 34060
rect 32088 34008 32094 34060
rect 32309 34051 32367 34057
rect 32309 34017 32321 34051
rect 32355 34048 32367 34051
rect 33962 34048 33968 34060
rect 32355 34020 33968 34048
rect 32355 34017 32367 34020
rect 32309 34011 32367 34017
rect 33962 34008 33968 34020
rect 34020 34008 34026 34060
rect 34790 34008 34796 34060
rect 34848 34048 34854 34060
rect 34977 34051 35035 34057
rect 34977 34048 34989 34051
rect 34848 34020 34989 34048
rect 34848 34008 34854 34020
rect 34977 34017 34989 34020
rect 35023 34048 35035 34051
rect 35618 34048 35624 34060
rect 35023 34020 35624 34048
rect 35023 34017 35035 34020
rect 34977 34011 35035 34017
rect 35618 34008 35624 34020
rect 35676 34008 35682 34060
rect 37274 34008 37280 34060
rect 37332 34048 37338 34060
rect 39574 34048 39580 34060
rect 37332 34020 39580 34048
rect 37332 34008 37338 34020
rect 39574 34008 39580 34020
rect 39632 34008 39638 34060
rect 40678 34008 40684 34060
rect 40736 34008 40742 34060
rect 41601 34051 41659 34057
rect 41601 34017 41613 34051
rect 41647 34048 41659 34051
rect 41690 34048 41696 34060
rect 41647 34020 41696 34048
rect 41647 34017 41659 34020
rect 41601 34011 41659 34017
rect 41690 34008 41696 34020
rect 41748 34008 41754 34060
rect 13386 33952 13492 33980
rect 14458 33940 14464 33992
rect 14516 33940 14522 33992
rect 14550 33940 14556 33992
rect 14608 33980 14614 33992
rect 15473 33983 15531 33989
rect 15473 33980 15485 33983
rect 14608 33952 15485 33980
rect 14608 33940 14614 33952
rect 15473 33949 15485 33952
rect 15519 33949 15531 33983
rect 15473 33943 15531 33949
rect 15654 33940 15660 33992
rect 15712 33940 15718 33992
rect 15838 33940 15844 33992
rect 15896 33940 15902 33992
rect 22094 33940 22100 33992
rect 22152 33940 22158 33992
rect 23569 33983 23627 33989
rect 23569 33949 23581 33983
rect 23615 33980 23627 33983
rect 23658 33980 23664 33992
rect 23615 33952 23664 33980
rect 23615 33949 23627 33952
rect 23569 33943 23627 33949
rect 23658 33940 23664 33952
rect 23716 33980 23722 33992
rect 24394 33980 24400 33992
rect 23716 33952 24400 33980
rect 23716 33940 23722 33952
rect 24394 33940 24400 33952
rect 24452 33940 24458 33992
rect 31021 33983 31079 33989
rect 31021 33980 31033 33983
rect 26712 33952 31033 33980
rect 26712 33924 26740 33952
rect 31021 33949 31033 33952
rect 31067 33980 31079 33983
rect 31110 33980 31116 33992
rect 31067 33952 31116 33980
rect 31067 33949 31079 33952
rect 31021 33943 31079 33949
rect 31110 33940 31116 33952
rect 31168 33940 31174 33992
rect 33410 33940 33416 33992
rect 33468 33940 33474 33992
rect 38654 33940 38660 33992
rect 38712 33940 38718 33992
rect 40589 33983 40647 33989
rect 40589 33949 40601 33983
rect 40635 33980 40647 33983
rect 40954 33980 40960 33992
rect 40635 33952 40960 33980
rect 40635 33949 40647 33952
rect 40589 33943 40647 33949
rect 40954 33940 40960 33952
rect 41012 33940 41018 33992
rect 41322 33940 41328 33992
rect 41380 33940 41386 33992
rect 11701 33915 11759 33921
rect 11701 33912 11713 33915
rect 11164 33884 11713 33912
rect 10413 33875 10471 33881
rect 11701 33881 11713 33884
rect 11747 33881 11759 33915
rect 11701 33875 11759 33881
rect 12253 33915 12311 33921
rect 12253 33881 12265 33915
rect 12299 33912 12311 33915
rect 12526 33912 12532 33924
rect 12299 33884 12532 33912
rect 12299 33881 12311 33884
rect 12253 33875 12311 33881
rect 12526 33872 12532 33884
rect 12584 33872 12590 33924
rect 19521 33915 19579 33921
rect 19521 33881 19533 33915
rect 19567 33912 19579 33915
rect 19794 33912 19800 33924
rect 19567 33884 19800 33912
rect 19567 33881 19579 33884
rect 19521 33875 19579 33881
rect 19794 33872 19800 33884
rect 19852 33872 19858 33924
rect 21450 33912 21456 33924
rect 20746 33884 21456 33912
rect 21450 33872 21456 33884
rect 21508 33912 21514 33924
rect 23324 33915 23382 33921
rect 21508 33884 21956 33912
rect 21508 33872 21514 33884
rect 5718 33804 5724 33856
rect 5776 33804 5782 33856
rect 8938 33804 8944 33856
rect 8996 33804 9002 33856
rect 10134 33804 10140 33856
rect 10192 33844 10198 33856
rect 10597 33847 10655 33853
rect 10597 33844 10609 33847
rect 10192 33816 10609 33844
rect 10192 33804 10198 33816
rect 10597 33813 10609 33816
rect 10643 33813 10655 33847
rect 10597 33807 10655 33813
rect 11330 33804 11336 33856
rect 11388 33844 11394 33856
rect 11491 33847 11549 33853
rect 11491 33844 11503 33847
rect 11388 33816 11503 33844
rect 11388 33804 11394 33816
rect 11491 33813 11503 33816
rect 11537 33813 11549 33847
rect 11491 33807 11549 33813
rect 14553 33847 14611 33853
rect 14553 33813 14565 33847
rect 14599 33844 14611 33847
rect 14921 33847 14979 33853
rect 14921 33844 14933 33847
rect 14599 33816 14933 33844
rect 14599 33813 14611 33816
rect 14553 33807 14611 33813
rect 14921 33813 14933 33816
rect 14967 33813 14979 33847
rect 14921 33807 14979 33813
rect 16761 33847 16819 33853
rect 16761 33813 16773 33847
rect 16807 33844 16819 33847
rect 17310 33844 17316 33856
rect 16807 33816 17316 33844
rect 16807 33813 16819 33816
rect 16761 33807 16819 33813
rect 17310 33804 17316 33816
rect 17368 33804 17374 33856
rect 21082 33804 21088 33856
rect 21140 33804 21146 33856
rect 21928 33853 21956 33884
rect 23324 33881 23336 33915
rect 23370 33912 23382 33915
rect 23934 33912 23940 33924
rect 23370 33884 23940 33912
rect 23370 33881 23382 33884
rect 23324 33875 23382 33881
rect 23934 33872 23940 33884
rect 23992 33872 23998 33924
rect 24664 33915 24722 33921
rect 24664 33881 24676 33915
rect 24710 33912 24722 33915
rect 24762 33912 24768 33924
rect 24710 33884 24768 33912
rect 24710 33881 24722 33884
rect 24664 33875 24722 33881
rect 24762 33872 24768 33884
rect 24820 33872 24826 33924
rect 26694 33872 26700 33924
rect 26752 33872 26758 33924
rect 27062 33872 27068 33924
rect 27120 33912 27126 33924
rect 27433 33915 27491 33921
rect 27433 33912 27445 33915
rect 27120 33884 27445 33912
rect 27120 33872 27126 33884
rect 27433 33881 27445 33884
rect 27479 33881 27491 33915
rect 27433 33875 27491 33881
rect 28261 33915 28319 33921
rect 28261 33881 28273 33915
rect 28307 33912 28319 33915
rect 28718 33912 28724 33924
rect 28307 33884 28724 33912
rect 28307 33881 28319 33884
rect 28261 33875 28319 33881
rect 28718 33872 28724 33884
rect 28776 33872 28782 33924
rect 30561 33915 30619 33921
rect 30561 33881 30573 33915
rect 30607 33912 30619 33915
rect 31570 33912 31576 33924
rect 30607 33884 31576 33912
rect 30607 33881 30619 33884
rect 30561 33875 30619 33881
rect 31570 33872 31576 33884
rect 31628 33872 31634 33924
rect 35253 33915 35311 33921
rect 35253 33881 35265 33915
rect 35299 33912 35311 33915
rect 35342 33912 35348 33924
rect 35299 33884 35348 33912
rect 35299 33881 35311 33884
rect 35253 33875 35311 33881
rect 35342 33872 35348 33884
rect 35400 33872 35406 33924
rect 35526 33872 35532 33924
rect 35584 33912 35590 33924
rect 35584 33884 35742 33912
rect 35584 33872 35590 33884
rect 37550 33872 37556 33924
rect 37608 33872 37614 33924
rect 41874 33912 41880 33924
rect 38856 33884 41880 33912
rect 21913 33847 21971 33853
rect 21913 33813 21925 33847
rect 21959 33813 21971 33847
rect 21913 33807 21971 33813
rect 22189 33847 22247 33853
rect 22189 33813 22201 33847
rect 22235 33844 22247 33847
rect 22370 33844 22376 33856
rect 22235 33816 22376 33844
rect 22235 33813 22247 33816
rect 22189 33807 22247 33813
rect 22370 33804 22376 33816
rect 22428 33844 22434 33856
rect 23198 33844 23204 33856
rect 22428 33816 23204 33844
rect 22428 33804 22434 33816
rect 23198 33804 23204 33816
rect 23256 33804 23262 33856
rect 25130 33804 25136 33856
rect 25188 33844 25194 33856
rect 25777 33847 25835 33853
rect 25777 33844 25789 33847
rect 25188 33816 25789 33844
rect 25188 33804 25194 33816
rect 25777 33813 25789 33816
rect 25823 33813 25835 33847
rect 25777 33807 25835 33813
rect 26234 33804 26240 33856
rect 26292 33804 26298 33856
rect 26326 33804 26332 33856
rect 26384 33804 26390 33856
rect 28350 33804 28356 33856
rect 28408 33804 28414 33856
rect 30653 33847 30711 33853
rect 30653 33813 30665 33847
rect 30699 33844 30711 33847
rect 31478 33844 31484 33856
rect 30699 33816 31484 33844
rect 30699 33813 30711 33816
rect 30653 33807 30711 33813
rect 31478 33804 31484 33816
rect 31536 33804 31542 33856
rect 36722 33804 36728 33856
rect 36780 33804 36786 33856
rect 36814 33804 36820 33856
rect 36872 33844 36878 33856
rect 38856 33844 38884 33884
rect 41874 33872 41880 33884
rect 41932 33872 41938 33924
rect 36872 33816 38884 33844
rect 40129 33847 40187 33853
rect 36872 33804 36878 33816
rect 40129 33813 40141 33847
rect 40175 33844 40187 33847
rect 40218 33844 40224 33856
rect 40175 33816 40224 33844
rect 40175 33813 40187 33816
rect 40129 33807 40187 33813
rect 40218 33804 40224 33816
rect 40276 33804 40282 33856
rect 40494 33804 40500 33856
rect 40552 33804 40558 33856
rect 41230 33804 41236 33856
rect 41288 33844 41294 33856
rect 41417 33847 41475 33853
rect 41417 33844 41429 33847
rect 41288 33816 41429 33844
rect 41288 33804 41294 33816
rect 41417 33813 41429 33816
rect 41463 33813 41475 33847
rect 41417 33807 41475 33813
rect 1104 33754 42504 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 42504 33754
rect 1104 33680 42504 33702
rect 3234 33640 3240 33652
rect 2332 33612 3240 33640
rect 2332 33581 2360 33612
rect 3234 33600 3240 33612
rect 3292 33600 3298 33652
rect 10962 33600 10968 33652
rect 11020 33640 11026 33652
rect 11241 33643 11299 33649
rect 11241 33640 11253 33643
rect 11020 33612 11253 33640
rect 11020 33600 11026 33612
rect 11241 33609 11253 33612
rect 11287 33609 11299 33643
rect 11241 33603 11299 33609
rect 12434 33600 12440 33652
rect 12492 33640 12498 33652
rect 12897 33643 12955 33649
rect 12897 33640 12909 33643
rect 12492 33612 12909 33640
rect 12492 33600 12498 33612
rect 12897 33609 12909 33612
rect 12943 33609 12955 33643
rect 12897 33603 12955 33609
rect 16574 33600 16580 33652
rect 16632 33640 16638 33652
rect 16669 33643 16727 33649
rect 16669 33640 16681 33643
rect 16632 33612 16681 33640
rect 16632 33600 16638 33612
rect 16669 33609 16681 33612
rect 16715 33609 16727 33643
rect 16669 33603 16727 33609
rect 18598 33600 18604 33652
rect 18656 33600 18662 33652
rect 19794 33600 19800 33652
rect 19852 33600 19858 33652
rect 20257 33643 20315 33649
rect 20257 33609 20269 33643
rect 20303 33640 20315 33643
rect 21082 33640 21088 33652
rect 20303 33612 21088 33640
rect 20303 33609 20315 33612
rect 20257 33603 20315 33609
rect 21082 33600 21088 33612
rect 21140 33600 21146 33652
rect 21821 33643 21879 33649
rect 21821 33609 21833 33643
rect 21867 33640 21879 33643
rect 21910 33640 21916 33652
rect 21867 33612 21916 33640
rect 21867 33609 21879 33612
rect 21821 33603 21879 33609
rect 21910 33600 21916 33612
rect 21968 33600 21974 33652
rect 23842 33600 23848 33652
rect 23900 33600 23906 33652
rect 23934 33600 23940 33652
rect 23992 33600 23998 33652
rect 24762 33600 24768 33652
rect 24820 33600 24826 33652
rect 26786 33600 26792 33652
rect 26844 33640 26850 33652
rect 26973 33643 27031 33649
rect 26973 33640 26985 33643
rect 26844 33612 26985 33640
rect 26844 33600 26850 33612
rect 26973 33609 26985 33612
rect 27019 33609 27031 33643
rect 26973 33603 27031 33609
rect 27893 33643 27951 33649
rect 27893 33609 27905 33643
rect 27939 33640 27951 33643
rect 27982 33640 27988 33652
rect 27939 33612 27988 33640
rect 27939 33609 27951 33612
rect 27893 33603 27951 33609
rect 27982 33600 27988 33612
rect 28040 33600 28046 33652
rect 30006 33600 30012 33652
rect 30064 33640 30070 33652
rect 30285 33643 30343 33649
rect 30285 33640 30297 33643
rect 30064 33612 30297 33640
rect 30064 33600 30070 33612
rect 30285 33609 30297 33612
rect 30331 33609 30343 33643
rect 30285 33603 30343 33609
rect 30745 33643 30803 33649
rect 30745 33609 30757 33643
rect 30791 33640 30803 33643
rect 31113 33643 31171 33649
rect 31113 33640 31125 33643
rect 30791 33612 31125 33640
rect 30791 33609 30803 33612
rect 30745 33603 30803 33609
rect 31113 33609 31125 33612
rect 31159 33609 31171 33643
rect 31113 33603 31171 33609
rect 31478 33600 31484 33652
rect 31536 33600 31542 33652
rect 31570 33600 31576 33652
rect 31628 33600 31634 33652
rect 33318 33600 33324 33652
rect 33376 33640 33382 33652
rect 33505 33643 33563 33649
rect 33505 33640 33517 33643
rect 33376 33612 33517 33640
rect 33376 33600 33382 33612
rect 33505 33609 33517 33612
rect 33551 33609 33563 33643
rect 33505 33603 33563 33609
rect 33873 33643 33931 33649
rect 33873 33609 33885 33643
rect 33919 33640 33931 33643
rect 34238 33640 34244 33652
rect 33919 33612 34244 33640
rect 33919 33609 33931 33612
rect 33873 33603 33931 33609
rect 34238 33600 34244 33612
rect 34296 33600 34302 33652
rect 34333 33643 34391 33649
rect 34333 33609 34345 33643
rect 34379 33640 34391 33643
rect 34422 33640 34428 33652
rect 34379 33612 34428 33640
rect 34379 33609 34391 33612
rect 34333 33603 34391 33609
rect 34422 33600 34428 33612
rect 34480 33600 34486 33652
rect 36262 33600 36268 33652
rect 36320 33640 36326 33652
rect 36357 33643 36415 33649
rect 36357 33640 36369 33643
rect 36320 33612 36369 33640
rect 36320 33600 36326 33612
rect 36357 33609 36369 33612
rect 36403 33609 36415 33643
rect 36357 33603 36415 33609
rect 37921 33643 37979 33649
rect 37921 33609 37933 33643
rect 37967 33640 37979 33643
rect 38102 33640 38108 33652
rect 37967 33612 38108 33640
rect 37967 33609 37979 33612
rect 37921 33603 37979 33609
rect 38102 33600 38108 33612
rect 38160 33600 38166 33652
rect 38749 33643 38807 33649
rect 38749 33609 38761 33643
rect 38795 33640 38807 33643
rect 39022 33640 39028 33652
rect 38795 33612 39028 33640
rect 38795 33609 38807 33612
rect 38749 33603 38807 33609
rect 39022 33600 39028 33612
rect 39080 33600 39086 33652
rect 41322 33600 41328 33652
rect 41380 33600 41386 33652
rect 41877 33643 41935 33649
rect 41877 33609 41889 33643
rect 41923 33640 41935 33643
rect 42150 33640 42156 33652
rect 41923 33612 42156 33640
rect 41923 33609 41935 33612
rect 41877 33603 41935 33609
rect 42150 33600 42156 33612
rect 42208 33600 42214 33652
rect 2317 33575 2375 33581
rect 2317 33541 2329 33575
rect 2363 33541 2375 33575
rect 2317 33535 2375 33541
rect 2777 33575 2835 33581
rect 2777 33541 2789 33575
rect 2823 33572 2835 33575
rect 3142 33572 3148 33584
rect 2823 33544 3148 33572
rect 2823 33541 2835 33544
rect 2777 33535 2835 33541
rect 3142 33532 3148 33544
rect 3200 33532 3206 33584
rect 3602 33532 3608 33584
rect 3660 33532 3666 33584
rect 5258 33572 5264 33584
rect 4908 33544 5264 33572
rect 1854 33464 1860 33516
rect 1912 33504 1918 33516
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1912 33476 2053 33504
rect 1912 33464 1918 33476
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 2056 33368 2084 33467
rect 2130 33464 2136 33516
rect 2188 33504 2194 33516
rect 4908 33513 4936 33544
rect 5258 33532 5264 33544
rect 5316 33532 5322 33584
rect 5813 33575 5871 33581
rect 5813 33541 5825 33575
rect 5859 33572 5871 33575
rect 5902 33572 5908 33584
rect 5859 33544 5908 33572
rect 5859 33541 5871 33544
rect 5813 33535 5871 33541
rect 5902 33532 5908 33544
rect 5960 33532 5966 33584
rect 7650 33532 7656 33584
rect 7708 33572 7714 33584
rect 8110 33572 8116 33584
rect 7708 33544 8116 33572
rect 7708 33532 7714 33544
rect 8110 33532 8116 33544
rect 8168 33532 8174 33584
rect 8294 33532 8300 33584
rect 8352 33572 8358 33584
rect 8389 33575 8447 33581
rect 8389 33572 8401 33575
rect 8352 33544 8401 33572
rect 8352 33532 8358 33544
rect 8389 33541 8401 33544
rect 8435 33572 8447 33575
rect 9582 33572 9588 33584
rect 8435 33544 9588 33572
rect 8435 33541 8447 33544
rect 8389 33535 8447 33541
rect 2593 33507 2651 33513
rect 2593 33504 2605 33507
rect 2188 33476 2605 33504
rect 2188 33464 2194 33476
rect 2593 33473 2605 33476
rect 2639 33473 2651 33507
rect 2593 33467 2651 33473
rect 2869 33507 2927 33513
rect 2869 33473 2881 33507
rect 2915 33473 2927 33507
rect 2869 33467 2927 33473
rect 4893 33507 4951 33513
rect 4893 33473 4905 33507
rect 4939 33473 4951 33507
rect 4893 33467 4951 33473
rect 2884 33368 2912 33467
rect 5350 33464 5356 33516
rect 5408 33464 5414 33516
rect 5442 33464 5448 33516
rect 5500 33464 5506 33516
rect 5534 33464 5540 33516
rect 5592 33504 5598 33516
rect 5629 33507 5687 33513
rect 5629 33504 5641 33507
rect 5592 33476 5641 33504
rect 5592 33464 5598 33476
rect 5629 33473 5641 33476
rect 5675 33473 5687 33507
rect 5629 33467 5687 33473
rect 8570 33464 8576 33516
rect 8628 33504 8634 33516
rect 9232 33513 9260 33544
rect 9582 33532 9588 33544
rect 9640 33532 9646 33584
rect 12161 33575 12219 33581
rect 12161 33541 12173 33575
rect 12207 33572 12219 33575
rect 13170 33572 13176 33584
rect 12207 33544 13176 33572
rect 12207 33541 12219 33544
rect 12161 33535 12219 33541
rect 13170 33532 13176 33544
rect 13228 33532 13234 33584
rect 8941 33507 8999 33513
rect 8941 33504 8953 33507
rect 8628 33476 8953 33504
rect 8628 33464 8634 33476
rect 8941 33473 8953 33476
rect 8987 33473 8999 33507
rect 8941 33467 8999 33473
rect 9217 33507 9275 33513
rect 9217 33473 9229 33507
rect 9263 33473 9275 33507
rect 9217 33467 9275 33473
rect 10594 33464 10600 33516
rect 10652 33464 10658 33516
rect 11057 33507 11115 33513
rect 11057 33473 11069 33507
rect 11103 33504 11115 33507
rect 11146 33504 11152 33516
rect 11103 33476 11152 33504
rect 11103 33473 11115 33476
rect 11057 33467 11115 33473
rect 11146 33464 11152 33476
rect 11204 33464 11210 33516
rect 11330 33464 11336 33516
rect 11388 33464 11394 33516
rect 11701 33507 11759 33513
rect 11701 33473 11713 33507
rect 11747 33504 11759 33507
rect 12434 33504 12440 33516
rect 11747 33476 12440 33504
rect 11747 33473 11759 33476
rect 11701 33467 11759 33473
rect 12434 33464 12440 33476
rect 12492 33464 12498 33516
rect 15933 33507 15991 33513
rect 15933 33473 15945 33507
rect 15979 33504 15991 33507
rect 16592 33504 16620 33600
rect 18616 33572 18644 33600
rect 18064 33544 18644 33572
rect 15979 33476 16620 33504
rect 15979 33473 15991 33476
rect 15933 33467 15991 33473
rect 17218 33464 17224 33516
rect 17276 33504 17282 33516
rect 18064 33513 18092 33544
rect 26234 33532 26240 33584
rect 26292 33572 26298 33584
rect 27246 33572 27252 33584
rect 26292 33544 27252 33572
rect 26292 33532 26298 33544
rect 27246 33532 27252 33544
rect 27304 33572 27310 33584
rect 27433 33575 27491 33581
rect 27433 33572 27445 33575
rect 27304 33544 27445 33572
rect 27304 33532 27310 33544
rect 27433 33541 27445 33544
rect 27479 33541 27491 33575
rect 27433 33535 27491 33541
rect 30653 33575 30711 33581
rect 30653 33541 30665 33575
rect 30699 33572 30711 33575
rect 31386 33572 31392 33584
rect 30699 33544 31392 33572
rect 30699 33541 30711 33544
rect 30653 33535 30711 33541
rect 31386 33532 31392 33544
rect 31444 33532 31450 33584
rect 32217 33575 32275 33581
rect 32217 33572 32229 33575
rect 31726 33544 32229 33572
rect 17782 33507 17840 33513
rect 17782 33504 17794 33507
rect 17276 33476 17794 33504
rect 17276 33464 17282 33476
rect 17782 33473 17794 33476
rect 17828 33473 17840 33507
rect 17782 33467 17840 33473
rect 18049 33507 18107 33513
rect 18049 33473 18061 33507
rect 18095 33473 18107 33507
rect 18049 33467 18107 33473
rect 18230 33464 18236 33516
rect 18288 33504 18294 33516
rect 18463 33507 18521 33513
rect 18463 33504 18475 33507
rect 18288 33476 18475 33504
rect 18288 33464 18294 33476
rect 18463 33473 18475 33476
rect 18509 33473 18521 33507
rect 18463 33467 18521 33473
rect 18601 33507 18659 33513
rect 18601 33473 18613 33507
rect 18647 33473 18659 33507
rect 18601 33467 18659 33473
rect 18693 33507 18751 33513
rect 18693 33473 18705 33507
rect 18739 33473 18751 33507
rect 18693 33467 18751 33473
rect 4614 33396 4620 33448
rect 4672 33396 4678 33448
rect 5166 33396 5172 33448
rect 5224 33396 5230 33448
rect 5258 33396 5264 33448
rect 5316 33396 5322 33448
rect 8662 33396 8668 33448
rect 8720 33396 8726 33448
rect 8849 33439 8907 33445
rect 8849 33405 8861 33439
rect 8895 33436 8907 33439
rect 9122 33436 9128 33448
rect 8895 33408 9128 33436
rect 8895 33405 8907 33408
rect 8849 33399 8907 33405
rect 9122 33396 9128 33408
rect 9180 33396 9186 33448
rect 9490 33396 9496 33448
rect 9548 33396 9554 33448
rect 10612 33436 10640 33464
rect 10612 33408 11192 33436
rect 2056 33340 2912 33368
rect 11054 33328 11060 33380
rect 11112 33328 11118 33380
rect 11164 33368 11192 33408
rect 11422 33396 11428 33448
rect 11480 33436 11486 33448
rect 11793 33439 11851 33445
rect 11793 33436 11805 33439
rect 11480 33408 11805 33436
rect 11480 33396 11486 33408
rect 11793 33405 11805 33408
rect 11839 33405 11851 33439
rect 11793 33399 11851 33405
rect 12342 33396 12348 33448
rect 12400 33396 12406 33448
rect 13078 33396 13084 33448
rect 13136 33396 13142 33448
rect 12710 33368 12716 33380
rect 11164 33340 12716 33368
rect 12710 33328 12716 33340
rect 12768 33328 12774 33380
rect 16485 33371 16543 33377
rect 16485 33337 16497 33371
rect 16531 33368 16543 33371
rect 16758 33368 16764 33380
rect 16531 33340 16764 33368
rect 16531 33337 16543 33340
rect 16485 33331 16543 33337
rect 16758 33328 16764 33340
rect 16816 33328 16822 33380
rect 18616 33368 18644 33467
rect 18708 33436 18736 33467
rect 18782 33464 18788 33516
rect 18840 33513 18846 33516
rect 18840 33507 18879 33513
rect 18867 33473 18879 33507
rect 18840 33467 18879 33473
rect 18840 33464 18846 33467
rect 18966 33464 18972 33516
rect 19024 33464 19030 33516
rect 19794 33464 19800 33516
rect 19852 33504 19858 33516
rect 20165 33507 20223 33513
rect 20165 33504 20177 33507
rect 19852 33476 20177 33504
rect 19852 33464 19858 33476
rect 20165 33473 20177 33476
rect 20211 33473 20223 33507
rect 20165 33467 20223 33473
rect 21358 33464 21364 33516
rect 21416 33504 21422 33516
rect 22373 33507 22431 33513
rect 22373 33504 22385 33507
rect 21416 33476 22385 33504
rect 21416 33464 21422 33476
rect 22373 33473 22385 33476
rect 22419 33473 22431 33507
rect 22373 33467 22431 33473
rect 23198 33464 23204 33516
rect 23256 33464 23262 33516
rect 23750 33464 23756 33516
rect 23808 33504 23814 33516
rect 24489 33507 24547 33513
rect 24489 33504 24501 33507
rect 23808 33476 24501 33504
rect 23808 33464 23814 33476
rect 24489 33473 24501 33476
rect 24535 33473 24547 33507
rect 24489 33467 24547 33473
rect 25133 33507 25191 33513
rect 25133 33473 25145 33507
rect 25179 33504 25191 33507
rect 25406 33504 25412 33516
rect 25179 33476 25412 33504
rect 25179 33473 25191 33476
rect 25133 33467 25191 33473
rect 25406 33464 25412 33476
rect 25464 33464 25470 33516
rect 26326 33464 26332 33516
rect 26384 33504 26390 33516
rect 26697 33507 26755 33513
rect 26697 33504 26709 33507
rect 26384 33476 26709 33504
rect 26384 33464 26390 33476
rect 26697 33473 26709 33476
rect 26743 33504 26755 33507
rect 27341 33507 27399 33513
rect 27341 33504 27353 33507
rect 26743 33476 27353 33504
rect 26743 33473 26755 33476
rect 26697 33467 26755 33473
rect 27341 33473 27353 33476
rect 27387 33473 27399 33507
rect 27341 33467 27399 33473
rect 28258 33464 28264 33516
rect 28316 33464 28322 33516
rect 28353 33507 28411 33513
rect 28353 33473 28365 33507
rect 28399 33504 28411 33507
rect 28718 33504 28724 33516
rect 28399 33476 28724 33504
rect 28399 33473 28411 33476
rect 28353 33467 28411 33473
rect 28718 33464 28724 33476
rect 28776 33464 28782 33516
rect 31726 33504 31754 33544
rect 32217 33541 32229 33544
rect 32263 33572 32275 33575
rect 36814 33572 36820 33584
rect 32263 33544 36820 33572
rect 32263 33541 32275 33544
rect 32217 33535 32275 33541
rect 36814 33532 36820 33544
rect 36872 33532 36878 33584
rect 39209 33575 39267 33581
rect 39209 33572 39221 33575
rect 38304 33544 39221 33572
rect 38304 33516 38332 33544
rect 39209 33541 39221 33544
rect 39255 33541 39267 33575
rect 39209 33535 39267 33541
rect 28828 33476 31754 33504
rect 20441 33439 20499 33445
rect 20441 33436 20453 33439
rect 18708 33408 20453 33436
rect 20441 33405 20453 33408
rect 20487 33436 20499 33439
rect 20714 33436 20720 33448
rect 20487 33408 20720 33436
rect 20487 33405 20499 33408
rect 20441 33399 20499 33405
rect 20714 33396 20720 33408
rect 20772 33396 20778 33448
rect 25222 33396 25228 33448
rect 25280 33396 25286 33448
rect 25314 33396 25320 33448
rect 25372 33436 25378 33448
rect 25958 33436 25964 33448
rect 25372 33408 25964 33436
rect 25372 33396 25378 33408
rect 25958 33396 25964 33408
rect 26016 33396 26022 33448
rect 26418 33396 26424 33448
rect 26476 33436 26482 33448
rect 27525 33439 27583 33445
rect 27525 33436 27537 33439
rect 26476 33408 27537 33436
rect 26476 33396 26482 33408
rect 27525 33405 27537 33408
rect 27571 33436 27583 33439
rect 28445 33439 28503 33445
rect 28445 33436 28457 33439
rect 27571 33408 28457 33436
rect 27571 33405 27583 33408
rect 27525 33399 27583 33405
rect 28445 33405 28457 33408
rect 28491 33436 28503 33439
rect 28828 33436 28856 33476
rect 33042 33464 33048 33516
rect 33100 33464 33106 33516
rect 33965 33507 34023 33513
rect 33965 33473 33977 33507
rect 34011 33504 34023 33507
rect 34146 33504 34152 33516
rect 34011 33476 34152 33504
rect 34011 33473 34023 33476
rect 33965 33467 34023 33473
rect 34146 33464 34152 33476
rect 34204 33504 34210 33516
rect 34701 33507 34759 33513
rect 34701 33504 34713 33507
rect 34204 33476 34713 33504
rect 34204 33464 34210 33476
rect 34701 33473 34713 33476
rect 34747 33473 34759 33507
rect 34701 33467 34759 33473
rect 38286 33464 38292 33516
rect 38344 33464 38350 33516
rect 38381 33507 38439 33513
rect 38381 33473 38393 33507
rect 38427 33504 38439 33507
rect 38654 33504 38660 33516
rect 38427 33476 38660 33504
rect 38427 33473 38439 33476
rect 38381 33467 38439 33473
rect 38654 33464 38660 33476
rect 38712 33504 38718 33516
rect 39117 33507 39175 33513
rect 39117 33504 39129 33507
rect 38712 33476 39129 33504
rect 38712 33464 38718 33476
rect 39117 33473 39129 33476
rect 39163 33473 39175 33507
rect 39117 33467 39175 33473
rect 39574 33464 39580 33516
rect 39632 33504 39638 33516
rect 40218 33513 40224 33516
rect 39945 33507 40003 33513
rect 39945 33504 39957 33507
rect 39632 33476 39957 33504
rect 39632 33464 39638 33476
rect 39945 33473 39957 33476
rect 39991 33473 40003 33507
rect 40212 33504 40224 33513
rect 40179 33476 40224 33504
rect 39945 33467 40003 33473
rect 40212 33467 40224 33476
rect 40218 33464 40224 33467
rect 40276 33464 40282 33516
rect 41598 33464 41604 33516
rect 41656 33504 41662 33516
rect 41785 33507 41843 33513
rect 41785 33504 41797 33507
rect 41656 33476 41797 33504
rect 41656 33464 41662 33476
rect 41785 33473 41797 33476
rect 41831 33473 41843 33507
rect 41785 33467 41843 33473
rect 28491 33408 28856 33436
rect 28491 33405 28503 33408
rect 28445 33399 28503 33405
rect 28902 33396 28908 33448
rect 28960 33436 28966 33448
rect 30837 33439 30895 33445
rect 30837 33436 30849 33439
rect 28960 33408 30849 33436
rect 28960 33396 28966 33408
rect 30837 33405 30849 33408
rect 30883 33405 30895 33439
rect 30837 33399 30895 33405
rect 20622 33368 20628 33380
rect 18616 33340 20628 33368
rect 20622 33328 20628 33340
rect 20680 33328 20686 33380
rect 30852 33368 30880 33399
rect 31662 33396 31668 33448
rect 31720 33436 31726 33448
rect 32493 33439 32551 33445
rect 32493 33436 32505 33439
rect 31720 33408 32505 33436
rect 31720 33396 31726 33408
rect 32493 33405 32505 33408
rect 32539 33436 32551 33439
rect 34057 33439 34115 33445
rect 34057 33436 34069 33439
rect 32539 33408 34069 33436
rect 32539 33405 32551 33408
rect 32493 33399 32551 33405
rect 34057 33405 34069 33408
rect 34103 33405 34115 33439
rect 34057 33399 34115 33405
rect 33226 33368 33232 33380
rect 30852 33340 33232 33368
rect 33226 33328 33232 33340
rect 33284 33328 33290 33380
rect 34072 33368 34100 33399
rect 34422 33396 34428 33448
rect 34480 33436 34486 33448
rect 34793 33439 34851 33445
rect 34793 33436 34805 33439
rect 34480 33408 34805 33436
rect 34480 33396 34486 33408
rect 34793 33405 34805 33408
rect 34839 33405 34851 33439
rect 34793 33399 34851 33405
rect 34977 33439 35035 33445
rect 34977 33405 34989 33439
rect 35023 33405 35035 33439
rect 34977 33399 35035 33405
rect 34992 33368 35020 33399
rect 36722 33396 36728 33448
rect 36780 33436 36786 33448
rect 36909 33439 36967 33445
rect 36909 33436 36921 33439
rect 36780 33408 36921 33436
rect 36780 33396 36786 33408
rect 36909 33405 36921 33408
rect 36955 33405 36967 33439
rect 36909 33399 36967 33405
rect 38565 33439 38623 33445
rect 38565 33405 38577 33439
rect 38611 33436 38623 33439
rect 39301 33439 39359 33445
rect 39301 33436 39313 33439
rect 38611 33408 39313 33436
rect 38611 33405 38623 33408
rect 38565 33399 38623 33405
rect 39301 33405 39313 33408
rect 39347 33405 39359 33439
rect 39301 33399 39359 33405
rect 38580 33368 38608 33399
rect 41966 33396 41972 33448
rect 42024 33396 42030 33448
rect 34072 33340 38608 33368
rect 40954 33328 40960 33380
rect 41012 33368 41018 33380
rect 41417 33371 41475 33377
rect 41417 33368 41429 33371
rect 41012 33340 41429 33368
rect 41012 33328 41018 33340
rect 41417 33337 41429 33340
rect 41463 33337 41475 33371
rect 41417 33331 41475 33337
rect 2222 33260 2228 33312
rect 2280 33300 2286 33312
rect 2317 33303 2375 33309
rect 2317 33300 2329 33303
rect 2280 33272 2329 33300
rect 2280 33260 2286 33272
rect 2317 33269 2329 33272
rect 2363 33269 2375 33303
rect 2317 33263 2375 33269
rect 2406 33260 2412 33312
rect 2464 33260 2470 33312
rect 3145 33303 3203 33309
rect 3145 33269 3157 33303
rect 3191 33300 3203 33303
rect 3326 33300 3332 33312
rect 3191 33272 3332 33300
rect 3191 33269 3203 33272
rect 3145 33263 3203 33269
rect 3326 33260 3332 33272
rect 3384 33260 3390 33312
rect 4982 33260 4988 33312
rect 5040 33260 5046 33312
rect 5810 33260 5816 33312
rect 5868 33300 5874 33312
rect 5997 33303 6055 33309
rect 5997 33300 6009 33303
rect 5868 33272 6009 33300
rect 5868 33260 5874 33272
rect 5997 33269 6009 33272
rect 6043 33269 6055 33303
rect 5997 33263 6055 33269
rect 8754 33260 8760 33312
rect 8812 33260 8818 33312
rect 10686 33260 10692 33312
rect 10744 33300 10750 33312
rect 10962 33300 10968 33312
rect 10744 33272 10968 33300
rect 10744 33260 10750 33272
rect 10962 33260 10968 33272
rect 11020 33260 11026 33312
rect 11514 33260 11520 33312
rect 11572 33260 11578 33312
rect 13630 33260 13636 33312
rect 13688 33260 13694 33312
rect 18138 33260 18144 33312
rect 18196 33300 18202 33312
rect 18325 33303 18383 33309
rect 18325 33300 18337 33303
rect 18196 33272 18337 33300
rect 18196 33260 18202 33272
rect 18325 33269 18337 33272
rect 18371 33269 18383 33303
rect 18325 33263 18383 33269
rect 26050 33260 26056 33312
rect 26108 33300 26114 33312
rect 26145 33303 26203 33309
rect 26145 33300 26157 33303
rect 26108 33272 26157 33300
rect 26108 33260 26114 33272
rect 26145 33269 26157 33272
rect 26191 33269 26203 33303
rect 26145 33263 26203 33269
rect 33321 33303 33379 33309
rect 33321 33269 33333 33303
rect 33367 33300 33379 33303
rect 34238 33300 34244 33312
rect 33367 33272 34244 33300
rect 33367 33269 33379 33272
rect 33321 33263 33379 33269
rect 34238 33260 34244 33272
rect 34296 33260 34302 33312
rect 1104 33210 42504 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 42504 33210
rect 1104 33136 42504 33158
rect 4614 33056 4620 33108
rect 4672 33096 4678 33108
rect 4709 33099 4767 33105
rect 4709 33096 4721 33099
rect 4672 33068 4721 33096
rect 4672 33056 4678 33068
rect 4709 33065 4721 33068
rect 4755 33065 4767 33099
rect 4709 33059 4767 33065
rect 4985 33099 5043 33105
rect 4985 33065 4997 33099
rect 5031 33096 5043 33099
rect 5074 33096 5080 33108
rect 5031 33068 5080 33096
rect 5031 33065 5043 33068
rect 4985 33059 5043 33065
rect 5074 33056 5080 33068
rect 5132 33056 5138 33108
rect 5442 33056 5448 33108
rect 5500 33096 5506 33108
rect 5537 33099 5595 33105
rect 5537 33096 5549 33099
rect 5500 33068 5549 33096
rect 5500 33056 5506 33068
rect 5537 33065 5549 33068
rect 5583 33096 5595 33099
rect 6546 33096 6552 33108
rect 5583 33068 6552 33096
rect 5583 33065 5595 33068
rect 5537 33059 5595 33065
rect 6546 33056 6552 33068
rect 6604 33056 6610 33108
rect 7006 33056 7012 33108
rect 7064 33096 7070 33108
rect 7561 33099 7619 33105
rect 7561 33096 7573 33099
rect 7064 33068 7573 33096
rect 7064 33056 7070 33068
rect 7561 33065 7573 33068
rect 7607 33065 7619 33099
rect 7561 33059 7619 33065
rect 9490 33056 9496 33108
rect 9548 33056 9554 33108
rect 9582 33056 9588 33108
rect 9640 33096 9646 33108
rect 9640 33068 11008 33096
rect 9640 33056 9646 33068
rect 3421 33031 3479 33037
rect 3421 32997 3433 33031
rect 3467 33028 3479 33031
rect 4798 33028 4804 33040
rect 3467 33000 4804 33028
rect 3467 32997 3479 33000
rect 3421 32991 3479 32997
rect 4798 32988 4804 33000
rect 4856 32988 4862 33040
rect 5721 33031 5779 33037
rect 5721 32997 5733 33031
rect 5767 33028 5779 33031
rect 5902 33028 5908 33040
rect 5767 33000 5908 33028
rect 5767 32997 5779 33000
rect 5721 32991 5779 32997
rect 2774 32920 2780 32972
rect 2832 32960 2838 32972
rect 3145 32963 3203 32969
rect 3145 32960 3157 32963
rect 2832 32932 3157 32960
rect 2832 32920 2838 32932
rect 3145 32929 3157 32932
rect 3191 32929 3203 32963
rect 3145 32923 3203 32929
rect 3605 32963 3663 32969
rect 3605 32929 3617 32963
rect 3651 32960 3663 32963
rect 4982 32960 4988 32972
rect 3651 32932 4988 32960
rect 3651 32929 3663 32932
rect 3605 32923 3663 32929
rect 4982 32920 4988 32932
rect 5040 32920 5046 32972
rect 5350 32960 5356 32972
rect 5092 32932 5356 32960
rect 3326 32852 3332 32904
rect 3384 32852 3390 32904
rect 4433 32895 4491 32901
rect 4433 32892 4445 32895
rect 3620 32864 4445 32892
rect 2314 32784 2320 32836
rect 2372 32784 2378 32836
rect 2866 32784 2872 32836
rect 2924 32784 2930 32836
rect 1397 32759 1455 32765
rect 1397 32725 1409 32759
rect 1443 32756 1455 32759
rect 2130 32756 2136 32768
rect 1443 32728 2136 32756
rect 1443 32725 1455 32728
rect 1397 32719 1455 32725
rect 2130 32716 2136 32728
rect 2188 32756 2194 32768
rect 2498 32756 2504 32768
rect 2188 32728 2504 32756
rect 2188 32716 2194 32728
rect 2498 32716 2504 32728
rect 2556 32716 2562 32768
rect 3344 32756 3372 32852
rect 3620 32833 3648 32864
rect 4433 32861 4445 32864
rect 4479 32861 4491 32895
rect 4433 32855 4491 32861
rect 4525 32895 4583 32901
rect 4525 32861 4537 32895
rect 4571 32861 4583 32895
rect 4525 32855 4583 32861
rect 3605 32827 3663 32833
rect 3605 32793 3617 32827
rect 3651 32793 3663 32827
rect 3605 32787 3663 32793
rect 4065 32827 4123 32833
rect 4065 32793 4077 32827
rect 4111 32793 4123 32827
rect 4065 32787 4123 32793
rect 4080 32756 4108 32787
rect 4154 32784 4160 32836
rect 4212 32784 4218 32836
rect 4540 32768 4568 32855
rect 4706 32852 4712 32904
rect 4764 32892 4770 32904
rect 5092 32892 5120 32932
rect 5350 32920 5356 32932
rect 5408 32920 5414 32972
rect 5736 32960 5764 32991
rect 5902 32988 5908 33000
rect 5960 32988 5966 33040
rect 10781 33031 10839 33037
rect 10781 33028 10793 33031
rect 9784 33000 10793 33028
rect 5460 32932 5764 32960
rect 7469 32963 7527 32969
rect 4764 32864 5120 32892
rect 5166 32895 5224 32901
rect 4764 32852 4770 32864
rect 5166 32861 5178 32895
rect 5212 32892 5224 32895
rect 5460 32892 5488 32932
rect 7469 32929 7481 32963
rect 7515 32960 7527 32963
rect 8294 32960 8300 32972
rect 7515 32932 8300 32960
rect 7515 32929 7527 32932
rect 7469 32923 7527 32929
rect 8294 32920 8300 32932
rect 8352 32920 8358 32972
rect 5212 32864 5488 32892
rect 5212 32861 5224 32864
rect 5166 32855 5224 32861
rect 5626 32852 5632 32904
rect 5684 32852 5690 32904
rect 7742 32852 7748 32904
rect 7800 32852 7806 32904
rect 7837 32895 7895 32901
rect 7837 32861 7849 32895
rect 7883 32892 7895 32895
rect 8754 32892 8760 32904
rect 7883 32864 8760 32892
rect 7883 32861 7895 32864
rect 7837 32855 7895 32861
rect 8754 32852 8760 32864
rect 8812 32852 8818 32904
rect 9784 32901 9812 33000
rect 10781 32997 10793 33000
rect 10827 32997 10839 33031
rect 10781 32991 10839 32997
rect 10226 32960 10232 32972
rect 9876 32932 10232 32960
rect 9876 32901 9904 32932
rect 10226 32920 10232 32932
rect 10284 32920 10290 32972
rect 10980 32969 11008 33068
rect 12342 33056 12348 33108
rect 12400 33056 12406 33108
rect 12437 33099 12495 33105
rect 12437 33065 12449 33099
rect 12483 33096 12495 33099
rect 13078 33096 13084 33108
rect 12483 33068 13084 33096
rect 12483 33065 12495 33068
rect 12437 33059 12495 33065
rect 13078 33056 13084 33068
rect 13136 33096 13142 33108
rect 13136 33068 14403 33096
rect 13136 33056 13142 33068
rect 10965 32963 11023 32969
rect 10965 32929 10977 32963
rect 11011 32929 11023 32963
rect 10965 32923 11023 32929
rect 14185 32963 14243 32969
rect 14185 32929 14197 32963
rect 14231 32929 14243 32963
rect 14185 32923 14243 32929
rect 9677 32895 9735 32901
rect 9677 32861 9689 32895
rect 9723 32861 9735 32895
rect 9677 32855 9735 32861
rect 9769 32895 9827 32901
rect 9769 32861 9781 32895
rect 9815 32861 9827 32895
rect 9769 32855 9827 32861
rect 9861 32895 9919 32901
rect 9861 32861 9873 32895
rect 9907 32861 9919 32895
rect 9861 32855 9919 32861
rect 5074 32784 5080 32836
rect 5132 32824 5138 32836
rect 5442 32824 5448 32836
rect 5132 32796 5448 32824
rect 5132 32784 5138 32796
rect 5442 32784 5448 32796
rect 5500 32784 5506 32836
rect 5902 32784 5908 32836
rect 5960 32824 5966 32836
rect 5960 32796 6026 32824
rect 5960 32784 5966 32796
rect 7190 32784 7196 32836
rect 7248 32784 7254 32836
rect 8110 32784 8116 32836
rect 8168 32784 8174 32836
rect 8205 32827 8263 32833
rect 8205 32793 8217 32827
rect 8251 32824 8263 32827
rect 8938 32824 8944 32836
rect 8251 32796 8944 32824
rect 8251 32793 8263 32796
rect 8205 32787 8263 32793
rect 8938 32784 8944 32796
rect 8996 32784 9002 32836
rect 4430 32756 4436 32768
rect 3344 32728 4436 32756
rect 4430 32716 4436 32728
rect 4488 32716 4494 32768
rect 4522 32716 4528 32768
rect 4580 32756 4586 32768
rect 5169 32759 5227 32765
rect 5169 32756 5181 32759
rect 4580 32728 5181 32756
rect 4580 32716 4586 32728
rect 5169 32725 5181 32728
rect 5215 32756 5227 32759
rect 5534 32756 5540 32768
rect 5215 32728 5540 32756
rect 5215 32725 5227 32728
rect 5169 32719 5227 32725
rect 5534 32716 5540 32728
rect 5592 32716 5598 32768
rect 9692 32756 9720 32855
rect 9950 32852 9956 32904
rect 10008 32901 10014 32904
rect 10008 32895 10037 32901
rect 10025 32861 10037 32895
rect 10008 32855 10037 32861
rect 10008 32852 10014 32855
rect 10134 32852 10140 32904
rect 10192 32852 10198 32904
rect 10413 32895 10471 32901
rect 10413 32861 10425 32895
rect 10459 32892 10471 32895
rect 10686 32892 10692 32904
rect 10459 32864 10692 32892
rect 10459 32861 10471 32864
rect 10413 32855 10471 32861
rect 10686 32852 10692 32864
rect 10744 32852 10750 32904
rect 10873 32895 10931 32901
rect 10873 32861 10885 32895
rect 10919 32861 10931 32895
rect 10873 32855 10931 32861
rect 11232 32895 11290 32901
rect 11232 32861 11244 32895
rect 11278 32892 11290 32895
rect 11514 32892 11520 32904
rect 11278 32864 11520 32892
rect 11278 32861 11290 32864
rect 11232 32855 11290 32861
rect 10594 32784 10600 32836
rect 10652 32824 10658 32836
rect 10888 32824 10916 32855
rect 11514 32852 11520 32864
rect 11572 32852 11578 32904
rect 13814 32852 13820 32904
rect 13872 32852 13878 32904
rect 11330 32824 11336 32836
rect 10652 32796 11336 32824
rect 10652 32784 10658 32796
rect 11330 32784 11336 32796
rect 11388 32784 11394 32836
rect 13572 32827 13630 32833
rect 13572 32793 13584 32827
rect 13618 32824 13630 32827
rect 13906 32824 13912 32836
rect 13618 32796 13912 32824
rect 13618 32793 13630 32796
rect 13572 32787 13630 32793
rect 13906 32784 13912 32796
rect 13964 32784 13970 32836
rect 10229 32759 10287 32765
rect 10229 32756 10241 32759
rect 9692 32728 10241 32756
rect 10229 32725 10241 32728
rect 10275 32725 10287 32759
rect 14200 32756 14228 32923
rect 14277 32895 14335 32901
rect 14277 32861 14289 32895
rect 14323 32861 14335 32895
rect 14375 32892 14403 33068
rect 17218 33056 17224 33108
rect 17276 33056 17282 33108
rect 18417 33099 18475 33105
rect 18417 33065 18429 33099
rect 18463 33096 18475 33099
rect 18782 33096 18788 33108
rect 18463 33068 18788 33096
rect 18463 33065 18475 33068
rect 18417 33059 18475 33065
rect 18782 33056 18788 33068
rect 18840 33056 18846 33108
rect 20898 33056 20904 33108
rect 20956 33096 20962 33108
rect 21085 33099 21143 33105
rect 21085 33096 21097 33099
rect 20956 33068 21097 33096
rect 20956 33056 20962 33068
rect 21085 33065 21097 33068
rect 21131 33096 21143 33099
rect 21266 33096 21272 33108
rect 21131 33068 21272 33096
rect 21131 33065 21143 33068
rect 21085 33059 21143 33065
rect 21266 33056 21272 33068
rect 21324 33056 21330 33108
rect 22738 33056 22744 33108
rect 22796 33096 22802 33108
rect 22925 33099 22983 33105
rect 22925 33096 22937 33099
rect 22796 33068 22937 33096
rect 22796 33056 22802 33068
rect 22925 33065 22937 33068
rect 22971 33096 22983 33099
rect 23106 33096 23112 33108
rect 22971 33068 23112 33096
rect 22971 33065 22983 33068
rect 22925 33059 22983 33065
rect 23106 33056 23112 33068
rect 23164 33056 23170 33108
rect 24581 33099 24639 33105
rect 24581 33065 24593 33099
rect 24627 33096 24639 33099
rect 25222 33096 25228 33108
rect 24627 33068 25228 33096
rect 24627 33065 24639 33068
rect 24581 33059 24639 33065
rect 25222 33056 25228 33068
rect 25280 33056 25286 33108
rect 26326 33056 26332 33108
rect 26384 33096 26390 33108
rect 26697 33099 26755 33105
rect 26697 33096 26709 33099
rect 26384 33068 26709 33096
rect 26384 33056 26390 33068
rect 26697 33065 26709 33068
rect 26743 33065 26755 33099
rect 26697 33059 26755 33065
rect 38286 33056 38292 33108
rect 38344 33096 38350 33108
rect 38473 33099 38531 33105
rect 38473 33096 38485 33099
rect 38344 33068 38485 33096
rect 38344 33056 38350 33068
rect 38473 33065 38485 33068
rect 38519 33065 38531 33099
rect 38473 33059 38531 33065
rect 14645 33031 14703 33037
rect 14645 32997 14657 33031
rect 14691 33028 14703 33031
rect 15289 33031 15347 33037
rect 14691 33000 14872 33028
rect 14691 32997 14703 33000
rect 14645 32991 14703 32997
rect 14844 32969 14872 33000
rect 15289 32997 15301 33031
rect 15335 33028 15347 33031
rect 15654 33028 15660 33040
rect 15335 33000 15660 33028
rect 15335 32997 15347 33000
rect 15289 32991 15347 32997
rect 15654 32988 15660 33000
rect 15712 32988 15718 33040
rect 17034 33028 17040 33040
rect 16684 33000 17040 33028
rect 14829 32963 14887 32969
rect 14829 32929 14841 32963
rect 14875 32929 14887 32963
rect 14829 32923 14887 32929
rect 15473 32963 15531 32969
rect 15473 32929 15485 32963
rect 15519 32960 15531 32963
rect 15838 32960 15844 32972
rect 15519 32932 15844 32960
rect 15519 32929 15531 32932
rect 15473 32923 15531 32929
rect 14921 32895 14979 32901
rect 14921 32892 14933 32895
rect 14375 32864 14933 32892
rect 14277 32855 14335 32861
rect 14921 32861 14933 32864
rect 14967 32861 14979 32895
rect 14921 32855 14979 32861
rect 14292 32824 14320 32855
rect 15470 32824 15476 32836
rect 14292 32796 15476 32824
rect 15470 32784 15476 32796
rect 15528 32784 15534 32836
rect 15194 32756 15200 32768
rect 14200 32728 15200 32756
rect 10229 32719 10287 32725
rect 15194 32716 15200 32728
rect 15252 32756 15258 32768
rect 15580 32756 15608 32932
rect 15838 32920 15844 32932
rect 15896 32920 15902 32972
rect 16574 32920 16580 32972
rect 16632 32960 16638 32972
rect 16684 32969 16712 33000
rect 17034 32988 17040 33000
rect 17092 32988 17098 33040
rect 23014 33028 23020 33040
rect 22572 33000 23020 33028
rect 16669 32963 16727 32969
rect 16669 32960 16681 32963
rect 16632 32932 16681 32960
rect 16632 32920 16638 32932
rect 16669 32929 16681 32932
rect 16715 32929 16727 32963
rect 16669 32923 16727 32929
rect 16758 32920 16764 32972
rect 16816 32920 16822 32972
rect 19337 32963 19395 32969
rect 19337 32960 19349 32963
rect 17788 32932 19349 32960
rect 17788 32901 17816 32932
rect 19337 32929 19349 32932
rect 19383 32960 19395 32963
rect 19610 32960 19616 32972
rect 19383 32932 19616 32960
rect 19383 32929 19395 32932
rect 19337 32923 19395 32929
rect 19610 32920 19616 32932
rect 19668 32960 19674 32972
rect 21177 32963 21235 32969
rect 21177 32960 21189 32963
rect 19668 32932 21189 32960
rect 19668 32920 19674 32932
rect 21177 32929 21189 32932
rect 21223 32929 21235 32963
rect 21177 32923 21235 32929
rect 17773 32895 17831 32901
rect 17773 32861 17785 32895
rect 17819 32892 17831 32895
rect 17862 32892 17868 32904
rect 17819 32864 17868 32892
rect 17819 32861 17831 32864
rect 17773 32855 17831 32861
rect 17862 32852 17868 32864
rect 17920 32852 17926 32904
rect 19061 32895 19119 32901
rect 19061 32861 19073 32895
rect 19107 32861 19119 32895
rect 22572 32878 22600 33000
rect 23014 32988 23020 33000
rect 23072 32988 23078 33040
rect 28258 32988 28264 33040
rect 28316 33028 28322 33040
rect 28537 33031 28595 33037
rect 28537 33028 28549 33031
rect 28316 33000 28549 33028
rect 28316 32988 28322 33000
rect 28537 32997 28549 33000
rect 28583 32997 28595 33031
rect 28537 32991 28595 32997
rect 32493 33031 32551 33037
rect 32493 32997 32505 33031
rect 32539 32997 32551 33031
rect 32493 32991 32551 32997
rect 24394 32920 24400 32972
rect 24452 32960 24458 32972
rect 28552 32960 28580 32991
rect 29181 32963 29239 32969
rect 29181 32960 29193 32963
rect 24452 32932 25360 32960
rect 28552 32932 29193 32960
rect 24452 32920 24458 32932
rect 23017 32895 23075 32901
rect 19061 32855 19119 32861
rect 23017 32861 23029 32895
rect 23063 32861 23075 32895
rect 23017 32855 23075 32861
rect 19076 32824 19104 32855
rect 19518 32824 19524 32836
rect 19076 32796 19524 32824
rect 19518 32784 19524 32796
rect 19576 32784 19582 32836
rect 19613 32827 19671 32833
rect 19613 32793 19625 32827
rect 19659 32793 19671 32827
rect 19613 32787 19671 32793
rect 15252 32728 15608 32756
rect 15252 32716 15258 32728
rect 16022 32716 16028 32768
rect 16080 32716 16086 32768
rect 16853 32759 16911 32765
rect 16853 32725 16865 32759
rect 16899 32756 16911 32759
rect 17770 32756 17776 32768
rect 16899 32728 17776 32756
rect 16899 32725 16911 32728
rect 16853 32719 16911 32725
rect 17770 32716 17776 32728
rect 17828 32716 17834 32768
rect 19628 32756 19656 32787
rect 20070 32784 20076 32836
rect 20128 32784 20134 32836
rect 21358 32824 21364 32836
rect 21008 32796 21364 32824
rect 21008 32756 21036 32796
rect 21358 32784 21364 32796
rect 21416 32784 21422 32836
rect 21450 32784 21456 32836
rect 21508 32784 21514 32836
rect 23032 32824 23060 32855
rect 25130 32852 25136 32904
rect 25188 32852 25194 32904
rect 25332 32901 25360 32932
rect 29181 32929 29193 32932
rect 29227 32929 29239 32963
rect 29181 32923 29239 32929
rect 29730 32920 29736 32972
rect 29788 32960 29794 32972
rect 31113 32963 31171 32969
rect 31113 32960 31125 32963
rect 29788 32932 31125 32960
rect 29788 32920 29794 32932
rect 31113 32929 31125 32932
rect 31159 32929 31171 32963
rect 32508 32960 32536 32991
rect 33229 32963 33287 32969
rect 33229 32960 33241 32963
rect 32508 32932 33241 32960
rect 31113 32923 31171 32929
rect 33229 32929 33241 32932
rect 33275 32960 33287 32963
rect 33594 32960 33600 32972
rect 33275 32932 33600 32960
rect 33275 32929 33287 32932
rect 33229 32923 33287 32929
rect 33594 32920 33600 32932
rect 33652 32920 33658 32972
rect 33962 32920 33968 32972
rect 34020 32960 34026 32972
rect 34238 32960 34244 32972
rect 34020 32932 34244 32960
rect 34020 32920 34026 32932
rect 34238 32920 34244 32932
rect 34296 32960 34302 32972
rect 35529 32963 35587 32969
rect 35529 32960 35541 32963
rect 34296 32932 35541 32960
rect 34296 32920 34302 32932
rect 35529 32929 35541 32932
rect 35575 32929 35587 32963
rect 38488 32960 38516 33059
rect 41230 33056 41236 33108
rect 41288 33096 41294 33108
rect 41693 33099 41751 33105
rect 41693 33096 41705 33099
rect 41288 33068 41705 33096
rect 41288 33056 41294 33068
rect 41693 33065 41705 33068
rect 41739 33065 41751 33099
rect 41693 33059 41751 33065
rect 39117 32963 39175 32969
rect 39117 32960 39129 32963
rect 38488 32932 39129 32960
rect 35529 32923 35587 32929
rect 39117 32929 39129 32932
rect 39163 32929 39175 32963
rect 39117 32923 39175 32929
rect 25317 32895 25375 32901
rect 25317 32861 25329 32895
rect 25363 32892 25375 32895
rect 27062 32892 27068 32904
rect 25363 32864 27068 32892
rect 25363 32861 25375 32864
rect 25317 32855 25375 32861
rect 27062 32852 27068 32864
rect 27120 32892 27126 32904
rect 27157 32895 27215 32901
rect 27157 32892 27169 32895
rect 27120 32864 27169 32892
rect 27120 32852 27126 32864
rect 27157 32861 27169 32864
rect 27203 32861 27215 32895
rect 27157 32855 27215 32861
rect 30650 32852 30656 32904
rect 30708 32852 30714 32904
rect 34698 32852 34704 32904
rect 34756 32892 34762 32904
rect 35434 32892 35440 32904
rect 34756 32864 35440 32892
rect 34756 32852 34762 32864
rect 35434 32852 35440 32864
rect 35492 32892 35498 32904
rect 36357 32895 36415 32901
rect 36357 32892 36369 32895
rect 35492 32864 36369 32892
rect 35492 32852 35498 32864
rect 36357 32861 36369 32864
rect 36403 32861 36415 32895
rect 36357 32855 36415 32861
rect 37093 32895 37151 32901
rect 37093 32861 37105 32895
rect 37139 32892 37151 32895
rect 37182 32892 37188 32904
rect 37139 32864 37188 32892
rect 37139 32861 37151 32864
rect 37093 32855 37151 32861
rect 37182 32852 37188 32864
rect 37240 32852 37246 32904
rect 39666 32852 39672 32904
rect 39724 32892 39730 32904
rect 40313 32895 40371 32901
rect 40313 32892 40325 32895
rect 39724 32864 40325 32892
rect 39724 32852 39730 32864
rect 40313 32861 40325 32864
rect 40359 32861 40371 32895
rect 40313 32855 40371 32861
rect 40580 32895 40638 32901
rect 40580 32861 40592 32895
rect 40626 32892 40638 32895
rect 40954 32892 40960 32904
rect 40626 32864 40960 32892
rect 40626 32861 40638 32864
rect 40580 32855 40638 32861
rect 40954 32852 40960 32864
rect 41012 32852 41018 32904
rect 22756 32796 23060 32824
rect 25584 32827 25642 32833
rect 19628 32728 21036 32756
rect 21726 32716 21732 32768
rect 21784 32756 21790 32768
rect 22756 32756 22784 32796
rect 25584 32793 25596 32827
rect 25630 32824 25642 32827
rect 25774 32824 25780 32836
rect 25630 32796 25780 32824
rect 25630 32793 25642 32796
rect 25584 32787 25642 32793
rect 25774 32784 25780 32796
rect 25832 32784 25838 32836
rect 27430 32833 27436 32836
rect 27424 32787 27436 32833
rect 27430 32784 27436 32787
rect 27488 32784 27494 32836
rect 28074 32784 28080 32836
rect 28132 32824 28138 32836
rect 28629 32827 28687 32833
rect 28629 32824 28641 32827
rect 28132 32796 28641 32824
rect 28132 32784 28138 32796
rect 28629 32793 28641 32796
rect 28675 32793 28687 32827
rect 28629 32787 28687 32793
rect 31380 32827 31438 32833
rect 31380 32793 31392 32827
rect 31426 32824 31438 32827
rect 32030 32824 32036 32836
rect 31426 32796 32036 32824
rect 31426 32793 31438 32796
rect 31380 32787 31438 32793
rect 32030 32784 32036 32796
rect 32088 32784 32094 32836
rect 34057 32827 34115 32833
rect 34057 32793 34069 32827
rect 34103 32824 34115 32827
rect 34330 32824 34336 32836
rect 34103 32796 34336 32824
rect 34103 32793 34115 32796
rect 34057 32787 34115 32793
rect 34330 32784 34336 32796
rect 34388 32784 34394 32836
rect 34606 32784 34612 32836
rect 34664 32824 34670 32836
rect 35345 32827 35403 32833
rect 35345 32824 35357 32827
rect 34664 32796 35357 32824
rect 34664 32784 34670 32796
rect 35345 32793 35357 32796
rect 35391 32793 35403 32827
rect 35345 32787 35403 32793
rect 37360 32827 37418 32833
rect 37360 32793 37372 32827
rect 37406 32824 37418 32827
rect 38102 32824 38108 32836
rect 37406 32796 38108 32824
rect 37406 32793 37418 32796
rect 37360 32787 37418 32793
rect 38102 32784 38108 32796
rect 38160 32784 38166 32836
rect 21784 32728 22784 32756
rect 23201 32759 23259 32765
rect 21784 32716 21790 32728
rect 23201 32725 23213 32759
rect 23247 32756 23259 32759
rect 23658 32756 23664 32768
rect 23247 32728 23664 32756
rect 23247 32725 23259 32728
rect 23201 32719 23259 32725
rect 23658 32716 23664 32728
rect 23716 32716 23722 32768
rect 30098 32716 30104 32768
rect 30156 32716 30162 32768
rect 32582 32716 32588 32768
rect 32640 32716 32646 32768
rect 33686 32716 33692 32768
rect 33744 32716 33750 32768
rect 34149 32759 34207 32765
rect 34149 32725 34161 32759
rect 34195 32756 34207 32759
rect 34882 32756 34888 32768
rect 34195 32728 34888 32756
rect 34195 32725 34207 32728
rect 34149 32719 34207 32725
rect 34882 32716 34888 32728
rect 34940 32716 34946 32768
rect 34974 32716 34980 32768
rect 35032 32716 35038 32768
rect 35437 32759 35495 32765
rect 35437 32725 35449 32759
rect 35483 32756 35495 32759
rect 35805 32759 35863 32765
rect 35805 32756 35817 32759
rect 35483 32728 35817 32756
rect 35483 32725 35495 32728
rect 35437 32719 35495 32725
rect 35805 32725 35817 32728
rect 35851 32725 35863 32759
rect 35805 32719 35863 32725
rect 38562 32716 38568 32768
rect 38620 32716 38626 32768
rect 1104 32666 42504 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 42504 32666
rect 1104 32592 42504 32614
rect 2777 32555 2835 32561
rect 2777 32521 2789 32555
rect 2823 32552 2835 32555
rect 2866 32552 2872 32564
rect 2823 32524 2872 32552
rect 2823 32521 2835 32524
rect 2777 32515 2835 32521
rect 2866 32512 2872 32524
rect 2924 32512 2930 32564
rect 3234 32512 3240 32564
rect 3292 32512 3298 32564
rect 4417 32555 4475 32561
rect 4417 32521 4429 32555
rect 4463 32552 4475 32555
rect 4522 32552 4528 32564
rect 4463 32524 4528 32552
rect 4463 32521 4475 32524
rect 4417 32515 4475 32521
rect 4522 32512 4528 32524
rect 4580 32512 4586 32564
rect 4982 32552 4988 32564
rect 4632 32524 4988 32552
rect 2406 32444 2412 32496
rect 2464 32444 2470 32496
rect 4632 32493 4660 32524
rect 4982 32512 4988 32524
rect 5040 32512 5046 32564
rect 5810 32552 5816 32564
rect 5644 32524 5816 32552
rect 4617 32487 4675 32493
rect 4617 32453 4629 32487
rect 4663 32453 4675 32487
rect 5350 32484 5356 32496
rect 4617 32447 4675 32453
rect 4708 32456 5356 32484
rect 2222 32376 2228 32428
rect 2280 32376 2286 32428
rect 2498 32376 2504 32428
rect 2556 32376 2562 32428
rect 2593 32419 2651 32425
rect 2593 32385 2605 32419
rect 2639 32385 2651 32419
rect 2593 32379 2651 32385
rect 2608 32280 2636 32379
rect 3142 32376 3148 32428
rect 3200 32376 3206 32428
rect 3418 32376 3424 32428
rect 3476 32416 3482 32428
rect 3513 32419 3571 32425
rect 3513 32416 3525 32419
rect 3476 32388 3525 32416
rect 3476 32376 3482 32388
rect 3513 32385 3525 32388
rect 3559 32416 3571 32419
rect 4708 32416 4736 32456
rect 5350 32444 5356 32456
rect 5408 32444 5414 32496
rect 5644 32493 5672 32524
rect 5810 32512 5816 32524
rect 5868 32512 5874 32564
rect 5997 32555 6055 32561
rect 5997 32521 6009 32555
rect 6043 32552 6055 32555
rect 7190 32552 7196 32564
rect 6043 32524 7196 32552
rect 6043 32521 6055 32524
rect 5997 32515 6055 32521
rect 7190 32512 7196 32524
rect 7248 32512 7254 32564
rect 8021 32555 8079 32561
rect 8021 32521 8033 32555
rect 8067 32552 8079 32555
rect 8110 32552 8116 32564
rect 8067 32524 8116 32552
rect 8067 32521 8079 32524
rect 8021 32515 8079 32521
rect 8110 32512 8116 32524
rect 8168 32552 8174 32564
rect 9950 32552 9956 32564
rect 8168 32524 9956 32552
rect 8168 32512 8174 32524
rect 9950 32512 9956 32524
rect 10008 32512 10014 32564
rect 21910 32552 21916 32564
rect 12084 32524 21916 32552
rect 12084 32493 12112 32524
rect 21910 32512 21916 32524
rect 21968 32552 21974 32564
rect 32122 32552 32128 32564
rect 21968 32524 32128 32552
rect 21968 32512 21974 32524
rect 32122 32512 32128 32524
rect 32180 32512 32186 32564
rect 34146 32512 34152 32564
rect 34204 32512 34210 32564
rect 34790 32512 34796 32564
rect 34848 32512 34854 32564
rect 34882 32512 34888 32564
rect 34940 32552 34946 32564
rect 35989 32555 36047 32561
rect 35989 32552 36001 32555
rect 34940 32524 36001 32552
rect 34940 32512 34946 32524
rect 35989 32521 36001 32524
rect 36035 32521 36047 32555
rect 35989 32515 36047 32521
rect 38654 32512 38660 32564
rect 38712 32512 38718 32564
rect 40862 32512 40868 32564
rect 40920 32552 40926 32564
rect 41049 32555 41107 32561
rect 41049 32552 41061 32555
rect 40920 32524 41061 32552
rect 40920 32512 40926 32524
rect 41049 32521 41061 32524
rect 41095 32552 41107 32555
rect 41095 32524 41736 32552
rect 41095 32521 41107 32524
rect 41049 32515 41107 32521
rect 5629 32487 5687 32493
rect 5629 32453 5641 32487
rect 5675 32453 5687 32487
rect 5629 32447 5687 32453
rect 12069 32487 12127 32493
rect 12069 32453 12081 32487
rect 12115 32453 12127 32487
rect 12069 32447 12127 32453
rect 12158 32444 12164 32496
rect 12216 32484 12222 32496
rect 13725 32487 13783 32493
rect 13725 32484 13737 32487
rect 12216 32456 13737 32484
rect 12216 32444 12222 32456
rect 13725 32453 13737 32456
rect 13771 32484 13783 32487
rect 16850 32484 16856 32496
rect 13771 32456 16856 32484
rect 13771 32453 13783 32456
rect 13725 32447 13783 32453
rect 16850 32444 16856 32456
rect 16908 32444 16914 32496
rect 18138 32444 18144 32496
rect 18196 32444 18202 32496
rect 20070 32484 20076 32496
rect 19366 32470 20076 32484
rect 19352 32456 20076 32470
rect 3559 32388 4736 32416
rect 3559 32385 3571 32388
rect 3513 32379 3571 32385
rect 4798 32376 4804 32428
rect 4856 32416 4862 32428
rect 4893 32419 4951 32425
rect 4893 32416 4905 32419
rect 4856 32388 4905 32416
rect 4856 32376 4862 32388
rect 4893 32385 4905 32388
rect 4939 32385 4951 32419
rect 4893 32379 4951 32385
rect 4982 32376 4988 32428
rect 5040 32376 5046 32428
rect 5442 32376 5448 32428
rect 5500 32376 5506 32428
rect 5721 32419 5779 32425
rect 5721 32385 5733 32419
rect 5767 32385 5779 32419
rect 5721 32379 5779 32385
rect 5813 32419 5871 32425
rect 5813 32385 5825 32419
rect 5859 32416 5871 32419
rect 6270 32416 6276 32428
rect 5859 32388 6276 32416
rect 5859 32385 5871 32388
rect 5813 32379 5871 32385
rect 3694 32308 3700 32360
rect 3752 32308 3758 32360
rect 4706 32308 4712 32360
rect 4764 32348 4770 32360
rect 5074 32348 5080 32360
rect 4764 32320 5080 32348
rect 4764 32308 4770 32320
rect 5074 32308 5080 32320
rect 5132 32308 5138 32360
rect 5169 32351 5227 32357
rect 5169 32317 5181 32351
rect 5215 32317 5227 32351
rect 5169 32311 5227 32317
rect 5736 32348 5764 32379
rect 6270 32376 6276 32388
rect 6328 32376 6334 32428
rect 6365 32419 6423 32425
rect 6365 32385 6377 32419
rect 6411 32385 6423 32419
rect 6365 32379 6423 32385
rect 5994 32348 6000 32360
rect 5736 32320 6000 32348
rect 3326 32280 3332 32292
rect 2608 32252 3332 32280
rect 3326 32240 3332 32252
rect 3384 32240 3390 32292
rect 5184 32280 5212 32311
rect 5534 32280 5540 32292
rect 4448 32252 5540 32280
rect 4062 32172 4068 32224
rect 4120 32212 4126 32224
rect 4448 32221 4476 32252
rect 5534 32240 5540 32252
rect 5592 32240 5598 32292
rect 4249 32215 4307 32221
rect 4249 32212 4261 32215
rect 4120 32184 4261 32212
rect 4120 32172 4126 32184
rect 4249 32181 4261 32184
rect 4295 32181 4307 32215
rect 4249 32175 4307 32181
rect 4433 32215 4491 32221
rect 4433 32181 4445 32215
rect 4479 32181 4491 32215
rect 4433 32175 4491 32181
rect 4706 32172 4712 32224
rect 4764 32172 4770 32224
rect 4982 32172 4988 32224
rect 5040 32212 5046 32224
rect 5258 32212 5264 32224
rect 5040 32184 5264 32212
rect 5040 32172 5046 32184
rect 5258 32172 5264 32184
rect 5316 32212 5322 32224
rect 5736 32212 5764 32320
rect 5994 32308 6000 32320
rect 6052 32308 6058 32360
rect 6086 32308 6092 32360
rect 6144 32348 6150 32360
rect 6380 32348 6408 32379
rect 6454 32376 6460 32428
rect 6512 32416 6518 32428
rect 7929 32419 7987 32425
rect 7929 32416 7941 32419
rect 6512 32388 7941 32416
rect 6512 32376 6518 32388
rect 7929 32385 7941 32388
rect 7975 32385 7987 32419
rect 7929 32379 7987 32385
rect 9858 32376 9864 32428
rect 9916 32416 9922 32428
rect 10137 32419 10195 32425
rect 10137 32416 10149 32419
rect 9916 32388 10149 32416
rect 9916 32376 9922 32388
rect 10137 32385 10149 32388
rect 10183 32416 10195 32419
rect 10594 32416 10600 32428
rect 10183 32388 10600 32416
rect 10183 32385 10195 32388
rect 10137 32379 10195 32385
rect 10594 32376 10600 32388
rect 10652 32376 10658 32428
rect 13906 32376 13912 32428
rect 13964 32376 13970 32428
rect 15562 32376 15568 32428
rect 15620 32416 15626 32428
rect 15850 32419 15908 32425
rect 15850 32416 15862 32419
rect 15620 32388 15862 32416
rect 15620 32376 15626 32388
rect 15850 32385 15862 32388
rect 15896 32385 15908 32419
rect 15850 32379 15908 32385
rect 16117 32419 16175 32425
rect 16117 32385 16129 32419
rect 16163 32416 16175 32419
rect 16390 32416 16396 32428
rect 16163 32388 16396 32416
rect 16163 32385 16175 32388
rect 16117 32379 16175 32385
rect 16390 32376 16396 32388
rect 16448 32416 16454 32428
rect 17681 32419 17739 32425
rect 17681 32416 17693 32419
rect 16448 32388 17693 32416
rect 16448 32376 16454 32388
rect 17681 32385 17693 32388
rect 17727 32416 17739 32419
rect 17862 32416 17868 32428
rect 17727 32388 17868 32416
rect 17727 32385 17739 32388
rect 17681 32379 17739 32385
rect 17862 32376 17868 32388
rect 17920 32376 17926 32428
rect 8662 32348 8668 32360
rect 6144 32320 8668 32348
rect 6144 32308 6150 32320
rect 8662 32308 8668 32320
rect 8720 32308 8726 32360
rect 14458 32308 14464 32360
rect 14516 32308 14522 32360
rect 18598 32308 18604 32360
rect 18656 32348 18662 32360
rect 19352 32348 19380 32456
rect 20070 32444 20076 32456
rect 20128 32444 20134 32496
rect 20622 32444 20628 32496
rect 20680 32444 20686 32496
rect 20806 32444 20812 32496
rect 20864 32484 20870 32496
rect 21177 32487 21235 32493
rect 21177 32484 21189 32487
rect 20864 32456 21189 32484
rect 20864 32444 20870 32456
rect 21177 32453 21189 32456
rect 21223 32453 21235 32487
rect 21177 32447 21235 32453
rect 21358 32444 21364 32496
rect 21416 32444 21422 32496
rect 22189 32487 22247 32493
rect 22189 32453 22201 32487
rect 22235 32484 22247 32487
rect 22370 32484 22376 32496
rect 22235 32456 22376 32484
rect 22235 32453 22247 32456
rect 22189 32447 22247 32453
rect 22370 32444 22376 32456
rect 22428 32444 22434 32496
rect 23014 32444 23020 32496
rect 23072 32444 23078 32496
rect 24026 32444 24032 32496
rect 24084 32484 24090 32496
rect 24397 32487 24455 32493
rect 24397 32484 24409 32487
rect 24084 32456 24409 32484
rect 24084 32444 24090 32456
rect 24397 32453 24409 32456
rect 24443 32453 24455 32487
rect 24397 32447 24455 32453
rect 26050 32444 26056 32496
rect 26108 32484 26114 32496
rect 26237 32487 26295 32493
rect 26237 32484 26249 32487
rect 26108 32456 26249 32484
rect 26108 32444 26114 32456
rect 26237 32453 26249 32456
rect 26283 32453 26295 32487
rect 26237 32447 26295 32453
rect 26326 32444 26332 32496
rect 26384 32444 26390 32496
rect 28810 32484 28816 32496
rect 28460 32456 28816 32484
rect 20530 32376 20536 32428
rect 20588 32376 20594 32428
rect 20714 32376 20720 32428
rect 20772 32376 20778 32428
rect 20898 32376 20904 32428
rect 20956 32376 20962 32428
rect 20993 32419 21051 32425
rect 20993 32385 21005 32419
rect 21039 32385 21051 32419
rect 20993 32379 21051 32385
rect 18656 32320 19380 32348
rect 19613 32351 19671 32357
rect 18656 32308 18662 32320
rect 19613 32317 19625 32351
rect 19659 32348 19671 32351
rect 19702 32348 19708 32360
rect 19659 32320 19708 32348
rect 19659 32317 19671 32320
rect 19613 32311 19671 32317
rect 19702 32308 19708 32320
rect 19760 32308 19766 32360
rect 21008 32348 21036 32379
rect 21818 32376 21824 32428
rect 21876 32416 21882 32428
rect 22051 32419 22109 32425
rect 22051 32416 22063 32419
rect 21876 32388 22063 32416
rect 21876 32376 21882 32388
rect 22051 32385 22063 32388
rect 22097 32385 22109 32419
rect 22051 32379 22109 32385
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32385 22339 32419
rect 22281 32379 22339 32385
rect 22465 32419 22523 32425
rect 22465 32385 22477 32419
rect 22511 32416 22523 32419
rect 22738 32416 22744 32428
rect 22511 32388 22744 32416
rect 22511 32385 22523 32388
rect 22465 32379 22523 32385
rect 20364 32320 21036 32348
rect 22296 32348 22324 32379
rect 22738 32376 22744 32388
rect 22796 32376 22802 32428
rect 24302 32376 24308 32428
rect 24360 32376 24366 32428
rect 24578 32376 24584 32428
rect 24636 32376 24642 32428
rect 25590 32376 25596 32428
rect 25648 32376 25654 32428
rect 26145 32419 26203 32425
rect 26145 32385 26157 32419
rect 26191 32416 26203 32419
rect 26344 32416 26372 32444
rect 26191 32388 26372 32416
rect 26191 32385 26203 32388
rect 26145 32379 26203 32385
rect 27154 32376 27160 32428
rect 27212 32416 27218 32428
rect 27985 32419 28043 32425
rect 27985 32416 27997 32419
rect 27212 32388 27997 32416
rect 27212 32376 27218 32388
rect 27985 32385 27997 32388
rect 28031 32385 28043 32419
rect 27985 32379 28043 32385
rect 28074 32376 28080 32428
rect 28132 32376 28138 32428
rect 28460 32425 28488 32456
rect 28810 32444 28816 32456
rect 28868 32484 28874 32496
rect 29730 32484 29736 32496
rect 28868 32456 29736 32484
rect 28868 32444 28874 32456
rect 29730 32444 29736 32456
rect 29788 32444 29794 32496
rect 30098 32444 30104 32496
rect 30156 32484 30162 32496
rect 30377 32487 30435 32493
rect 30377 32484 30389 32487
rect 30156 32456 30389 32484
rect 30156 32444 30162 32456
rect 30377 32453 30389 32456
rect 30423 32453 30435 32487
rect 34808 32484 34836 32512
rect 30377 32447 30435 32453
rect 34532 32456 34836 32484
rect 28445 32419 28503 32425
rect 28445 32385 28457 32419
rect 28491 32385 28503 32419
rect 28445 32379 28503 32385
rect 28712 32419 28770 32425
rect 28712 32385 28724 32419
rect 28758 32416 28770 32419
rect 28758 32388 29960 32416
rect 28758 32385 28770 32388
rect 28712 32379 28770 32385
rect 23658 32348 23664 32360
rect 22296 32320 23664 32348
rect 6546 32240 6552 32292
rect 6604 32240 6610 32292
rect 13170 32240 13176 32292
rect 13228 32280 13234 32292
rect 20364 32289 20392 32320
rect 20349 32283 20407 32289
rect 13228 32252 15240 32280
rect 13228 32240 13234 32252
rect 5316 32184 5764 32212
rect 5316 32172 5322 32184
rect 9582 32172 9588 32224
rect 9640 32212 9646 32224
rect 10045 32215 10103 32221
rect 10045 32212 10057 32215
rect 9640 32184 10057 32212
rect 9640 32172 9646 32184
rect 10045 32181 10057 32184
rect 10091 32181 10103 32215
rect 10045 32175 10103 32181
rect 14737 32215 14795 32221
rect 14737 32181 14749 32215
rect 14783 32212 14795 32215
rect 15102 32212 15108 32224
rect 14783 32184 15108 32212
rect 14783 32181 14795 32184
rect 14737 32175 14795 32181
rect 15102 32172 15108 32184
rect 15160 32172 15166 32224
rect 15212 32212 15240 32252
rect 20349 32249 20361 32283
rect 20395 32249 20407 32283
rect 20349 32243 20407 32249
rect 20714 32240 20720 32292
rect 20772 32280 20778 32292
rect 22296 32280 22324 32320
rect 23658 32308 23664 32320
rect 23716 32308 23722 32360
rect 24029 32351 24087 32357
rect 24029 32317 24041 32351
rect 24075 32348 24087 32351
rect 24765 32351 24823 32357
rect 24765 32348 24777 32351
rect 24075 32320 24777 32348
rect 24075 32317 24087 32320
rect 24029 32311 24087 32317
rect 24765 32317 24777 32320
rect 24811 32317 24823 32351
rect 24765 32311 24823 32317
rect 26050 32308 26056 32360
rect 26108 32348 26114 32360
rect 26329 32351 26387 32357
rect 26329 32348 26341 32351
rect 26108 32320 26341 32348
rect 26108 32308 26114 32320
rect 26329 32317 26341 32320
rect 26375 32317 26387 32351
rect 26329 32311 26387 32317
rect 28261 32351 28319 32357
rect 28261 32317 28273 32351
rect 28307 32317 28319 32351
rect 28261 32311 28319 32317
rect 20772 32252 22324 32280
rect 20772 32240 20778 32252
rect 25774 32240 25780 32292
rect 25832 32240 25838 32292
rect 27430 32240 27436 32292
rect 27488 32280 27494 32292
rect 27617 32283 27675 32289
rect 27617 32280 27629 32283
rect 27488 32252 27629 32280
rect 27488 32240 27494 32252
rect 27617 32249 27629 32252
rect 27663 32249 27675 32283
rect 27617 32243 27675 32249
rect 16114 32212 16120 32224
rect 15212 32184 16120 32212
rect 16114 32172 16120 32184
rect 16172 32172 16178 32224
rect 21913 32215 21971 32221
rect 21913 32181 21925 32215
rect 21959 32212 21971 32215
rect 22002 32212 22008 32224
rect 21959 32184 22008 32212
rect 21959 32181 21971 32184
rect 21913 32175 21971 32181
rect 22002 32172 22008 32184
rect 22060 32172 22066 32224
rect 22554 32172 22560 32224
rect 22612 32172 22618 32224
rect 25038 32172 25044 32224
rect 25096 32172 25102 32224
rect 28276 32212 28304 32311
rect 29932 32289 29960 32388
rect 30190 32376 30196 32428
rect 30248 32416 30254 32428
rect 30285 32419 30343 32425
rect 30285 32416 30297 32419
rect 30248 32388 30297 32416
rect 30248 32376 30254 32388
rect 30285 32385 30297 32388
rect 30331 32385 30343 32419
rect 30285 32379 30343 32385
rect 31478 32376 31484 32428
rect 31536 32416 31542 32428
rect 31573 32419 31631 32425
rect 31573 32416 31585 32419
rect 31536 32388 31585 32416
rect 31536 32376 31542 32388
rect 31573 32385 31585 32388
rect 31619 32385 31631 32419
rect 31573 32379 31631 32385
rect 33036 32419 33094 32425
rect 33036 32385 33048 32419
rect 33082 32416 33094 32419
rect 33318 32416 33324 32428
rect 33082 32388 33324 32416
rect 33082 32385 33094 32388
rect 33036 32379 33094 32385
rect 33318 32376 33324 32388
rect 33376 32376 33382 32428
rect 34532 32425 34560 32456
rect 34974 32444 34980 32496
rect 35032 32444 35038 32496
rect 34517 32419 34575 32425
rect 34517 32385 34529 32419
rect 34563 32385 34575 32419
rect 34517 32379 34575 32385
rect 34784 32419 34842 32425
rect 34784 32385 34796 32419
rect 34830 32416 34842 32419
rect 34992 32416 35020 32444
rect 34830 32388 35020 32416
rect 34830 32385 34842 32388
rect 34784 32379 34842 32385
rect 37366 32376 37372 32428
rect 37424 32416 37430 32428
rect 37533 32419 37591 32425
rect 37533 32416 37545 32419
rect 37424 32388 37545 32416
rect 37424 32376 37430 32388
rect 37533 32385 37545 32388
rect 37579 32385 37591 32419
rect 38672 32416 38700 32512
rect 39301 32419 39359 32425
rect 39301 32416 39313 32419
rect 38672 32388 39313 32416
rect 37533 32379 37591 32385
rect 39301 32385 39313 32388
rect 39347 32385 39359 32419
rect 39301 32379 39359 32385
rect 39666 32376 39672 32428
rect 39724 32376 39730 32428
rect 39942 32425 39948 32428
rect 39936 32379 39948 32425
rect 39942 32376 39948 32379
rect 40000 32376 40006 32428
rect 41708 32425 41736 32524
rect 41693 32419 41751 32425
rect 41693 32385 41705 32419
rect 41739 32385 41751 32419
rect 41693 32379 41751 32385
rect 41877 32419 41935 32425
rect 41877 32385 41889 32419
rect 41923 32416 41935 32419
rect 42150 32416 42156 32428
rect 41923 32388 42156 32416
rect 41923 32385 41935 32388
rect 41877 32379 41935 32385
rect 42150 32376 42156 32388
rect 42208 32376 42214 32428
rect 30469 32351 30527 32357
rect 30469 32348 30481 32351
rect 30300 32320 30481 32348
rect 30300 32292 30328 32320
rect 30469 32317 30481 32320
rect 30515 32317 30527 32351
rect 30469 32311 30527 32317
rect 32766 32308 32772 32360
rect 32824 32308 32830 32360
rect 36541 32351 36599 32357
rect 36541 32317 36553 32351
rect 36587 32317 36599 32351
rect 36541 32311 36599 32317
rect 29917 32283 29975 32289
rect 29917 32249 29929 32283
rect 29963 32249 29975 32283
rect 29917 32243 29975 32249
rect 30282 32240 30288 32292
rect 30340 32240 30346 32292
rect 36556 32280 36584 32311
rect 37274 32308 37280 32360
rect 37332 32308 37338 32360
rect 35452 32252 36584 32280
rect 29178 32212 29184 32224
rect 28276 32184 29184 32212
rect 29178 32172 29184 32184
rect 29236 32172 29242 32224
rect 29825 32215 29883 32221
rect 29825 32181 29837 32215
rect 29871 32212 29883 32215
rect 30650 32212 30656 32224
rect 29871 32184 30656 32212
rect 29871 32181 29883 32184
rect 29825 32175 29883 32181
rect 30650 32172 30656 32184
rect 30708 32172 30714 32224
rect 31018 32172 31024 32224
rect 31076 32172 31082 32224
rect 34422 32172 34428 32224
rect 34480 32212 34486 32224
rect 35452 32212 35480 32252
rect 34480 32184 35480 32212
rect 34480 32172 34486 32184
rect 35526 32172 35532 32224
rect 35584 32212 35590 32224
rect 35897 32215 35955 32221
rect 35897 32212 35909 32215
rect 35584 32184 35909 32212
rect 35584 32172 35590 32184
rect 35897 32181 35909 32184
rect 35943 32181 35955 32215
rect 37292 32212 37320 32308
rect 37918 32212 37924 32224
rect 37292 32184 37924 32212
rect 35897 32175 35955 32181
rect 37918 32172 37924 32184
rect 37976 32172 37982 32224
rect 38746 32172 38752 32224
rect 38804 32172 38810 32224
rect 41138 32172 41144 32224
rect 41196 32172 41202 32224
rect 42058 32172 42064 32224
rect 42116 32172 42122 32224
rect 1104 32122 42504 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 42504 32122
rect 1104 32048 42504 32070
rect 4614 31968 4620 32020
rect 4672 31968 4678 32020
rect 5166 32008 5172 32020
rect 4724 31980 5172 32008
rect 3694 31900 3700 31952
rect 3752 31940 3758 31952
rect 4724 31940 4752 31980
rect 5166 31968 5172 31980
rect 5224 31968 5230 32020
rect 5350 31968 5356 32020
rect 5408 32008 5414 32020
rect 5445 32011 5503 32017
rect 5445 32008 5457 32011
rect 5408 31980 5457 32008
rect 5408 31968 5414 31980
rect 5445 31977 5457 31980
rect 5491 31977 5503 32011
rect 5445 31971 5503 31977
rect 5626 31968 5632 32020
rect 5684 31968 5690 32020
rect 7650 31968 7656 32020
rect 7708 32008 7714 32020
rect 11514 32008 11520 32020
rect 7708 31980 11520 32008
rect 7708 31968 7714 31980
rect 11514 31968 11520 31980
rect 11572 31968 11578 32020
rect 13817 32011 13875 32017
rect 13817 31977 13829 32011
rect 13863 32008 13875 32011
rect 14458 32008 14464 32020
rect 13863 31980 14464 32008
rect 13863 31977 13875 31980
rect 13817 31971 13875 31977
rect 14458 31968 14464 31980
rect 14516 31968 14522 32020
rect 15470 31968 15476 32020
rect 15528 31968 15534 32020
rect 15562 31968 15568 32020
rect 15620 31968 15626 32020
rect 16390 32008 16396 32020
rect 16040 31980 16396 32008
rect 3752 31912 4752 31940
rect 8128 31912 9260 31940
rect 3752 31900 3758 31912
rect 3326 31832 3332 31884
rect 3384 31872 3390 31884
rect 3970 31872 3976 31884
rect 3384 31844 3976 31872
rect 3384 31832 3390 31844
rect 3970 31832 3976 31844
rect 4028 31872 4034 31884
rect 6270 31872 6276 31884
rect 4028 31844 6276 31872
rect 4028 31832 4034 31844
rect 6270 31832 6276 31844
rect 6328 31832 6334 31884
rect 2866 31764 2872 31816
rect 2924 31804 2930 31816
rect 3237 31807 3295 31813
rect 3237 31804 3249 31807
rect 2924 31776 3249 31804
rect 2924 31764 2930 31776
rect 3237 31773 3249 31776
rect 3283 31773 3295 31807
rect 3237 31767 3295 31773
rect 4798 31764 4804 31816
rect 4856 31764 4862 31816
rect 4985 31807 5043 31813
rect 4985 31773 4997 31807
rect 5031 31804 5043 31807
rect 5074 31804 5080 31816
rect 5031 31776 5080 31804
rect 5031 31773 5043 31776
rect 4985 31767 5043 31773
rect 5074 31764 5080 31776
rect 5132 31764 5138 31816
rect 5350 31764 5356 31816
rect 5408 31804 5414 31816
rect 6454 31804 6460 31816
rect 5408 31776 6460 31804
rect 5408 31764 5414 31776
rect 6454 31764 6460 31776
rect 6512 31764 6518 31816
rect 6638 31764 6644 31816
rect 6696 31804 6702 31816
rect 6733 31807 6791 31813
rect 6733 31804 6745 31807
rect 6696 31776 6745 31804
rect 6696 31764 6702 31776
rect 6733 31773 6745 31776
rect 6779 31773 6791 31807
rect 8128 31790 8156 31912
rect 8294 31832 8300 31884
rect 8352 31872 8358 31884
rect 9125 31875 9183 31881
rect 9125 31872 9137 31875
rect 8352 31844 9137 31872
rect 8352 31832 8358 31844
rect 9125 31841 9137 31844
rect 9171 31841 9183 31875
rect 9232 31872 9260 31912
rect 9232 31844 10548 31872
rect 9125 31835 9183 31841
rect 10520 31816 10548 31844
rect 13170 31832 13176 31884
rect 13228 31832 13234 31884
rect 13357 31875 13415 31881
rect 13357 31841 13369 31875
rect 13403 31872 13415 31875
rect 13630 31872 13636 31884
rect 13403 31844 13636 31872
rect 13403 31841 13415 31844
rect 13357 31835 13415 31841
rect 13630 31832 13636 31844
rect 13688 31832 13694 31884
rect 16040 31872 16068 31980
rect 16390 31968 16396 31980
rect 16448 31968 16454 32020
rect 17770 31968 17776 32020
rect 17828 32008 17834 32020
rect 18141 32011 18199 32017
rect 18141 32008 18153 32011
rect 17828 31980 18153 32008
rect 17828 31968 17834 31980
rect 18141 31977 18153 31980
rect 18187 31977 18199 32011
rect 18141 31971 18199 31977
rect 19981 32011 20039 32017
rect 19981 31977 19993 32011
rect 20027 32008 20039 32011
rect 20346 32008 20352 32020
rect 20027 31980 20352 32008
rect 20027 31977 20039 31980
rect 19981 31971 20039 31977
rect 20346 31968 20352 31980
rect 20404 32008 20410 32020
rect 20530 32008 20536 32020
rect 20404 31980 20536 32008
rect 20404 31968 20410 31980
rect 20530 31968 20536 31980
rect 20588 31968 20594 32020
rect 21450 31968 21456 32020
rect 21508 32008 21514 32020
rect 22281 32011 22339 32017
rect 22281 32008 22293 32011
rect 21508 31980 22293 32008
rect 21508 31968 21514 31980
rect 22281 31977 22293 31980
rect 22327 31977 22339 32011
rect 22281 31971 22339 31977
rect 22554 31968 22560 32020
rect 22612 32008 22618 32020
rect 23474 32008 23480 32020
rect 22612 31980 23480 32008
rect 22612 31968 22618 31980
rect 23474 31968 23480 31980
rect 23532 31968 23538 32020
rect 24026 31968 24032 32020
rect 24084 31968 24090 32020
rect 24412 31980 25360 32008
rect 21542 31900 21548 31952
rect 21600 31940 21606 31952
rect 24412 31940 24440 31980
rect 21600 31912 24440 31940
rect 25332 31940 25360 31980
rect 25590 31968 25596 32020
rect 25648 32008 25654 32020
rect 25777 32011 25835 32017
rect 25777 32008 25789 32011
rect 25648 31980 25789 32008
rect 25648 31968 25654 31980
rect 25777 31977 25789 31980
rect 25823 31977 25835 32011
rect 25777 31971 25835 31977
rect 25884 31980 26832 32008
rect 25884 31940 25912 31980
rect 25332 31912 25912 31940
rect 26804 31940 26832 31980
rect 27246 31968 27252 32020
rect 27304 31968 27310 32020
rect 31113 32011 31171 32017
rect 27356 31980 28948 32008
rect 27356 31940 27384 31980
rect 26804 31912 27384 31940
rect 21600 31900 21606 31912
rect 28718 31900 28724 31952
rect 28776 31900 28782 31952
rect 15948 31844 16068 31872
rect 16209 31875 16267 31881
rect 6733 31767 6791 31773
rect 10502 31764 10508 31816
rect 10560 31764 10566 31816
rect 11517 31807 11575 31813
rect 11517 31804 11529 31807
rect 10888 31776 11529 31804
rect 5258 31696 5264 31748
rect 5316 31696 5322 31748
rect 7006 31696 7012 31748
rect 7064 31696 7070 31748
rect 9398 31696 9404 31748
rect 9456 31696 9462 31748
rect 10888 31680 10916 31776
rect 11517 31773 11529 31776
rect 11563 31773 11575 31807
rect 11517 31767 11575 31773
rect 11606 31764 11612 31816
rect 11664 31804 11670 31816
rect 12069 31807 12127 31813
rect 12069 31804 12081 31807
rect 11664 31776 12081 31804
rect 11664 31764 11670 31776
rect 12069 31773 12081 31776
rect 12115 31804 12127 31807
rect 12158 31804 12164 31816
rect 12115 31776 12164 31804
rect 12115 31773 12127 31776
rect 12069 31767 12127 31773
rect 12158 31764 12164 31776
rect 12216 31764 12222 31816
rect 13814 31764 13820 31816
rect 13872 31804 13878 31816
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13872 31776 14105 31804
rect 13872 31764 13878 31776
rect 14093 31773 14105 31776
rect 14139 31804 14151 31807
rect 15948 31804 15976 31844
rect 16209 31841 16221 31875
rect 16255 31841 16267 31875
rect 16209 31835 16267 31841
rect 14139 31776 15976 31804
rect 14139 31773 14151 31776
rect 14093 31767 14151 31773
rect 16022 31764 16028 31816
rect 16080 31764 16086 31816
rect 16114 31764 16120 31816
rect 16172 31804 16178 31816
rect 16224 31804 16252 31835
rect 16390 31832 16396 31884
rect 16448 31832 16454 31884
rect 19429 31875 19487 31881
rect 19429 31841 19441 31875
rect 19475 31872 19487 31875
rect 19702 31872 19708 31884
rect 19475 31844 19708 31872
rect 19475 31841 19487 31844
rect 19429 31835 19487 31841
rect 19702 31832 19708 31844
rect 19760 31832 19766 31884
rect 20622 31832 20628 31884
rect 20680 31872 20686 31884
rect 22370 31872 22376 31884
rect 20680 31844 22376 31872
rect 20680 31832 20686 31844
rect 22370 31832 22376 31844
rect 22428 31872 22434 31884
rect 22738 31872 22744 31884
rect 22428 31844 22744 31872
rect 22428 31832 22434 31844
rect 22738 31832 22744 31844
rect 22796 31832 22802 31884
rect 16172 31776 16252 31804
rect 21913 31807 21971 31813
rect 16172 31764 16178 31776
rect 21913 31773 21925 31807
rect 21959 31804 21971 31807
rect 22002 31804 22008 31816
rect 21959 31776 22008 31804
rect 21959 31773 21971 31776
rect 21913 31767 21971 31773
rect 22002 31764 22008 31776
rect 22060 31764 22066 31816
rect 22756 31804 22784 31832
rect 22756 31776 23428 31804
rect 14360 31739 14418 31745
rect 14360 31705 14372 31739
rect 14406 31736 14418 31739
rect 14458 31736 14464 31748
rect 14406 31708 14464 31736
rect 14406 31705 14418 31708
rect 14360 31699 14418 31705
rect 14458 31696 14464 31708
rect 14516 31696 14522 31748
rect 16132 31736 16160 31764
rect 16574 31736 16580 31748
rect 16132 31708 16580 31736
rect 16574 31696 16580 31708
rect 16632 31696 16638 31748
rect 16666 31696 16672 31748
rect 16724 31696 16730 31748
rect 18138 31736 18144 31748
rect 17894 31708 18144 31736
rect 18138 31696 18144 31708
rect 18196 31736 18202 31748
rect 18598 31736 18604 31748
rect 18196 31708 18604 31736
rect 18196 31696 18202 31708
rect 18598 31696 18604 31708
rect 18656 31696 18662 31748
rect 19334 31696 19340 31748
rect 19392 31736 19398 31748
rect 19613 31739 19671 31745
rect 19613 31736 19625 31739
rect 19392 31708 19625 31736
rect 19392 31696 19398 31708
rect 19613 31705 19625 31708
rect 19659 31705 19671 31739
rect 19613 31699 19671 31705
rect 22094 31696 22100 31748
rect 22152 31696 22158 31748
rect 23400 31736 23428 31776
rect 23474 31764 23480 31816
rect 23532 31764 23538 31816
rect 23658 31764 23664 31816
rect 23716 31764 23722 31816
rect 23761 31807 23819 31813
rect 23761 31773 23773 31807
rect 23807 31773 23819 31807
rect 23869 31807 23927 31813
rect 23869 31804 23881 31807
rect 23761 31767 23819 31773
rect 23860 31773 23881 31804
rect 23915 31773 23927 31807
rect 23860 31767 23927 31773
rect 24397 31807 24455 31813
rect 24397 31773 24409 31807
rect 24443 31804 24455 31807
rect 25774 31804 25780 31816
rect 24443 31776 25780 31804
rect 24443 31773 24455 31776
rect 24397 31767 24455 31773
rect 23768 31736 23796 31767
rect 23400 31708 23796 31736
rect 23860 31736 23888 31767
rect 25774 31764 25780 31776
rect 25832 31804 25838 31816
rect 25869 31807 25927 31813
rect 25869 31804 25881 31807
rect 25832 31776 25881 31804
rect 25832 31764 25838 31776
rect 25869 31773 25881 31776
rect 25915 31804 25927 31807
rect 27062 31804 27068 31816
rect 25915 31776 27068 31804
rect 25915 31773 25927 31776
rect 25869 31767 25927 31773
rect 27062 31764 27068 31776
rect 27120 31804 27126 31816
rect 27341 31807 27399 31813
rect 27341 31804 27353 31807
rect 27120 31776 27353 31804
rect 27120 31764 27126 31776
rect 27341 31773 27353 31776
rect 27387 31804 27399 31807
rect 28810 31804 28816 31816
rect 27387 31776 28816 31804
rect 27387 31773 27399 31776
rect 27341 31767 27399 31773
rect 28810 31764 28816 31776
rect 28868 31764 28874 31816
rect 24026 31736 24032 31748
rect 23860 31708 24032 31736
rect 24026 31696 24032 31708
rect 24084 31696 24090 31748
rect 24664 31739 24722 31745
rect 24664 31705 24676 31739
rect 24710 31736 24722 31739
rect 24854 31736 24860 31748
rect 24710 31708 24860 31736
rect 24710 31705 24722 31708
rect 24664 31699 24722 31705
rect 24854 31696 24860 31708
rect 24912 31696 24918 31748
rect 26142 31745 26148 31748
rect 26136 31699 26148 31745
rect 26142 31696 26148 31699
rect 26200 31696 26206 31748
rect 27608 31739 27666 31745
rect 27608 31705 27620 31739
rect 27654 31736 27666 31739
rect 27706 31736 27712 31748
rect 27654 31708 27712 31736
rect 27654 31705 27666 31708
rect 27608 31699 27666 31705
rect 27706 31696 27712 31708
rect 27764 31696 27770 31748
rect 28920 31745 28948 31980
rect 31113 31977 31125 32011
rect 31159 32008 31171 32011
rect 31478 32008 31484 32020
rect 31159 31980 31484 32008
rect 31159 31977 31171 31980
rect 31113 31971 31171 31977
rect 31478 31968 31484 31980
rect 31536 31968 31542 32020
rect 33962 31968 33968 32020
rect 34020 31968 34026 32020
rect 34422 31968 34428 32020
rect 34480 31968 34486 32020
rect 37277 32011 37335 32017
rect 37277 31977 37289 32011
rect 37323 32008 37335 32011
rect 37366 32008 37372 32020
rect 37323 31980 37372 32008
rect 37323 31977 37335 31980
rect 37277 31971 37335 31977
rect 37366 31968 37372 31980
rect 37424 31968 37430 32020
rect 38102 31968 38108 32020
rect 38160 31968 38166 32020
rect 39853 32011 39911 32017
rect 39853 31977 39865 32011
rect 39899 32008 39911 32011
rect 39942 32008 39948 32020
rect 39899 31980 39948 32008
rect 39899 31977 39911 31980
rect 39853 31971 39911 31977
rect 39942 31968 39948 31980
rect 40000 31968 40006 32020
rect 31202 31900 31208 31952
rect 31260 31940 31266 31952
rect 31570 31940 31576 31952
rect 31260 31912 31576 31940
rect 31260 31900 31266 31912
rect 31570 31900 31576 31912
rect 31628 31900 31634 31952
rect 33980 31940 34008 31968
rect 38746 31940 38752 31952
rect 33980 31912 35204 31940
rect 34790 31832 34796 31884
rect 34848 31872 34854 31884
rect 35069 31875 35127 31881
rect 35069 31872 35081 31875
rect 34848 31844 35081 31872
rect 34848 31832 34854 31844
rect 35069 31841 35081 31844
rect 35115 31841 35127 31875
rect 35176 31872 35204 31912
rect 37752 31912 38752 31940
rect 37752 31881 37780 31912
rect 38746 31900 38752 31912
rect 38804 31900 38810 31952
rect 41138 31940 41144 31952
rect 40328 31912 41144 31940
rect 37737 31875 37795 31881
rect 35176 31844 37688 31872
rect 35069 31835 35127 31841
rect 28994 31764 29000 31816
rect 29052 31804 29058 31816
rect 29733 31807 29791 31813
rect 29733 31804 29745 31807
rect 29052 31776 29745 31804
rect 29052 31764 29058 31776
rect 29733 31773 29745 31776
rect 29779 31773 29791 31807
rect 29733 31767 29791 31773
rect 30000 31807 30058 31813
rect 30000 31773 30012 31807
rect 30046 31804 30058 31807
rect 30374 31804 30380 31816
rect 30046 31776 30380 31804
rect 30046 31773 30058 31776
rect 30000 31767 30058 31773
rect 30374 31764 30380 31776
rect 30432 31764 30438 31816
rect 31754 31764 31760 31816
rect 31812 31804 31818 31816
rect 32585 31807 32643 31813
rect 32585 31804 32597 31807
rect 31812 31776 32597 31804
rect 31812 31764 31818 31776
rect 32585 31773 32597 31776
rect 32631 31804 32643 31807
rect 32766 31804 32772 31816
rect 32631 31776 32772 31804
rect 32631 31773 32643 31776
rect 32585 31767 32643 31773
rect 32766 31764 32772 31776
rect 32824 31804 32830 31816
rect 33045 31807 33103 31813
rect 33045 31804 33057 31807
rect 32824 31776 33057 31804
rect 32824 31764 32830 31776
rect 33045 31773 33057 31776
rect 33091 31773 33103 31807
rect 33045 31767 33103 31773
rect 33312 31807 33370 31813
rect 33312 31773 33324 31807
rect 33358 31804 33370 31807
rect 33686 31804 33692 31816
rect 33358 31776 33692 31804
rect 33358 31773 33370 31776
rect 33312 31767 33370 31773
rect 33686 31764 33692 31776
rect 33744 31764 33750 31816
rect 37660 31804 37688 31844
rect 37737 31841 37749 31875
rect 37783 31841 37795 31875
rect 37737 31835 37795 31841
rect 37829 31875 37887 31881
rect 37829 31841 37841 31875
rect 37875 31841 37887 31875
rect 37829 31835 37887 31841
rect 37844 31804 37872 31835
rect 38562 31832 38568 31884
rect 38620 31832 38626 31884
rect 38657 31875 38715 31881
rect 38657 31841 38669 31875
rect 38703 31841 38715 31875
rect 38657 31835 38715 31841
rect 39117 31875 39175 31881
rect 39117 31841 39129 31875
rect 39163 31872 39175 31875
rect 39482 31872 39488 31884
rect 39163 31844 39488 31872
rect 39163 31841 39175 31844
rect 39117 31835 39175 31841
rect 38672 31804 38700 31835
rect 39482 31832 39488 31844
rect 39540 31832 39546 31884
rect 40328 31881 40356 31912
rect 41138 31900 41144 31912
rect 41196 31900 41202 31952
rect 40313 31875 40371 31881
rect 39592 31844 40264 31872
rect 38930 31804 38936 31816
rect 37660 31776 38936 31804
rect 38930 31764 38936 31776
rect 38988 31804 38994 31816
rect 39592 31804 39620 31844
rect 38988 31776 39620 31804
rect 39669 31807 39727 31813
rect 38988 31764 38994 31776
rect 39669 31773 39681 31807
rect 39715 31804 39727 31807
rect 39942 31804 39948 31816
rect 39715 31776 39948 31804
rect 39715 31773 39727 31776
rect 39669 31767 39727 31773
rect 39942 31764 39948 31776
rect 40000 31764 40006 31816
rect 40236 31804 40264 31844
rect 40313 31841 40325 31875
rect 40359 31841 40371 31875
rect 40313 31835 40371 31841
rect 40405 31875 40463 31881
rect 40405 31841 40417 31875
rect 40451 31841 40463 31875
rect 40405 31835 40463 31841
rect 40420 31804 40448 31835
rect 40678 31832 40684 31884
rect 40736 31872 40742 31884
rect 41509 31875 41567 31881
rect 41509 31872 41521 31875
rect 40736 31844 41521 31872
rect 40736 31832 40742 31844
rect 41509 31841 41521 31844
rect 41555 31841 41567 31875
rect 41509 31835 41567 31841
rect 40494 31804 40500 31816
rect 40236 31776 40500 31804
rect 40494 31764 40500 31776
rect 40552 31764 40558 31816
rect 40770 31764 40776 31816
rect 40828 31764 40834 31816
rect 41414 31764 41420 31816
rect 41472 31764 41478 31816
rect 42150 31764 42156 31816
rect 42208 31764 42214 31816
rect 28905 31739 28963 31745
rect 28905 31705 28917 31739
rect 28951 31705 28963 31739
rect 28905 31699 28963 31705
rect 29178 31696 29184 31748
rect 29236 31736 29242 31748
rect 29273 31739 29331 31745
rect 29273 31736 29285 31739
rect 29236 31708 29285 31736
rect 29236 31696 29242 31708
rect 29273 31705 29285 31708
rect 29319 31736 29331 31739
rect 30282 31736 30288 31748
rect 29319 31708 30288 31736
rect 29319 31705 29331 31708
rect 29273 31699 29331 31705
rect 30282 31696 30288 31708
rect 30340 31696 30346 31748
rect 31938 31696 31944 31748
rect 31996 31736 32002 31748
rect 32318 31739 32376 31745
rect 32318 31736 32330 31739
rect 31996 31708 32330 31736
rect 31996 31696 32002 31708
rect 32318 31705 32330 31708
rect 32364 31705 32376 31739
rect 32318 31699 32376 31705
rect 35342 31696 35348 31748
rect 35400 31696 35406 31748
rect 35452 31708 35834 31736
rect 3326 31628 3332 31680
rect 3384 31628 3390 31680
rect 5166 31628 5172 31680
rect 5224 31668 5230 31680
rect 5461 31671 5519 31677
rect 5461 31668 5473 31671
rect 5224 31640 5473 31668
rect 5224 31628 5230 31640
rect 5461 31637 5473 31640
rect 5507 31637 5519 31671
rect 5461 31631 5519 31637
rect 8478 31628 8484 31680
rect 8536 31668 8542 31680
rect 10410 31668 10416 31680
rect 8536 31640 10416 31668
rect 8536 31628 8542 31640
rect 10410 31628 10416 31640
rect 10468 31628 10474 31680
rect 10870 31628 10876 31680
rect 10928 31628 10934 31680
rect 10962 31628 10968 31680
rect 11020 31628 11026 31680
rect 13446 31628 13452 31680
rect 13504 31628 13510 31680
rect 15930 31628 15936 31680
rect 15988 31628 15994 31680
rect 17586 31628 17592 31680
rect 17644 31668 17650 31680
rect 19518 31668 19524 31680
rect 17644 31640 19524 31668
rect 17644 31628 17650 31640
rect 19518 31628 19524 31640
rect 19576 31628 19582 31680
rect 28810 31628 28816 31680
rect 28868 31668 28874 31680
rect 28994 31668 29000 31680
rect 28868 31640 29000 31668
rect 28868 31628 28874 31640
rect 28994 31628 29000 31640
rect 29052 31628 29058 31680
rect 33502 31628 33508 31680
rect 33560 31668 33566 31680
rect 35452 31668 35480 31708
rect 33560 31640 35480 31668
rect 33560 31628 33566 31640
rect 36814 31628 36820 31680
rect 36872 31668 36878 31680
rect 37645 31671 37703 31677
rect 37645 31668 37657 31671
rect 36872 31640 37657 31668
rect 36872 31628 36878 31640
rect 37645 31637 37657 31640
rect 37691 31637 37703 31671
rect 37645 31631 37703 31637
rect 38470 31628 38476 31680
rect 38528 31628 38534 31680
rect 38654 31628 38660 31680
rect 38712 31668 38718 31680
rect 40221 31671 40279 31677
rect 40221 31668 40233 31671
rect 38712 31640 40233 31668
rect 38712 31628 38718 31640
rect 40221 31637 40233 31640
rect 40267 31637 40279 31671
rect 40221 31631 40279 31637
rect 1104 31578 42504 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 42504 31578
rect 1104 31504 42504 31526
rect 4062 31424 4068 31476
rect 4120 31464 4126 31476
rect 6178 31464 6184 31476
rect 4120 31436 6184 31464
rect 4120 31424 4126 31436
rect 6178 31424 6184 31436
rect 6236 31424 6242 31476
rect 7006 31424 7012 31476
rect 7064 31464 7070 31476
rect 7377 31467 7435 31473
rect 7377 31464 7389 31467
rect 7064 31436 7389 31464
rect 7064 31424 7070 31436
rect 7377 31433 7389 31436
rect 7423 31433 7435 31467
rect 8662 31464 8668 31476
rect 7377 31427 7435 31433
rect 7760 31436 8668 31464
rect 2406 31356 2412 31408
rect 2464 31356 2470 31408
rect 5902 31396 5908 31408
rect 5474 31368 5908 31396
rect 5902 31356 5908 31368
rect 5960 31356 5966 31408
rect 7760 31405 7788 31436
rect 8662 31424 8668 31436
rect 8720 31464 8726 31476
rect 9122 31464 9128 31476
rect 8720 31436 9128 31464
rect 8720 31424 8726 31436
rect 9122 31424 9128 31436
rect 9180 31424 9186 31476
rect 9309 31467 9367 31473
rect 9309 31433 9321 31467
rect 9355 31464 9367 31467
rect 9398 31464 9404 31476
rect 9355 31436 9404 31464
rect 9355 31433 9367 31436
rect 9309 31427 9367 31433
rect 9398 31424 9404 31436
rect 9456 31424 9462 31476
rect 14458 31424 14464 31476
rect 14516 31424 14522 31476
rect 15930 31424 15936 31476
rect 15988 31464 15994 31476
rect 16482 31464 16488 31476
rect 15988 31436 16488 31464
rect 15988 31424 15994 31436
rect 16482 31424 16488 31436
rect 16540 31464 16546 31476
rect 16945 31467 17003 31473
rect 16945 31464 16957 31467
rect 16540 31436 16957 31464
rect 16540 31424 16546 31436
rect 16945 31433 16957 31436
rect 16991 31433 17003 31467
rect 16945 31427 17003 31433
rect 17586 31424 17592 31476
rect 17644 31464 17650 31476
rect 17773 31467 17831 31473
rect 17773 31464 17785 31467
rect 17644 31436 17785 31464
rect 17644 31424 17650 31436
rect 17773 31433 17785 31436
rect 17819 31433 17831 31467
rect 21542 31464 21548 31476
rect 17773 31427 17831 31433
rect 17972 31436 21548 31464
rect 7745 31399 7803 31405
rect 7745 31365 7757 31399
rect 7791 31365 7803 31399
rect 7745 31359 7803 31365
rect 7883 31399 7941 31405
rect 7883 31365 7895 31399
rect 7929 31396 7941 31399
rect 8110 31396 8116 31408
rect 7929 31368 8116 31396
rect 7929 31365 7941 31368
rect 7883 31359 7941 31365
rect 8110 31356 8116 31368
rect 8168 31356 8174 31408
rect 8202 31356 8208 31408
rect 8260 31396 8266 31408
rect 8481 31399 8539 31405
rect 8481 31396 8493 31399
rect 8260 31368 8493 31396
rect 8260 31356 8266 31368
rect 8481 31365 8493 31368
rect 8527 31365 8539 31399
rect 8481 31359 8539 31365
rect 3050 31288 3056 31340
rect 3108 31328 3114 31340
rect 3694 31328 3700 31340
rect 3108 31300 3700 31328
rect 3108 31288 3114 31300
rect 3694 31288 3700 31300
rect 3752 31288 3758 31340
rect 7561 31331 7619 31337
rect 7561 31297 7573 31331
rect 7607 31297 7619 31331
rect 7561 31291 7619 31297
rect 7653 31331 7711 31337
rect 7653 31297 7665 31331
rect 7699 31297 7711 31331
rect 7653 31291 7711 31297
rect 8297 31331 8355 31337
rect 8297 31297 8309 31331
rect 8343 31297 8355 31331
rect 8496 31328 8524 31359
rect 8754 31356 8760 31408
rect 8812 31396 8818 31408
rect 9033 31399 9091 31405
rect 9033 31396 9045 31399
rect 8812 31368 9045 31396
rect 8812 31356 8818 31368
rect 9033 31365 9045 31368
rect 9079 31365 9091 31399
rect 9033 31359 9091 31365
rect 9582 31356 9588 31408
rect 9640 31356 9646 31408
rect 9677 31399 9735 31405
rect 9677 31365 9689 31399
rect 9723 31365 9735 31399
rect 9677 31359 9735 31365
rect 9815 31399 9873 31405
rect 9815 31365 9827 31399
rect 9861 31396 9873 31399
rect 9950 31396 9956 31408
rect 9861 31368 9956 31396
rect 9861 31365 9873 31368
rect 9815 31359 9873 31365
rect 8849 31331 8907 31337
rect 8849 31328 8861 31331
rect 8496 31300 8861 31328
rect 8297 31291 8355 31297
rect 8849 31297 8861 31300
rect 8895 31297 8907 31331
rect 8849 31291 8907 31297
rect 8941 31331 8999 31337
rect 8941 31297 8953 31331
rect 8987 31297 8999 31331
rect 8941 31291 8999 31297
rect 1397 31263 1455 31269
rect 1397 31229 1409 31263
rect 1443 31229 1455 31263
rect 1397 31223 1455 31229
rect 1673 31263 1731 31269
rect 1673 31229 1685 31263
rect 1719 31260 1731 31263
rect 2038 31260 2044 31272
rect 1719 31232 2044 31260
rect 1719 31229 1731 31232
rect 1673 31223 1731 31229
rect 1412 31136 1440 31223
rect 2038 31220 2044 31232
rect 2096 31220 2102 31272
rect 3145 31263 3203 31269
rect 3145 31229 3157 31263
rect 3191 31260 3203 31263
rect 3234 31260 3240 31272
rect 3191 31232 3240 31260
rect 3191 31229 3203 31232
rect 3145 31223 3203 31229
rect 3234 31220 3240 31232
rect 3292 31260 3298 31272
rect 3789 31263 3847 31269
rect 3789 31260 3801 31263
rect 3292 31232 3801 31260
rect 3292 31220 3298 31232
rect 3789 31229 3801 31232
rect 3835 31229 3847 31263
rect 3789 31223 3847 31229
rect 3973 31263 4031 31269
rect 3973 31229 3985 31263
rect 4019 31229 4031 31263
rect 3973 31223 4031 31229
rect 4249 31263 4307 31269
rect 4249 31229 4261 31263
rect 4295 31260 4307 31263
rect 4706 31260 4712 31272
rect 4295 31232 4712 31260
rect 4295 31229 4307 31232
rect 4249 31223 4307 31229
rect 3988 31192 4016 31223
rect 4706 31220 4712 31232
rect 4764 31220 4770 31272
rect 2746 31164 4016 31192
rect 7576 31192 7604 31291
rect 7668 31260 7696 31291
rect 7834 31260 7840 31272
rect 7668 31232 7840 31260
rect 7834 31220 7840 31232
rect 7892 31220 7898 31272
rect 8021 31263 8079 31269
rect 8021 31229 8033 31263
rect 8067 31260 8079 31263
rect 8312 31260 8340 31291
rect 8067 31232 8524 31260
rect 8067 31229 8079 31232
rect 8021 31223 8079 31229
rect 8496 31204 8524 31232
rect 8113 31195 8171 31201
rect 8113 31192 8125 31195
rect 7576 31164 8125 31192
rect 2746 31136 2774 31164
rect 1394 31084 1400 31136
rect 1452 31124 1458 31136
rect 2682 31124 2688 31136
rect 1452 31096 2688 31124
rect 1452 31084 1458 31096
rect 2682 31084 2688 31096
rect 2740 31096 2774 31136
rect 2740 31084 2746 31096
rect 2958 31084 2964 31136
rect 3016 31124 3022 31136
rect 3237 31127 3295 31133
rect 3237 31124 3249 31127
rect 3016 31096 3249 31124
rect 3016 31084 3022 31096
rect 3237 31093 3249 31096
rect 3283 31093 3295 31127
rect 3988 31124 4016 31164
rect 8113 31161 8125 31164
rect 8159 31161 8171 31195
rect 8113 31155 8171 31161
rect 8478 31152 8484 31204
rect 8536 31192 8542 31204
rect 8665 31195 8723 31201
rect 8665 31192 8677 31195
rect 8536 31164 8677 31192
rect 8536 31152 8542 31164
rect 8665 31161 8677 31164
rect 8711 31161 8723 31195
rect 8665 31155 8723 31161
rect 4614 31124 4620 31136
rect 3988 31096 4620 31124
rect 3237 31087 3295 31093
rect 4614 31084 4620 31096
rect 4672 31084 4678 31136
rect 5626 31084 5632 31136
rect 5684 31124 5690 31136
rect 5721 31127 5779 31133
rect 5721 31124 5733 31127
rect 5684 31096 5733 31124
rect 5684 31084 5690 31096
rect 5721 31093 5733 31096
rect 5767 31093 5779 31127
rect 8956 31124 8984 31291
rect 9490 31288 9496 31340
rect 9548 31288 9554 31340
rect 9122 31220 9128 31272
rect 9180 31260 9186 31272
rect 9692 31260 9720 31359
rect 9950 31356 9956 31368
rect 10008 31356 10014 31408
rect 12894 31356 12900 31408
rect 12952 31356 12958 31408
rect 15378 31356 15384 31408
rect 15436 31396 15442 31408
rect 16117 31399 16175 31405
rect 16117 31396 16129 31399
rect 15436 31368 16129 31396
rect 15436 31356 15442 31368
rect 16117 31365 16129 31368
rect 16163 31396 16175 31399
rect 17972 31396 18000 31436
rect 21542 31424 21548 31436
rect 21600 31424 21606 31476
rect 21634 31424 21640 31476
rect 21692 31464 21698 31476
rect 22097 31467 22155 31473
rect 22097 31464 22109 31467
rect 21692 31436 22109 31464
rect 21692 31424 21698 31436
rect 22097 31433 22109 31436
rect 22143 31464 22155 31467
rect 22186 31464 22192 31476
rect 22143 31436 22192 31464
rect 22143 31433 22155 31436
rect 22097 31427 22155 31433
rect 22186 31424 22192 31436
rect 22244 31424 22250 31476
rect 23290 31424 23296 31476
rect 23348 31464 23354 31476
rect 23937 31467 23995 31473
rect 23937 31464 23949 31467
rect 23348 31436 23949 31464
rect 23348 31424 23354 31436
rect 23937 31433 23949 31436
rect 23983 31433 23995 31467
rect 23937 31427 23995 31433
rect 24854 31424 24860 31476
rect 24912 31424 24918 31476
rect 25038 31424 25044 31476
rect 25096 31464 25102 31476
rect 25317 31467 25375 31473
rect 25317 31464 25329 31467
rect 25096 31436 25329 31464
rect 25096 31424 25102 31436
rect 25317 31433 25329 31436
rect 25363 31433 25375 31467
rect 25317 31427 25375 31433
rect 26053 31467 26111 31473
rect 26053 31433 26065 31467
rect 26099 31464 26111 31467
rect 26142 31464 26148 31476
rect 26099 31436 26148 31464
rect 26099 31433 26111 31436
rect 26053 31427 26111 31433
rect 26142 31424 26148 31436
rect 26200 31424 26206 31476
rect 30374 31424 30380 31476
rect 30432 31424 30438 31476
rect 30837 31467 30895 31473
rect 30837 31433 30849 31467
rect 30883 31464 30895 31467
rect 31018 31464 31024 31476
rect 30883 31436 31024 31464
rect 30883 31433 30895 31436
rect 30837 31427 30895 31433
rect 31018 31424 31024 31436
rect 31076 31424 31082 31476
rect 31205 31467 31263 31473
rect 31205 31433 31217 31467
rect 31251 31464 31263 31467
rect 31938 31464 31944 31476
rect 31251 31436 31944 31464
rect 31251 31433 31263 31436
rect 31205 31427 31263 31433
rect 31938 31424 31944 31436
rect 31996 31424 32002 31476
rect 32030 31424 32036 31476
rect 32088 31464 32094 31476
rect 32125 31467 32183 31473
rect 32125 31464 32137 31467
rect 32088 31436 32137 31464
rect 32088 31424 32094 31436
rect 32125 31433 32137 31436
rect 32171 31433 32183 31467
rect 32125 31427 32183 31433
rect 32582 31424 32588 31476
rect 32640 31424 32646 31476
rect 33318 31424 33324 31476
rect 33376 31424 33382 31476
rect 33689 31467 33747 31473
rect 33689 31433 33701 31467
rect 33735 31464 33747 31467
rect 33778 31464 33784 31476
rect 33735 31436 33784 31464
rect 33735 31433 33747 31436
rect 33689 31427 33747 31433
rect 33778 31424 33784 31436
rect 33836 31424 33842 31476
rect 41046 31424 41052 31476
rect 41104 31464 41110 31476
rect 41104 31436 41414 31464
rect 41104 31424 41110 31436
rect 16163 31368 18000 31396
rect 16163 31365 16175 31368
rect 16117 31359 16175 31365
rect 19150 31356 19156 31408
rect 19208 31396 19214 31408
rect 19245 31399 19303 31405
rect 19245 31396 19257 31399
rect 19208 31368 19257 31396
rect 19208 31356 19214 31368
rect 19245 31365 19257 31368
rect 19291 31365 19303 31399
rect 19245 31359 19303 31365
rect 23382 31356 23388 31408
rect 23440 31396 23446 31408
rect 26421 31399 26479 31405
rect 23440 31368 25452 31396
rect 23440 31356 23446 31368
rect 10962 31328 10968 31340
rect 10152 31300 10968 31328
rect 9180 31232 9720 31260
rect 9953 31263 10011 31269
rect 9180 31220 9186 31232
rect 9953 31229 9965 31263
rect 9999 31260 10011 31263
rect 10152 31260 10180 31300
rect 10962 31288 10968 31300
rect 11020 31288 11026 31340
rect 13446 31288 13452 31340
rect 13504 31288 13510 31340
rect 14829 31331 14887 31337
rect 14829 31297 14841 31331
rect 14875 31297 14887 31331
rect 14829 31291 14887 31297
rect 14921 31331 14979 31337
rect 14921 31297 14933 31331
rect 14967 31328 14979 31331
rect 15289 31331 15347 31337
rect 15289 31328 15301 31331
rect 14967 31300 15301 31328
rect 14967 31297 14979 31300
rect 14921 31291 14979 31297
rect 15289 31297 15301 31300
rect 15335 31297 15347 31331
rect 15289 31291 15347 31297
rect 9999 31232 10180 31260
rect 9999 31229 10011 31232
rect 9953 31223 10011 31229
rect 10226 31220 10232 31272
rect 10284 31220 10290 31272
rect 10321 31263 10379 31269
rect 10321 31229 10333 31263
rect 10367 31229 10379 31263
rect 10321 31223 10379 31229
rect 9217 31195 9275 31201
rect 9217 31161 9229 31195
rect 9263 31192 9275 31195
rect 9766 31192 9772 31204
rect 9263 31164 9772 31192
rect 9263 31161 9275 31164
rect 9217 31155 9275 31161
rect 9766 31152 9772 31164
rect 9824 31152 9830 31204
rect 9858 31152 9864 31204
rect 9916 31192 9922 31204
rect 10045 31195 10103 31201
rect 10045 31192 10057 31195
rect 9916 31164 10057 31192
rect 9916 31152 9922 31164
rect 10045 31161 10057 31164
rect 10091 31161 10103 31195
rect 10045 31155 10103 31161
rect 10134 31152 10140 31204
rect 10192 31192 10198 31204
rect 10336 31192 10364 31223
rect 10410 31220 10416 31272
rect 10468 31220 10474 31272
rect 10505 31263 10563 31269
rect 10505 31229 10517 31263
rect 10551 31260 10563 31263
rect 10870 31260 10876 31272
rect 10551 31232 10876 31260
rect 10551 31229 10563 31232
rect 10505 31223 10563 31229
rect 10192 31164 10364 31192
rect 10192 31152 10198 31164
rect 10520 31124 10548 31223
rect 10870 31220 10876 31232
rect 10928 31220 10934 31272
rect 11606 31220 11612 31272
rect 11664 31220 11670 31272
rect 11885 31263 11943 31269
rect 11885 31229 11897 31263
rect 11931 31260 11943 31263
rect 12618 31260 12624 31272
rect 11931 31232 12624 31260
rect 11931 31229 11943 31232
rect 11885 31223 11943 31229
rect 12618 31220 12624 31232
rect 12676 31220 12682 31272
rect 13357 31263 13415 31269
rect 13357 31229 13369 31263
rect 13403 31260 13415 31263
rect 13464 31260 13492 31288
rect 14001 31263 14059 31269
rect 14001 31260 14013 31263
rect 13403 31232 14013 31260
rect 13403 31229 13415 31232
rect 13357 31223 13415 31229
rect 14001 31229 14013 31232
rect 14047 31229 14059 31263
rect 14001 31223 14059 31229
rect 12986 31152 12992 31204
rect 13044 31192 13050 31204
rect 13449 31195 13507 31201
rect 13449 31192 13461 31195
rect 13044 31164 13461 31192
rect 13044 31152 13050 31164
rect 13449 31161 13461 31164
rect 13495 31161 13507 31195
rect 14844 31192 14872 31291
rect 15470 31288 15476 31340
rect 15528 31328 15534 31340
rect 15841 31331 15899 31337
rect 15841 31328 15853 31331
rect 15528 31300 15853 31328
rect 15528 31288 15534 31300
rect 15841 31297 15853 31300
rect 15887 31297 15899 31331
rect 15841 31291 15899 31297
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31297 17095 31331
rect 17037 31291 17095 31297
rect 15105 31263 15163 31269
rect 15105 31229 15117 31263
rect 15151 31260 15163 31263
rect 16393 31263 16451 31269
rect 16393 31260 16405 31263
rect 15151 31232 16405 31260
rect 15151 31229 15163 31232
rect 15105 31223 15163 31229
rect 16393 31229 16405 31232
rect 16439 31260 16451 31263
rect 16574 31260 16580 31272
rect 16439 31232 16580 31260
rect 16439 31229 16451 31232
rect 16393 31223 16451 31229
rect 16574 31220 16580 31232
rect 16632 31220 16638 31272
rect 16850 31220 16856 31272
rect 16908 31220 16914 31272
rect 17052 31192 17080 31291
rect 18138 31288 18144 31340
rect 18196 31288 18202 31340
rect 19521 31331 19579 31337
rect 19521 31297 19533 31331
rect 19567 31328 19579 31331
rect 19610 31328 19616 31340
rect 19567 31300 19616 31328
rect 19567 31297 19579 31300
rect 19521 31291 19579 31297
rect 19610 31288 19616 31300
rect 19668 31288 19674 31340
rect 21174 31288 21180 31340
rect 21232 31328 21238 31340
rect 22189 31331 22247 31337
rect 22189 31328 22201 31331
rect 21232 31300 22201 31328
rect 21232 31288 21238 31300
rect 22189 31297 22201 31300
rect 22235 31328 22247 31331
rect 22278 31328 22284 31340
rect 22235 31300 22284 31328
rect 22235 31297 22247 31300
rect 22189 31291 22247 31297
rect 22278 31288 22284 31300
rect 22336 31288 22342 31340
rect 23845 31331 23903 31337
rect 23845 31297 23857 31331
rect 23891 31328 23903 31331
rect 24118 31328 24124 31340
rect 23891 31300 24124 31328
rect 23891 31297 23903 31300
rect 23845 31291 23903 31297
rect 24118 31288 24124 31300
rect 24176 31288 24182 31340
rect 25222 31288 25228 31340
rect 25280 31288 25286 31340
rect 19702 31260 19708 31272
rect 14844 31164 17080 31192
rect 17328 31232 19708 31260
rect 13449 31155 13507 31161
rect 16592 31136 16620 31164
rect 8956 31096 10548 31124
rect 5721 31087 5779 31093
rect 16574 31084 16580 31136
rect 16632 31084 16638 31136
rect 16850 31084 16856 31136
rect 16908 31124 16914 31136
rect 17328 31124 17356 31232
rect 19702 31220 19708 31232
rect 19760 31260 19766 31272
rect 21913 31263 21971 31269
rect 21913 31260 21925 31263
rect 19760 31232 21925 31260
rect 19760 31220 19766 31232
rect 21913 31229 21925 31232
rect 21959 31260 21971 31263
rect 24029 31263 24087 31269
rect 24029 31260 24041 31263
rect 21959 31232 24041 31260
rect 21959 31229 21971 31232
rect 21913 31223 21971 31229
rect 24029 31229 24041 31232
rect 24075 31260 24087 31263
rect 24210 31260 24216 31272
rect 24075 31232 24216 31260
rect 24075 31229 24087 31232
rect 24029 31223 24087 31229
rect 24210 31220 24216 31232
rect 24268 31220 24274 31272
rect 25424 31269 25452 31368
rect 26421 31365 26433 31399
rect 26467 31396 26479 31399
rect 26786 31396 26792 31408
rect 26467 31368 26792 31396
rect 26467 31365 26479 31368
rect 26421 31359 26479 31365
rect 26786 31356 26792 31368
rect 26844 31356 26850 31408
rect 28077 31399 28135 31405
rect 28077 31365 28089 31399
rect 28123 31396 28135 31399
rect 28350 31396 28356 31408
rect 28123 31368 28356 31396
rect 28123 31365 28135 31368
rect 28077 31359 28135 31365
rect 28350 31356 28356 31368
rect 28408 31356 28414 31408
rect 29178 31396 29184 31408
rect 28920 31368 29184 31396
rect 26513 31331 26571 31337
rect 26513 31297 26525 31331
rect 26559 31328 26571 31331
rect 26973 31331 27031 31337
rect 26973 31328 26985 31331
rect 26559 31300 26985 31328
rect 26559 31297 26571 31300
rect 26513 31291 26571 31297
rect 26973 31297 26985 31300
rect 27019 31297 27031 31331
rect 26973 31291 27031 31297
rect 27246 31288 27252 31340
rect 27304 31328 27310 31340
rect 27525 31331 27583 31337
rect 27525 31328 27537 31331
rect 27304 31300 27537 31328
rect 27304 31288 27310 31300
rect 27525 31297 27537 31300
rect 27571 31297 27583 31331
rect 27525 31291 27583 31297
rect 28810 31288 28816 31340
rect 28868 31288 28874 31340
rect 25409 31263 25467 31269
rect 25409 31229 25421 31263
rect 25455 31229 25467 31263
rect 25409 31223 25467 31229
rect 26050 31220 26056 31272
rect 26108 31260 26114 31272
rect 26605 31263 26663 31269
rect 26605 31260 26617 31263
rect 26108 31232 26617 31260
rect 26108 31220 26114 31232
rect 26605 31229 26617 31232
rect 26651 31229 26663 31263
rect 26605 31223 26663 31229
rect 28166 31220 28172 31272
rect 28224 31220 28230 31272
rect 28353 31263 28411 31269
rect 28353 31229 28365 31263
rect 28399 31260 28411 31263
rect 28920 31260 28948 31368
rect 29178 31356 29184 31368
rect 29236 31356 29242 31408
rect 29454 31356 29460 31408
rect 29512 31396 29518 31408
rect 30190 31396 30196 31408
rect 29512 31368 30196 31396
rect 29512 31356 29518 31368
rect 30190 31356 30196 31368
rect 30248 31356 30254 31408
rect 31573 31399 31631 31405
rect 31573 31365 31585 31399
rect 31619 31396 31631 31399
rect 33134 31396 33140 31408
rect 31619 31368 33140 31396
rect 31619 31365 31631 31368
rect 31573 31359 31631 31365
rect 33134 31356 33140 31368
rect 33192 31356 33198 31408
rect 37918 31356 37924 31408
rect 37976 31396 37982 31408
rect 40402 31396 40408 31408
rect 37976 31368 39344 31396
rect 37976 31356 37982 31368
rect 29080 31331 29138 31337
rect 29080 31297 29092 31331
rect 29126 31328 29138 31331
rect 29546 31328 29552 31340
rect 29126 31300 29552 31328
rect 29126 31297 29138 31300
rect 29080 31291 29138 31297
rect 29546 31288 29552 31300
rect 29604 31288 29610 31340
rect 30745 31331 30803 31337
rect 30745 31297 30757 31331
rect 30791 31328 30803 31331
rect 32398 31328 32404 31340
rect 30791 31300 32404 31328
rect 30791 31297 30803 31300
rect 30745 31291 30803 31297
rect 32398 31288 32404 31300
rect 32456 31288 32462 31340
rect 32493 31331 32551 31337
rect 32493 31297 32505 31331
rect 32539 31328 32551 31331
rect 32674 31328 32680 31340
rect 32539 31300 32680 31328
rect 32539 31297 32551 31300
rect 32493 31291 32551 31297
rect 32674 31288 32680 31300
rect 32732 31288 32738 31340
rect 33781 31331 33839 31337
rect 33781 31297 33793 31331
rect 33827 31328 33839 31331
rect 34149 31331 34207 31337
rect 34149 31328 34161 31331
rect 33827 31300 34161 31328
rect 33827 31297 33839 31300
rect 33781 31291 33839 31297
rect 34149 31297 34161 31300
rect 34195 31297 34207 31331
rect 34149 31291 34207 31297
rect 34238 31288 34244 31340
rect 34296 31328 34302 31340
rect 39316 31337 39344 31368
rect 39868 31368 40408 31396
rect 34701 31331 34759 31337
rect 34701 31328 34713 31331
rect 34296 31300 34713 31328
rect 34296 31288 34302 31300
rect 34701 31297 34713 31300
rect 34747 31297 34759 31331
rect 34701 31291 34759 31297
rect 39045 31331 39103 31337
rect 39045 31297 39057 31331
rect 39091 31328 39103 31331
rect 39301 31331 39359 31337
rect 39091 31300 39252 31328
rect 39091 31297 39103 31300
rect 39045 31291 39103 31297
rect 28399 31232 28948 31260
rect 31021 31263 31079 31269
rect 28399 31229 28411 31232
rect 28353 31223 28411 31229
rect 31021 31229 31033 31263
rect 31067 31229 31079 31263
rect 31021 31223 31079 31229
rect 30282 31152 30288 31204
rect 30340 31192 30346 31204
rect 31036 31192 31064 31223
rect 31662 31220 31668 31272
rect 31720 31220 31726 31272
rect 31849 31263 31907 31269
rect 31849 31229 31861 31263
rect 31895 31260 31907 31263
rect 32769 31263 32827 31269
rect 32769 31260 32781 31263
rect 31895 31232 32781 31260
rect 31895 31229 31907 31232
rect 31849 31223 31907 31229
rect 32769 31229 32781 31232
rect 32815 31260 32827 31263
rect 33042 31260 33048 31272
rect 32815 31232 33048 31260
rect 32815 31229 32827 31232
rect 32769 31223 32827 31229
rect 31864 31192 31892 31223
rect 33042 31220 33048 31232
rect 33100 31220 33106 31272
rect 33962 31220 33968 31272
rect 34020 31220 34026 31272
rect 39224 31260 39252 31300
rect 39301 31297 39313 31331
rect 39347 31328 39359 31331
rect 39666 31328 39672 31340
rect 39724 31337 39730 31340
rect 39347 31300 39672 31328
rect 39347 31297 39359 31300
rect 39301 31291 39359 31297
rect 39666 31288 39672 31300
rect 39724 31328 39734 31337
rect 39868 31328 39896 31368
rect 40402 31356 40408 31368
rect 40460 31356 40466 31408
rect 39724 31300 39896 31328
rect 39936 31331 39994 31337
rect 39724 31291 39734 31300
rect 39936 31297 39948 31331
rect 39982 31328 39994 31331
rect 40954 31328 40960 31340
rect 39982 31300 40960 31328
rect 39982 31297 39994 31300
rect 39936 31291 39994 31297
rect 39724 31288 39730 31291
rect 40954 31288 40960 31300
rect 41012 31288 41018 31340
rect 41386 31328 41414 31436
rect 41785 31331 41843 31337
rect 41785 31328 41797 31331
rect 41386 31300 41797 31328
rect 41785 31297 41797 31300
rect 41831 31297 41843 31331
rect 41785 31291 41843 31297
rect 39224 31232 39712 31260
rect 30340 31164 31892 31192
rect 30340 31152 30346 31164
rect 16908 31096 17356 31124
rect 16908 31084 16914 31096
rect 17402 31084 17408 31136
rect 17460 31124 17466 31136
rect 18230 31124 18236 31136
rect 17460 31096 18236 31124
rect 17460 31084 17466 31096
rect 18230 31084 18236 31096
rect 18288 31084 18294 31136
rect 21818 31084 21824 31136
rect 21876 31124 21882 31136
rect 22557 31127 22615 31133
rect 22557 31124 22569 31127
rect 21876 31096 22569 31124
rect 21876 31084 21882 31096
rect 22557 31093 22569 31096
rect 22603 31124 22615 31127
rect 22646 31124 22652 31136
rect 22603 31096 22652 31124
rect 22603 31093 22615 31096
rect 22557 31087 22615 31093
rect 22646 31084 22652 31096
rect 22704 31084 22710 31136
rect 23477 31127 23535 31133
rect 23477 31093 23489 31127
rect 23523 31124 23535 31127
rect 24026 31124 24032 31136
rect 23523 31096 24032 31124
rect 23523 31093 23535 31096
rect 23477 31087 23535 31093
rect 24026 31084 24032 31096
rect 24084 31084 24090 31136
rect 27709 31127 27767 31133
rect 27709 31093 27721 31127
rect 27755 31124 27767 31127
rect 28258 31124 28264 31136
rect 27755 31096 28264 31124
rect 27755 31093 27767 31096
rect 27709 31087 27767 31093
rect 28258 31084 28264 31096
rect 28316 31084 28322 31136
rect 30193 31127 30251 31133
rect 30193 31093 30205 31127
rect 30239 31124 30251 31127
rect 30926 31124 30932 31136
rect 30239 31096 30932 31124
rect 30239 31093 30251 31096
rect 30193 31087 30251 31093
rect 30926 31084 30932 31096
rect 30984 31084 30990 31136
rect 37921 31127 37979 31133
rect 37921 31093 37933 31127
rect 37967 31124 37979 31127
rect 39482 31124 39488 31136
rect 37967 31096 39488 31124
rect 37967 31093 37979 31096
rect 37921 31087 37979 31093
rect 39482 31084 39488 31096
rect 39540 31084 39546 31136
rect 39684 31124 39712 31232
rect 40034 31124 40040 31136
rect 39684 31096 40040 31124
rect 40034 31084 40040 31096
rect 40092 31084 40098 31136
rect 41230 31084 41236 31136
rect 41288 31084 41294 31136
rect 1104 31034 42504 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 42504 31034
rect 1104 30960 42504 30982
rect 1765 30923 1823 30929
rect 1765 30889 1777 30923
rect 1811 30889 1823 30923
rect 1765 30883 1823 30889
rect 1949 30923 2007 30929
rect 1949 30889 1961 30923
rect 1995 30920 2007 30923
rect 2866 30920 2872 30932
rect 1995 30892 2872 30920
rect 1995 30889 2007 30892
rect 1949 30883 2007 30889
rect 1780 30852 1808 30883
rect 2866 30880 2872 30892
rect 2924 30880 2930 30932
rect 4341 30923 4399 30929
rect 4341 30889 4353 30923
rect 4387 30920 4399 30923
rect 4706 30920 4712 30932
rect 4387 30892 4712 30920
rect 4387 30889 4399 30892
rect 4341 30883 4399 30889
rect 4706 30880 4712 30892
rect 4764 30880 4770 30932
rect 5166 30880 5172 30932
rect 5224 30920 5230 30932
rect 5810 30920 5816 30932
rect 5224 30892 5816 30920
rect 5224 30880 5230 30892
rect 5810 30880 5816 30892
rect 5868 30880 5874 30932
rect 7834 30880 7840 30932
rect 7892 30880 7898 30932
rect 8754 30880 8760 30932
rect 8812 30920 8818 30932
rect 10226 30920 10232 30932
rect 8812 30892 10232 30920
rect 8812 30880 8818 30892
rect 10226 30880 10232 30892
rect 10284 30920 10290 30932
rect 10689 30923 10747 30929
rect 10689 30920 10701 30923
rect 10284 30892 10701 30920
rect 10284 30880 10290 30892
rect 10689 30889 10701 30892
rect 10735 30889 10747 30923
rect 10689 30883 10747 30889
rect 12618 30880 12624 30932
rect 12676 30880 12682 30932
rect 16666 30880 16672 30932
rect 16724 30920 16730 30932
rect 17037 30923 17095 30929
rect 17037 30920 17049 30923
rect 16724 30892 17049 30920
rect 16724 30880 16730 30892
rect 17037 30889 17049 30892
rect 17083 30889 17095 30923
rect 19886 30920 19892 30932
rect 17037 30883 17095 30889
rect 18524 30892 19892 30920
rect 2590 30852 2596 30864
rect 1780 30824 2596 30852
rect 2590 30812 2596 30824
rect 2648 30812 2654 30864
rect 5442 30852 5448 30864
rect 3896 30824 5448 30852
rect 2038 30744 2044 30796
rect 2096 30744 2102 30796
rect 2869 30787 2927 30793
rect 2869 30784 2881 30787
rect 2240 30756 2881 30784
rect 2240 30725 2268 30756
rect 2869 30753 2881 30756
rect 2915 30753 2927 30787
rect 2869 30747 2927 30753
rect 2958 30744 2964 30796
rect 3016 30744 3022 30796
rect 3050 30744 3056 30796
rect 3108 30744 3114 30796
rect 3145 30787 3203 30793
rect 3145 30753 3157 30787
rect 3191 30784 3203 30787
rect 3418 30784 3424 30796
rect 3191 30756 3424 30784
rect 3191 30753 3203 30756
rect 3145 30747 3203 30753
rect 3418 30744 3424 30756
rect 3476 30744 3482 30796
rect 3896 30793 3924 30824
rect 5442 30812 5448 30824
rect 5500 30812 5506 30864
rect 5629 30855 5687 30861
rect 5629 30821 5641 30855
rect 5675 30852 5687 30855
rect 5718 30852 5724 30864
rect 5675 30824 5724 30852
rect 5675 30821 5687 30824
rect 5629 30815 5687 30821
rect 5718 30812 5724 30824
rect 5776 30812 5782 30864
rect 18325 30855 18383 30861
rect 18325 30852 18337 30855
rect 17328 30824 18337 30852
rect 3881 30787 3939 30793
rect 3881 30753 3893 30787
rect 3927 30753 3939 30787
rect 3881 30747 3939 30753
rect 3973 30787 4031 30793
rect 3973 30753 3985 30787
rect 4019 30784 4031 30787
rect 4798 30784 4804 30796
rect 4019 30756 4804 30784
rect 4019 30753 4031 30756
rect 3973 30747 4031 30753
rect 4798 30744 4804 30756
rect 4856 30744 4862 30796
rect 6638 30784 6644 30796
rect 4908 30756 6644 30784
rect 2225 30719 2283 30725
rect 1811 30685 1869 30691
rect 1811 30682 1823 30685
rect 1578 30608 1584 30660
rect 1636 30608 1642 30660
rect 1796 30651 1823 30682
rect 1857 30660 1869 30685
rect 2225 30685 2237 30719
rect 2271 30685 2283 30719
rect 2225 30679 2283 30685
rect 2685 30719 2743 30725
rect 2685 30685 2697 30719
rect 2731 30716 2743 30719
rect 2976 30716 3004 30744
rect 2731 30688 3004 30716
rect 2731 30685 2743 30688
rect 2685 30679 2743 30685
rect 3234 30676 3240 30728
rect 3292 30676 3298 30728
rect 3329 30719 3387 30725
rect 3329 30685 3341 30719
rect 3375 30685 3387 30719
rect 3329 30679 3387 30685
rect 4065 30719 4123 30725
rect 4065 30685 4077 30719
rect 4111 30685 4123 30719
rect 4065 30679 4123 30685
rect 4157 30719 4215 30725
rect 4157 30685 4169 30719
rect 4203 30685 4215 30719
rect 4157 30679 4215 30685
rect 1857 30651 1860 30660
rect 1796 30620 1860 30651
rect 1854 30608 1860 30620
rect 1912 30608 1918 30660
rect 2317 30651 2375 30657
rect 2317 30617 2329 30651
rect 2363 30617 2375 30651
rect 2317 30611 2375 30617
rect 2332 30580 2360 30611
rect 2406 30608 2412 30660
rect 2464 30608 2470 30660
rect 2547 30651 2605 30657
rect 2547 30617 2559 30651
rect 2593 30648 2605 30651
rect 2958 30648 2964 30660
rect 2593 30620 2964 30648
rect 2593 30617 2605 30620
rect 2547 30611 2605 30617
rect 2958 30608 2964 30620
rect 3016 30608 3022 30660
rect 3344 30648 3372 30679
rect 3878 30648 3884 30660
rect 3344 30620 3884 30648
rect 3878 30608 3884 30620
rect 3936 30608 3942 30660
rect 3326 30580 3332 30592
rect 2332 30552 3332 30580
rect 3326 30540 3332 30552
rect 3384 30540 3390 30592
rect 4080 30580 4108 30679
rect 4172 30648 4200 30679
rect 4614 30676 4620 30728
rect 4672 30716 4678 30728
rect 4908 30725 4936 30756
rect 6638 30744 6644 30756
rect 6696 30784 6702 30796
rect 8941 30787 8999 30793
rect 8941 30784 8953 30787
rect 6696 30756 8953 30784
rect 6696 30744 6702 30756
rect 8941 30753 8953 30756
rect 8987 30753 8999 30787
rect 8941 30747 8999 30753
rect 13265 30787 13323 30793
rect 13265 30753 13277 30787
rect 13311 30784 13323 30787
rect 13354 30784 13360 30796
rect 13311 30756 13360 30784
rect 13311 30753 13323 30756
rect 13265 30747 13323 30753
rect 13354 30744 13360 30756
rect 13412 30744 13418 30796
rect 4893 30719 4951 30725
rect 4893 30716 4905 30719
rect 4672 30688 4905 30716
rect 4672 30676 4678 30688
rect 4893 30685 4905 30688
rect 4939 30685 4951 30719
rect 4893 30679 4951 30685
rect 5077 30719 5135 30725
rect 5077 30685 5089 30719
rect 5123 30716 5135 30719
rect 5166 30716 5172 30728
rect 5123 30688 5172 30716
rect 5123 30685 5135 30688
rect 5077 30679 5135 30685
rect 5166 30676 5172 30688
rect 5224 30676 5230 30728
rect 5537 30719 5595 30725
rect 5537 30685 5549 30719
rect 5583 30716 5595 30719
rect 5718 30716 5724 30728
rect 5583 30688 5724 30716
rect 5583 30685 5595 30688
rect 5537 30679 5595 30685
rect 5718 30676 5724 30688
rect 5776 30676 5782 30728
rect 5810 30676 5816 30728
rect 5868 30676 5874 30728
rect 6178 30676 6184 30728
rect 6236 30676 6242 30728
rect 7745 30719 7803 30725
rect 7745 30685 7757 30719
rect 7791 30685 7803 30719
rect 7745 30679 7803 30685
rect 7929 30719 7987 30725
rect 7929 30685 7941 30719
rect 7975 30716 7987 30719
rect 8478 30716 8484 30728
rect 7975 30688 8484 30716
rect 7975 30685 7987 30688
rect 7929 30679 7987 30685
rect 4706 30648 4712 30660
rect 4172 30620 4712 30648
rect 4706 30608 4712 30620
rect 4764 30608 4770 30660
rect 6273 30651 6331 30657
rect 6273 30648 6285 30651
rect 4816 30620 6285 30648
rect 4816 30580 4844 30620
rect 6273 30617 6285 30620
rect 6319 30617 6331 30651
rect 7760 30648 7788 30679
rect 8478 30676 8484 30688
rect 8536 30676 8542 30728
rect 8754 30676 8760 30728
rect 8812 30676 8818 30728
rect 12986 30676 12992 30728
rect 13044 30676 13050 30728
rect 13446 30676 13452 30728
rect 13504 30676 13510 30728
rect 13538 30676 13544 30728
rect 13596 30716 13602 30728
rect 13633 30719 13691 30725
rect 13633 30716 13645 30719
rect 13596 30688 13645 30716
rect 13596 30676 13602 30688
rect 13633 30685 13645 30688
rect 13679 30685 13691 30719
rect 13633 30679 13691 30685
rect 17218 30676 17224 30728
rect 17276 30676 17282 30728
rect 17328 30725 17356 30824
rect 18325 30821 18337 30824
rect 18371 30821 18383 30855
rect 18325 30815 18383 30821
rect 17494 30744 17500 30796
rect 17552 30784 17558 30796
rect 18524 30784 18552 30892
rect 19886 30880 19892 30892
rect 19944 30920 19950 30932
rect 21542 30920 21548 30932
rect 19944 30892 21548 30920
rect 19944 30880 19950 30892
rect 21542 30880 21548 30892
rect 21600 30880 21606 30932
rect 22094 30880 22100 30932
rect 22152 30880 22158 30932
rect 23845 30923 23903 30929
rect 23845 30889 23857 30923
rect 23891 30920 23903 30923
rect 24578 30920 24584 30932
rect 23891 30892 24584 30920
rect 23891 30889 23903 30892
rect 23845 30883 23903 30889
rect 24578 30880 24584 30892
rect 24636 30880 24642 30932
rect 24679 30892 27108 30920
rect 18874 30812 18880 30864
rect 18932 30852 18938 30864
rect 19702 30852 19708 30864
rect 18932 30824 19708 30852
rect 18932 30812 18938 30824
rect 19702 30812 19708 30824
rect 19760 30812 19766 30864
rect 20254 30852 20260 30864
rect 19812 30824 20260 30852
rect 19426 30784 19432 30796
rect 17552 30756 18552 30784
rect 18616 30756 19432 30784
rect 17552 30744 17558 30756
rect 17313 30719 17371 30725
rect 17313 30685 17325 30719
rect 17359 30685 17371 30719
rect 17313 30679 17371 30685
rect 17589 30719 17647 30725
rect 17589 30685 17601 30719
rect 17635 30716 17647 30719
rect 17862 30716 17868 30728
rect 17635 30688 17868 30716
rect 17635 30685 17647 30688
rect 17589 30679 17647 30685
rect 17862 30676 17868 30688
rect 17920 30676 17926 30728
rect 18616 30725 18644 30756
rect 19426 30744 19432 30756
rect 19484 30784 19490 30796
rect 19812 30784 19840 30824
rect 20254 30812 20260 30824
rect 20312 30812 20318 30864
rect 22186 30852 22192 30864
rect 20456 30824 22192 30852
rect 19484 30756 19840 30784
rect 19484 30744 19490 30756
rect 19886 30744 19892 30796
rect 19944 30744 19950 30796
rect 19978 30744 19984 30796
rect 20036 30784 20042 30796
rect 20456 30784 20484 30824
rect 22186 30812 22192 30824
rect 22244 30812 22250 30864
rect 23658 30812 23664 30864
rect 23716 30852 23722 30864
rect 24679 30852 24707 30892
rect 23716 30824 24707 30852
rect 27080 30852 27108 30892
rect 27706 30880 27712 30932
rect 27764 30880 27770 30932
rect 28166 30880 28172 30932
rect 28224 30920 28230 30932
rect 28445 30923 28503 30929
rect 28445 30920 28457 30923
rect 28224 30892 28457 30920
rect 28224 30880 28230 30892
rect 28445 30889 28457 30892
rect 28491 30889 28503 30923
rect 28445 30883 28503 30889
rect 29546 30880 29552 30932
rect 29604 30880 29610 30932
rect 31662 30880 31668 30932
rect 31720 30920 31726 30932
rect 31941 30923 31999 30929
rect 31941 30920 31953 30923
rect 31720 30892 31953 30920
rect 31720 30880 31726 30892
rect 31941 30889 31953 30892
rect 31987 30889 31999 30923
rect 31941 30883 31999 30889
rect 35253 30923 35311 30929
rect 35253 30889 35265 30923
rect 35299 30920 35311 30923
rect 35342 30920 35348 30932
rect 35299 30892 35348 30920
rect 35299 30889 35311 30892
rect 35253 30883 35311 30889
rect 35342 30880 35348 30892
rect 35400 30880 35406 30932
rect 38838 30880 38844 30932
rect 38896 30920 38902 30932
rect 39209 30923 39267 30929
rect 39209 30920 39221 30923
rect 38896 30892 39221 30920
rect 38896 30880 38902 30892
rect 39209 30889 39221 30892
rect 39255 30920 39267 30923
rect 39482 30920 39488 30932
rect 39255 30892 39488 30920
rect 39255 30889 39267 30892
rect 39209 30883 39267 30889
rect 39482 30880 39488 30892
rect 39540 30880 39546 30932
rect 41414 30880 41420 30932
rect 41472 30920 41478 30932
rect 41782 30920 41788 30932
rect 41472 30892 41788 30920
rect 41472 30880 41478 30892
rect 41782 30880 41788 30892
rect 41840 30920 41846 30932
rect 42153 30923 42211 30929
rect 42153 30920 42165 30923
rect 41840 30892 42165 30920
rect 41840 30880 41846 30892
rect 42153 30889 42165 30892
rect 42199 30889 42211 30923
rect 42153 30883 42211 30889
rect 27080 30824 32168 30852
rect 23716 30812 23722 30824
rect 20036 30756 20484 30784
rect 20036 30744 20042 30756
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30685 18567 30719
rect 18509 30679 18567 30685
rect 18601 30719 18659 30725
rect 18601 30685 18613 30719
rect 18647 30685 18659 30719
rect 18601 30679 18659 30685
rect 18693 30719 18751 30725
rect 18693 30685 18705 30719
rect 18739 30716 18751 30719
rect 18782 30716 18788 30728
rect 18739 30688 18788 30716
rect 18739 30685 18751 30688
rect 18693 30679 18751 30685
rect 8202 30648 8208 30660
rect 7760 30620 8208 30648
rect 6273 30611 6331 30617
rect 8202 30608 8208 30620
rect 8260 30648 8266 30660
rect 8573 30651 8631 30657
rect 8573 30648 8585 30651
rect 8260 30620 8585 30648
rect 8260 30608 8266 30620
rect 8573 30617 8585 30620
rect 8619 30648 8631 30651
rect 8619 30620 9168 30648
rect 8619 30617 8631 30620
rect 8573 30611 8631 30617
rect 4080 30552 4844 30580
rect 5169 30583 5227 30589
rect 5169 30549 5181 30583
rect 5215 30580 5227 30583
rect 5810 30580 5816 30592
rect 5215 30552 5816 30580
rect 5215 30549 5227 30552
rect 5169 30543 5227 30549
rect 5810 30540 5816 30552
rect 5868 30540 5874 30592
rect 5997 30583 6055 30589
rect 5997 30549 6009 30583
rect 6043 30580 6055 30583
rect 6546 30580 6552 30592
rect 6043 30552 6552 30580
rect 6043 30549 6055 30552
rect 5997 30543 6055 30549
rect 6546 30540 6552 30552
rect 6604 30540 6610 30592
rect 8662 30540 8668 30592
rect 8720 30540 8726 30592
rect 9140 30580 9168 30620
rect 9214 30608 9220 30660
rect 9272 30608 9278 30660
rect 10502 30648 10508 30660
rect 10442 30620 10508 30648
rect 10502 30608 10508 30620
rect 10560 30648 10566 30660
rect 10962 30648 10968 30660
rect 10560 30620 10968 30648
rect 10560 30608 10566 30620
rect 10962 30608 10968 30620
rect 11020 30608 11026 30660
rect 18046 30608 18052 30660
rect 18104 30648 18110 30660
rect 18141 30651 18199 30657
rect 18141 30648 18153 30651
rect 18104 30620 18153 30648
rect 18104 30608 18110 30620
rect 18141 30617 18153 30620
rect 18187 30617 18199 30651
rect 18524 30648 18552 30679
rect 18782 30676 18788 30688
rect 18840 30676 18846 30728
rect 18877 30719 18935 30725
rect 18877 30685 18889 30719
rect 18923 30716 18935 30719
rect 19058 30716 19064 30728
rect 18923 30688 19064 30716
rect 18923 30685 18935 30688
rect 18877 30679 18935 30685
rect 19058 30676 19064 30688
rect 19116 30676 19122 30728
rect 19610 30676 19616 30728
rect 19668 30676 19674 30728
rect 19702 30676 19708 30728
rect 19760 30716 19766 30728
rect 20364 30725 20392 30756
rect 20622 30744 20628 30796
rect 20680 30784 20686 30796
rect 22281 30787 22339 30793
rect 22281 30784 22293 30787
rect 20680 30756 22293 30784
rect 20680 30744 20686 30756
rect 20073 30719 20131 30725
rect 20073 30716 20085 30719
rect 19760 30688 20085 30716
rect 19760 30676 19766 30688
rect 20073 30685 20085 30688
rect 20119 30685 20131 30719
rect 20073 30679 20131 30685
rect 20166 30719 20224 30725
rect 20166 30685 20178 30719
rect 20212 30685 20224 30719
rect 20166 30679 20224 30685
rect 20349 30719 20407 30725
rect 20349 30685 20361 30719
rect 20395 30685 20407 30719
rect 20349 30679 20407 30685
rect 19628 30648 19656 30676
rect 18524 30620 19656 30648
rect 18141 30611 18199 30617
rect 19886 30608 19892 30660
rect 19944 30648 19950 30660
rect 20180 30648 20208 30679
rect 20438 30676 20444 30728
rect 20496 30676 20502 30728
rect 20530 30676 20536 30728
rect 20588 30725 20594 30728
rect 20588 30716 20596 30725
rect 20588 30688 21036 30716
rect 20588 30679 20596 30688
rect 20588 30676 20594 30679
rect 19944 30620 20208 30648
rect 19944 30608 19950 30620
rect 10134 30580 10140 30592
rect 9140 30552 10140 30580
rect 10134 30540 10140 30552
rect 10192 30540 10198 30592
rect 13081 30583 13139 30589
rect 13081 30549 13093 30583
rect 13127 30580 13139 30583
rect 13170 30580 13176 30592
rect 13127 30552 13176 30580
rect 13127 30549 13139 30552
rect 13081 30543 13139 30549
rect 13170 30540 13176 30552
rect 13228 30540 13234 30592
rect 13541 30583 13599 30589
rect 13541 30549 13553 30583
rect 13587 30580 13599 30583
rect 15194 30580 15200 30592
rect 13587 30552 15200 30580
rect 13587 30549 13599 30552
rect 13541 30543 13599 30549
rect 15194 30540 15200 30552
rect 15252 30540 15258 30592
rect 17586 30540 17592 30592
rect 17644 30580 17650 30592
rect 17865 30583 17923 30589
rect 17865 30580 17877 30583
rect 17644 30552 17877 30580
rect 17644 30540 17650 30552
rect 17865 30549 17877 30552
rect 17911 30580 17923 30583
rect 18414 30580 18420 30592
rect 17911 30552 18420 30580
rect 17911 30549 17923 30552
rect 17865 30543 17923 30549
rect 18414 30540 18420 30552
rect 18472 30540 18478 30592
rect 19150 30540 19156 30592
rect 19208 30580 19214 30592
rect 19245 30583 19303 30589
rect 19245 30580 19257 30583
rect 19208 30552 19257 30580
rect 19208 30540 19214 30552
rect 19245 30549 19257 30552
rect 19291 30549 19303 30583
rect 19245 30543 19303 30549
rect 19518 30540 19524 30592
rect 19576 30580 19582 30592
rect 19613 30583 19671 30589
rect 19613 30580 19625 30583
rect 19576 30552 19625 30580
rect 19576 30540 19582 30552
rect 19613 30549 19625 30552
rect 19659 30549 19671 30583
rect 19613 30543 19671 30549
rect 19705 30583 19763 30589
rect 19705 30549 19717 30583
rect 19751 30580 19763 30583
rect 20717 30583 20775 30589
rect 20717 30580 20729 30583
rect 19751 30552 20729 30580
rect 19751 30549 19763 30552
rect 19705 30543 19763 30549
rect 20717 30549 20729 30552
rect 20763 30549 20775 30583
rect 21008 30580 21036 30688
rect 21082 30676 21088 30728
rect 21140 30716 21146 30728
rect 21545 30719 21603 30725
rect 21545 30716 21557 30719
rect 21140 30688 21557 30716
rect 21140 30676 21146 30688
rect 21545 30685 21557 30688
rect 21591 30685 21603 30719
rect 21545 30679 21603 30685
rect 21735 30657 21763 30756
rect 22281 30753 22293 30756
rect 22327 30784 22339 30787
rect 25682 30784 25688 30796
rect 22327 30756 25688 30784
rect 22327 30753 22339 30756
rect 22281 30747 22339 30753
rect 21913 30719 21971 30725
rect 21913 30685 21925 30719
rect 21959 30716 21971 30719
rect 22002 30716 22008 30728
rect 21959 30688 22008 30716
rect 21959 30685 21971 30688
rect 21913 30679 21971 30685
rect 22002 30676 22008 30688
rect 22060 30716 22066 30728
rect 23293 30719 23351 30725
rect 22060 30688 22692 30716
rect 22060 30676 22066 30688
rect 21729 30651 21787 30657
rect 21729 30617 21741 30651
rect 21775 30617 21787 30651
rect 21729 30611 21787 30617
rect 21818 30608 21824 30660
rect 21876 30648 21882 30660
rect 22462 30648 22468 30660
rect 21876 30620 22468 30648
rect 21876 30608 21882 30620
rect 22462 30608 22468 30620
rect 22520 30608 22526 30660
rect 22557 30651 22615 30657
rect 22557 30617 22569 30651
rect 22603 30617 22615 30651
rect 22664 30648 22692 30688
rect 23293 30685 23305 30719
rect 23339 30716 23351 30719
rect 23382 30716 23388 30728
rect 23339 30688 23388 30716
rect 23339 30685 23351 30688
rect 23293 30679 23351 30685
rect 23382 30676 23388 30688
rect 23440 30676 23446 30728
rect 23492 30725 23520 30756
rect 25682 30744 25688 30756
rect 25740 30744 25746 30796
rect 25774 30744 25780 30796
rect 25832 30744 25838 30796
rect 28258 30744 28264 30796
rect 28316 30744 28322 30796
rect 28718 30744 28724 30796
rect 28776 30784 28782 30796
rect 28997 30787 29055 30793
rect 28997 30784 29009 30787
rect 28776 30756 29009 30784
rect 28776 30744 28782 30756
rect 28997 30753 29009 30756
rect 29043 30753 29055 30787
rect 28997 30747 29055 30753
rect 30193 30787 30251 30793
rect 30193 30753 30205 30787
rect 30239 30784 30251 30787
rect 30282 30784 30288 30796
rect 30239 30756 30288 30784
rect 30239 30753 30251 30756
rect 30193 30747 30251 30753
rect 30282 30744 30288 30756
rect 30340 30744 30346 30796
rect 30926 30744 30932 30796
rect 30984 30744 30990 30796
rect 31202 30744 31208 30796
rect 31260 30784 31266 30796
rect 31297 30787 31355 30793
rect 31297 30784 31309 30787
rect 31260 30756 31309 30784
rect 31260 30744 31266 30756
rect 31297 30753 31309 30756
rect 31343 30753 31355 30787
rect 31297 30747 31355 30753
rect 31754 30744 31760 30796
rect 31812 30784 31818 30796
rect 32033 30787 32091 30793
rect 32033 30784 32045 30787
rect 31812 30756 32045 30784
rect 31812 30744 31818 30756
rect 32033 30753 32045 30756
rect 32079 30753 32091 30787
rect 32140 30784 32168 30824
rect 32140 30756 35020 30784
rect 32033 30747 32091 30753
rect 23477 30719 23535 30725
rect 23477 30685 23489 30719
rect 23523 30685 23535 30719
rect 23477 30679 23535 30685
rect 23566 30676 23572 30728
rect 23624 30676 23630 30728
rect 23661 30719 23719 30725
rect 23661 30685 23673 30719
rect 23707 30716 23719 30719
rect 25314 30716 25320 30728
rect 23707 30688 25320 30716
rect 23707 30685 23719 30688
rect 23661 30679 23719 30685
rect 23676 30648 23704 30679
rect 25314 30676 25320 30688
rect 25372 30676 25378 30728
rect 33410 30676 33416 30728
rect 33468 30676 33474 30728
rect 22664 30620 23704 30648
rect 26053 30651 26111 30657
rect 22557 30611 22615 30617
rect 26053 30617 26065 30651
rect 26099 30617 26111 30651
rect 28626 30648 28632 30660
rect 27278 30620 28632 30648
rect 26053 30611 26111 30617
rect 22002 30580 22008 30592
rect 21008 30552 22008 30580
rect 20717 30543 20775 30549
rect 22002 30540 22008 30552
rect 22060 30540 22066 30592
rect 22370 30540 22376 30592
rect 22428 30580 22434 30592
rect 22572 30580 22600 30611
rect 22428 30552 22600 30580
rect 26068 30580 26096 30611
rect 28626 30608 28632 30620
rect 28684 30608 28690 30660
rect 29917 30651 29975 30657
rect 29917 30617 29929 30651
rect 29963 30648 29975 30651
rect 30098 30648 30104 30660
rect 29963 30620 30104 30648
rect 29963 30617 29975 30620
rect 29917 30611 29975 30617
rect 30098 30608 30104 30620
rect 30156 30608 30162 30660
rect 32306 30608 32312 30660
rect 32364 30608 32370 30660
rect 26234 30580 26240 30592
rect 26068 30552 26240 30580
rect 22428 30540 22434 30552
rect 26234 30540 26240 30552
rect 26292 30540 26298 30592
rect 26786 30540 26792 30592
rect 26844 30580 26850 30592
rect 27525 30583 27583 30589
rect 27525 30580 27537 30583
rect 26844 30552 27537 30580
rect 26844 30540 26850 30552
rect 27525 30549 27537 30552
rect 27571 30549 27583 30583
rect 27525 30543 27583 30549
rect 30009 30583 30067 30589
rect 30009 30549 30021 30583
rect 30055 30580 30067 30583
rect 30377 30583 30435 30589
rect 30377 30580 30389 30583
rect 30055 30552 30389 30580
rect 30055 30549 30067 30552
rect 30009 30543 30067 30549
rect 30377 30549 30389 30552
rect 30423 30549 30435 30583
rect 30377 30543 30435 30549
rect 33134 30540 33140 30592
rect 33192 30580 33198 30592
rect 33781 30583 33839 30589
rect 33781 30580 33793 30583
rect 33192 30552 33793 30580
rect 33192 30540 33198 30552
rect 33781 30549 33793 30552
rect 33827 30549 33839 30583
rect 34992 30580 35020 30756
rect 35710 30744 35716 30796
rect 35768 30744 35774 30796
rect 40678 30784 40684 30796
rect 39960 30756 40684 30784
rect 35066 30676 35072 30728
rect 35124 30716 35130 30728
rect 35437 30719 35495 30725
rect 35437 30716 35449 30719
rect 35124 30688 35449 30716
rect 35124 30676 35130 30688
rect 35437 30685 35449 30688
rect 35483 30685 35495 30719
rect 35437 30679 35495 30685
rect 35526 30676 35532 30728
rect 35584 30676 35590 30728
rect 35805 30719 35863 30725
rect 35805 30685 35817 30719
rect 35851 30716 35863 30719
rect 36814 30716 36820 30728
rect 35851 30688 36820 30716
rect 35851 30685 35863 30688
rect 35805 30679 35863 30685
rect 35342 30608 35348 30660
rect 35400 30648 35406 30660
rect 35820 30648 35848 30679
rect 36814 30676 36820 30688
rect 36872 30716 36878 30728
rect 37734 30716 37740 30728
rect 36872 30688 37740 30716
rect 36872 30676 36878 30688
rect 37734 30676 37740 30688
rect 37792 30676 37798 30728
rect 37829 30719 37887 30725
rect 37829 30685 37841 30719
rect 37875 30716 37887 30719
rect 37918 30716 37924 30728
rect 37875 30688 37924 30716
rect 37875 30685 37887 30688
rect 37829 30679 37887 30685
rect 37918 30676 37924 30688
rect 37976 30676 37982 30728
rect 39960 30725 39988 30756
rect 40678 30744 40684 30756
rect 40736 30744 40742 30796
rect 39853 30719 39911 30725
rect 39853 30716 39865 30719
rect 38028 30688 39865 30716
rect 35400 30620 35848 30648
rect 35400 30608 35406 30620
rect 38028 30580 38056 30688
rect 38304 30660 38332 30688
rect 39853 30685 39865 30688
rect 39899 30685 39911 30719
rect 39853 30679 39911 30685
rect 39945 30719 40003 30725
rect 39945 30685 39957 30719
rect 39991 30685 40003 30719
rect 39945 30679 40003 30685
rect 40126 30676 40132 30728
rect 40184 30676 40190 30728
rect 40402 30676 40408 30728
rect 40460 30676 40466 30728
rect 38096 30651 38154 30657
rect 38096 30617 38108 30651
rect 38142 30648 38154 30651
rect 38194 30648 38200 30660
rect 38142 30620 38200 30648
rect 38142 30617 38154 30620
rect 38096 30611 38154 30617
rect 38194 30608 38200 30620
rect 38252 30608 38258 30660
rect 38286 30608 38292 30660
rect 38344 30608 38350 30660
rect 39868 30620 40448 30648
rect 39868 30592 39896 30620
rect 34992 30552 38056 30580
rect 33781 30543 33839 30549
rect 39850 30540 39856 30592
rect 39908 30540 39914 30592
rect 40310 30540 40316 30592
rect 40368 30540 40374 30592
rect 40420 30580 40448 30620
rect 40678 30608 40684 30660
rect 40736 30608 40742 30660
rect 40788 30620 41170 30648
rect 40788 30580 40816 30620
rect 40420 30552 40816 30580
rect 1104 30490 42504 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 42504 30490
rect 1104 30416 42504 30438
rect 2406 30336 2412 30388
rect 2464 30336 2470 30388
rect 4062 30376 4068 30388
rect 2516 30348 4068 30376
rect 1854 30268 1860 30320
rect 1912 30308 1918 30320
rect 2516 30308 2544 30348
rect 1912 30280 2544 30308
rect 1912 30268 1918 30280
rect 2590 30200 2596 30252
rect 2648 30200 2654 30252
rect 2777 30243 2835 30249
rect 2777 30209 2789 30243
rect 2823 30209 2835 30243
rect 2777 30203 2835 30209
rect 2869 30243 2927 30249
rect 2869 30209 2881 30243
rect 2915 30240 2927 30243
rect 2976 30240 3004 30348
rect 4062 30336 4068 30348
rect 4120 30336 4126 30388
rect 5810 30336 5816 30388
rect 5868 30336 5874 30388
rect 8849 30379 8907 30385
rect 8849 30345 8861 30379
rect 8895 30376 8907 30379
rect 9214 30376 9220 30388
rect 8895 30348 9220 30376
rect 8895 30345 8907 30348
rect 8849 30339 8907 30345
rect 9214 30336 9220 30348
rect 9272 30336 9278 30388
rect 16482 30336 16488 30388
rect 16540 30376 16546 30388
rect 16540 30348 17080 30376
rect 16540 30336 16546 30348
rect 3234 30268 3240 30320
rect 3292 30268 3298 30320
rect 3329 30311 3387 30317
rect 3329 30277 3341 30311
rect 3375 30308 3387 30311
rect 4154 30308 4160 30320
rect 3375 30280 4160 30308
rect 3375 30277 3387 30280
rect 3329 30271 3387 30277
rect 4154 30268 4160 30280
rect 4212 30268 4218 30320
rect 4614 30268 4620 30320
rect 4672 30268 4678 30320
rect 5442 30268 5448 30320
rect 5500 30268 5506 30320
rect 8662 30268 8668 30320
rect 8720 30308 8726 30320
rect 9125 30311 9183 30317
rect 9125 30308 9137 30311
rect 8720 30280 9137 30308
rect 8720 30268 8726 30280
rect 9125 30277 9137 30280
rect 9171 30277 9183 30311
rect 14918 30308 14924 30320
rect 9125 30271 9183 30277
rect 14752 30280 14924 30308
rect 2915 30212 3004 30240
rect 3145 30243 3203 30249
rect 2915 30209 2927 30212
rect 2869 30203 2927 30209
rect 3145 30209 3157 30243
rect 3191 30240 3203 30243
rect 4065 30243 4123 30249
rect 3191 30212 3648 30240
rect 3191 30209 3203 30212
rect 3145 30203 3203 30209
rect 1578 30132 1584 30184
rect 1636 30172 1642 30184
rect 2498 30172 2504 30184
rect 1636 30144 2504 30172
rect 1636 30132 1642 30144
rect 2498 30132 2504 30144
rect 2556 30172 2562 30184
rect 2792 30172 2820 30203
rect 3620 30184 3648 30212
rect 4065 30209 4077 30243
rect 4111 30209 4123 30243
rect 4065 30203 4123 30209
rect 2961 30175 3019 30181
rect 2961 30172 2973 30175
rect 2556 30144 2973 30172
rect 2556 30132 2562 30144
rect 2961 30141 2973 30144
rect 3007 30141 3019 30175
rect 2961 30135 3019 30141
rect 3602 30132 3608 30184
rect 3660 30132 3666 30184
rect 4080 30172 4108 30203
rect 5258 30200 5264 30252
rect 5316 30240 5322 30252
rect 5353 30243 5411 30249
rect 5353 30240 5365 30243
rect 5316 30212 5365 30240
rect 5316 30200 5322 30212
rect 5353 30209 5365 30212
rect 5399 30209 5411 30243
rect 5353 30203 5411 30209
rect 6546 30200 6552 30252
rect 6604 30200 6610 30252
rect 6822 30200 6828 30252
rect 6880 30200 6886 30252
rect 9030 30200 9036 30252
rect 9088 30200 9094 30252
rect 9214 30200 9220 30252
rect 9272 30200 9278 30252
rect 9335 30243 9393 30249
rect 9335 30240 9347 30243
rect 9324 30209 9347 30240
rect 9381 30209 9393 30243
rect 9324 30203 9393 30209
rect 5534 30172 5540 30184
rect 4080 30144 5540 30172
rect 5534 30132 5540 30144
rect 5592 30132 5598 30184
rect 5626 30132 5632 30184
rect 5684 30132 5690 30184
rect 5718 30132 5724 30184
rect 5776 30132 5782 30184
rect 5994 30132 6000 30184
rect 6052 30132 6058 30184
rect 6089 30175 6147 30181
rect 6089 30141 6101 30175
rect 6135 30172 6147 30175
rect 6178 30172 6184 30184
rect 6135 30144 6184 30172
rect 6135 30141 6147 30144
rect 6089 30135 6147 30141
rect 6178 30132 6184 30144
rect 6236 30132 6242 30184
rect 6270 30132 6276 30184
rect 6328 30172 6334 30184
rect 9324 30172 9352 30203
rect 10226 30200 10232 30252
rect 10284 30240 10290 30252
rect 10413 30243 10471 30249
rect 10413 30240 10425 30243
rect 10284 30212 10425 30240
rect 10284 30200 10290 30212
rect 10413 30209 10425 30212
rect 10459 30209 10471 30243
rect 10413 30203 10471 30209
rect 11606 30200 11612 30252
rect 11664 30200 11670 30252
rect 12986 30200 12992 30252
rect 13044 30200 13050 30252
rect 13538 30200 13544 30252
rect 13596 30200 13602 30252
rect 13633 30243 13691 30249
rect 13633 30209 13645 30243
rect 13679 30240 13691 30243
rect 13906 30240 13912 30252
rect 13679 30212 13912 30240
rect 13679 30209 13691 30212
rect 13633 30203 13691 30209
rect 13906 30200 13912 30212
rect 13964 30200 13970 30252
rect 14752 30249 14780 30280
rect 14918 30268 14924 30280
rect 14976 30268 14982 30320
rect 16666 30308 16672 30320
rect 16238 30280 16672 30308
rect 16666 30268 16672 30280
rect 16724 30268 16730 30320
rect 17052 30308 17080 30348
rect 17218 30336 17224 30388
rect 17276 30376 17282 30388
rect 17405 30379 17463 30385
rect 17405 30376 17417 30379
rect 17276 30348 17417 30376
rect 17276 30336 17282 30348
rect 17405 30345 17417 30348
rect 17451 30345 17463 30379
rect 17405 30339 17463 30345
rect 19426 30336 19432 30388
rect 19484 30336 19490 30388
rect 19610 30336 19616 30388
rect 19668 30376 19674 30388
rect 19978 30376 19984 30388
rect 19668 30348 19984 30376
rect 19668 30336 19674 30348
rect 19978 30336 19984 30348
rect 20036 30336 20042 30388
rect 20622 30376 20628 30388
rect 20088 30348 20628 30376
rect 19444 30308 19472 30336
rect 19521 30311 19579 30317
rect 19521 30308 19533 30311
rect 17052 30280 18828 30308
rect 19444 30280 19533 30308
rect 14001 30243 14059 30249
rect 14001 30209 14013 30243
rect 14047 30209 14059 30243
rect 14001 30203 14059 30209
rect 14737 30243 14795 30249
rect 14737 30209 14749 30243
rect 14783 30209 14795 30243
rect 17052 30240 17080 30280
rect 17221 30243 17279 30249
rect 17221 30240 17233 30243
rect 17052 30212 17233 30240
rect 14737 30203 14795 30209
rect 17221 30209 17233 30212
rect 17267 30209 17279 30243
rect 17221 30203 17279 30209
rect 6328 30144 9352 30172
rect 9493 30175 9551 30181
rect 6328 30132 6334 30144
rect 9493 30141 9505 30175
rect 9539 30172 9551 30175
rect 9861 30175 9919 30181
rect 9861 30172 9873 30175
rect 9539 30144 9873 30172
rect 9539 30141 9551 30144
rect 9493 30135 9551 30141
rect 9861 30141 9873 30144
rect 9907 30141 9919 30175
rect 9861 30135 9919 30141
rect 11885 30175 11943 30181
rect 11885 30141 11897 30175
rect 11931 30172 11943 30175
rect 13078 30172 13084 30184
rect 11931 30144 13084 30172
rect 11931 30141 11943 30144
rect 11885 30135 11943 30141
rect 13078 30132 13084 30144
rect 13136 30132 13142 30184
rect 13814 30132 13820 30184
rect 13872 30172 13878 30184
rect 14016 30172 14044 30203
rect 17586 30200 17592 30252
rect 17644 30200 17650 30252
rect 17678 30200 17684 30252
rect 17736 30200 17742 30252
rect 17862 30200 17868 30252
rect 17920 30240 17926 30252
rect 18800 30249 18828 30280
rect 19521 30277 19533 30280
rect 19567 30277 19579 30311
rect 19521 30271 19579 30277
rect 17957 30243 18015 30249
rect 17957 30240 17969 30243
rect 17920 30212 17969 30240
rect 17920 30200 17926 30212
rect 17957 30209 17969 30212
rect 18003 30209 18015 30243
rect 17957 30203 18015 30209
rect 18509 30243 18567 30249
rect 18509 30209 18521 30243
rect 18555 30209 18567 30243
rect 18509 30203 18567 30209
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 13872 30144 14044 30172
rect 15013 30175 15071 30181
rect 13872 30132 13878 30144
rect 15013 30141 15025 30175
rect 15059 30172 15071 30175
rect 16298 30172 16304 30184
rect 15059 30144 16304 30172
rect 15059 30141 15071 30144
rect 15013 30135 15071 30141
rect 16298 30132 16304 30144
rect 16356 30132 16362 30184
rect 17310 30132 17316 30184
rect 17368 30172 17374 30184
rect 18524 30172 18552 30203
rect 19150 30200 19156 30252
rect 19208 30200 19214 30252
rect 19628 30249 19656 30336
rect 19246 30243 19304 30249
rect 19246 30209 19258 30243
rect 19292 30209 19304 30243
rect 19246 30203 19304 30209
rect 19429 30243 19487 30249
rect 19429 30209 19441 30243
rect 19475 30209 19487 30243
rect 19429 30203 19487 30209
rect 19618 30243 19676 30249
rect 19618 30209 19630 30243
rect 19664 30209 19676 30243
rect 19618 30203 19676 30209
rect 17368 30144 18552 30172
rect 17368 30132 17374 30144
rect 19058 30132 19064 30184
rect 19116 30172 19122 30184
rect 19261 30172 19289 30203
rect 19116 30144 19289 30172
rect 19444 30172 19472 30203
rect 19886 30200 19892 30252
rect 19944 30200 19950 30252
rect 20088 30249 20116 30348
rect 20622 30336 20628 30348
rect 20680 30336 20686 30388
rect 21082 30336 21088 30388
rect 21140 30376 21146 30388
rect 21140 30348 22360 30376
rect 21140 30336 21146 30348
rect 20165 30311 20223 30317
rect 20165 30277 20177 30311
rect 20211 30308 20223 30311
rect 20438 30308 20444 30320
rect 20211 30280 20444 30308
rect 20211 30277 20223 30280
rect 20165 30271 20223 30277
rect 20438 30268 20444 30280
rect 20496 30268 20502 30320
rect 21818 30268 21824 30320
rect 21876 30308 21882 30320
rect 22097 30311 22155 30317
rect 22097 30308 22109 30311
rect 21876 30280 22109 30308
rect 21876 30268 21882 30280
rect 22097 30277 22109 30280
rect 22143 30277 22155 30311
rect 22097 30271 22155 30277
rect 20073 30243 20131 30249
rect 20073 30209 20085 30243
rect 20119 30209 20131 30243
rect 20257 30243 20315 30249
rect 20257 30240 20269 30243
rect 20073 30203 20131 30209
rect 20180 30212 20269 30240
rect 20088 30172 20116 30203
rect 20180 30184 20208 30212
rect 20257 30209 20269 30212
rect 20303 30240 20315 30243
rect 20530 30240 20536 30252
rect 20303 30212 20536 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 20530 30200 20536 30212
rect 20588 30200 20594 30252
rect 21266 30200 21272 30252
rect 21324 30200 21330 30252
rect 21361 30243 21419 30249
rect 21361 30209 21373 30243
rect 21407 30209 21419 30243
rect 21361 30203 21419 30209
rect 19444 30144 20116 30172
rect 19116 30132 19122 30144
rect 20162 30132 20168 30184
rect 20220 30132 20226 30184
rect 2590 30064 2596 30116
rect 2648 30104 2654 30116
rect 3234 30104 3240 30116
rect 2648 30076 3240 30104
rect 2648 30064 2654 30076
rect 3234 30064 3240 30076
rect 3292 30064 3298 30116
rect 3513 30107 3571 30113
rect 3513 30073 3525 30107
rect 3559 30104 3571 30107
rect 4614 30104 4620 30116
rect 3559 30076 4620 30104
rect 3559 30073 3571 30076
rect 3513 30067 3571 30073
rect 4614 30064 4620 30076
rect 4672 30104 4678 30116
rect 5166 30104 5172 30116
rect 4672 30076 5172 30104
rect 4672 30064 4678 30076
rect 5166 30064 5172 30076
rect 5224 30064 5230 30116
rect 5442 30064 5448 30116
rect 5500 30104 5506 30116
rect 6641 30107 6699 30113
rect 6641 30104 6653 30107
rect 5500 30076 6653 30104
rect 5500 30064 5506 30076
rect 6641 30073 6653 30076
rect 6687 30073 6699 30107
rect 6641 30067 6699 30073
rect 6733 30107 6791 30113
rect 6733 30073 6745 30107
rect 6779 30073 6791 30107
rect 6733 30067 6791 30073
rect 3878 29996 3884 30048
rect 3936 30036 3942 30048
rect 5810 30036 5816 30048
rect 3936 30008 5816 30036
rect 3936 29996 3942 30008
rect 5810 29996 5816 30008
rect 5868 29996 5874 30048
rect 5902 29996 5908 30048
rect 5960 30036 5966 30048
rect 6365 30039 6423 30045
rect 6365 30036 6377 30039
rect 5960 30008 6377 30036
rect 5960 29996 5966 30008
rect 6365 30005 6377 30008
rect 6411 30005 6423 30039
rect 6365 29999 6423 30005
rect 6454 29996 6460 30048
rect 6512 30036 6518 30048
rect 6748 30036 6776 30067
rect 17034 30064 17040 30116
rect 17092 30104 17098 30116
rect 18690 30104 18696 30116
rect 17092 30076 18696 30104
rect 17092 30064 17098 30076
rect 18690 30064 18696 30076
rect 18748 30064 18754 30116
rect 19794 30064 19800 30116
rect 19852 30064 19858 30116
rect 20441 30107 20499 30113
rect 20441 30073 20453 30107
rect 20487 30104 20499 30107
rect 20806 30104 20812 30116
rect 20487 30076 20812 30104
rect 20487 30073 20499 30076
rect 20441 30067 20499 30073
rect 20806 30064 20812 30076
rect 20864 30064 20870 30116
rect 21376 30104 21404 30203
rect 21634 30200 21640 30252
rect 21692 30200 21698 30252
rect 22002 30249 22008 30252
rect 22000 30240 22008 30249
rect 21963 30212 22008 30240
rect 22000 30203 22008 30212
rect 22002 30200 22008 30203
rect 22060 30200 22066 30252
rect 22186 30200 22192 30252
rect 22244 30200 22250 30252
rect 22332 30249 22360 30348
rect 23014 30336 23020 30388
rect 23072 30376 23078 30388
rect 23072 30348 24348 30376
rect 23072 30336 23078 30348
rect 24320 30308 24348 30348
rect 25682 30336 25688 30388
rect 25740 30376 25746 30388
rect 27798 30376 27804 30388
rect 25740 30348 27804 30376
rect 25740 30336 25746 30348
rect 27798 30336 27804 30348
rect 27856 30336 27862 30388
rect 32306 30336 32312 30388
rect 32364 30376 32370 30388
rect 32493 30379 32551 30385
rect 32493 30376 32505 30379
rect 32364 30348 32505 30376
rect 32364 30336 32370 30348
rect 32493 30345 32505 30348
rect 32539 30345 32551 30379
rect 32493 30339 32551 30345
rect 35066 30336 35072 30388
rect 35124 30336 35130 30388
rect 35434 30336 35440 30388
rect 35492 30376 35498 30388
rect 35529 30379 35587 30385
rect 35529 30376 35541 30379
rect 35492 30348 35541 30376
rect 35492 30336 35498 30348
rect 35529 30345 35541 30348
rect 35575 30345 35587 30379
rect 36354 30376 36360 30388
rect 35529 30339 35587 30345
rect 35723 30348 36360 30376
rect 26142 30308 26148 30320
rect 24242 30280 26148 30308
rect 26142 30268 26148 30280
rect 26200 30268 26206 30320
rect 26234 30268 26240 30320
rect 26292 30268 26298 30320
rect 34698 30317 34704 30320
rect 34685 30311 34704 30317
rect 34685 30277 34697 30311
rect 34685 30271 34704 30277
rect 34698 30268 34704 30271
rect 34756 30268 34762 30320
rect 34885 30311 34943 30317
rect 34885 30277 34897 30311
rect 34931 30308 34943 30311
rect 34931 30280 35572 30308
rect 34931 30277 34943 30280
rect 34885 30271 34943 30277
rect 22317 30243 22375 30249
rect 22317 30209 22329 30243
rect 22363 30209 22375 30243
rect 22317 30203 22375 30209
rect 22462 30200 22468 30252
rect 22520 30200 22526 30252
rect 26421 30243 26479 30249
rect 26421 30209 26433 30243
rect 26467 30209 26479 30243
rect 26421 30203 26479 30209
rect 21542 30132 21548 30184
rect 21600 30172 21606 30184
rect 23201 30175 23259 30181
rect 21600 30144 22232 30172
rect 21600 30132 21606 30144
rect 21821 30107 21879 30113
rect 21821 30104 21833 30107
rect 21008 30076 21312 30104
rect 21376 30076 21833 30104
rect 6512 30008 6776 30036
rect 13357 30039 13415 30045
rect 6512 29996 6518 30008
rect 13357 30005 13369 30039
rect 13403 30036 13415 30039
rect 13998 30036 14004 30048
rect 13403 30008 14004 30036
rect 13403 30005 13415 30008
rect 13357 29999 13415 30005
rect 13998 29996 14004 30008
rect 14056 29996 14062 30048
rect 14185 30039 14243 30045
rect 14185 30005 14197 30039
rect 14231 30036 14243 30039
rect 15378 30036 15384 30048
rect 14231 30008 15384 30036
rect 14231 30005 14243 30008
rect 14185 29999 14243 30005
rect 15378 29996 15384 30008
rect 15436 29996 15442 30048
rect 16669 30039 16727 30045
rect 16669 30005 16681 30039
rect 16715 30036 16727 30039
rect 16758 30036 16764 30048
rect 16715 30008 16764 30036
rect 16715 30005 16727 30008
rect 16669 29999 16727 30005
rect 16758 29996 16764 30008
rect 16816 29996 16822 30048
rect 17126 29996 17132 30048
rect 17184 30036 17190 30048
rect 17865 30039 17923 30045
rect 17865 30036 17877 30039
rect 17184 30008 17877 30036
rect 17184 29996 17190 30008
rect 17865 30005 17877 30008
rect 17911 30036 17923 30039
rect 18230 30036 18236 30048
rect 17911 30008 18236 30036
rect 17911 30005 17923 30008
rect 17865 29999 17923 30005
rect 18230 29996 18236 30008
rect 18288 29996 18294 30048
rect 18322 29996 18328 30048
rect 18380 29996 18386 30048
rect 18414 29996 18420 30048
rect 18472 30036 18478 30048
rect 21008 30036 21036 30076
rect 18472 30008 21036 30036
rect 21085 30039 21143 30045
rect 18472 29996 18478 30008
rect 21085 30005 21097 30039
rect 21131 30036 21143 30039
rect 21174 30036 21180 30048
rect 21131 30008 21180 30036
rect 21131 30005 21143 30008
rect 21085 29999 21143 30005
rect 21174 29996 21180 30008
rect 21232 29996 21238 30048
rect 21284 30036 21312 30076
rect 21821 30073 21833 30076
rect 21867 30073 21879 30107
rect 22204 30104 22232 30144
rect 23201 30141 23213 30175
rect 23247 30172 23259 30175
rect 23290 30172 23296 30184
rect 23247 30144 23296 30172
rect 23247 30141 23259 30144
rect 23201 30135 23259 30141
rect 23290 30132 23296 30144
rect 23348 30132 23354 30184
rect 24578 30132 24584 30184
rect 24636 30172 24642 30184
rect 24673 30175 24731 30181
rect 24673 30172 24685 30175
rect 24636 30144 24685 30172
rect 24636 30132 24642 30144
rect 24673 30141 24685 30144
rect 24719 30141 24731 30175
rect 24673 30135 24731 30141
rect 24949 30175 25007 30181
rect 24949 30141 24961 30175
rect 24995 30141 25007 30175
rect 26436 30172 26464 30203
rect 26510 30200 26516 30252
rect 26568 30200 26574 30252
rect 26786 30200 26792 30252
rect 26844 30200 26850 30252
rect 31665 30243 31723 30249
rect 31665 30209 31677 30243
rect 31711 30240 31723 30243
rect 31754 30240 31760 30252
rect 31711 30212 31760 30240
rect 31711 30209 31723 30212
rect 31665 30203 31723 30209
rect 31754 30200 31760 30212
rect 31812 30200 31818 30252
rect 32677 30243 32735 30249
rect 32677 30209 32689 30243
rect 32723 30209 32735 30243
rect 32677 30203 32735 30209
rect 32769 30243 32827 30249
rect 32769 30209 32781 30243
rect 32815 30240 32827 30243
rect 32950 30240 32956 30252
rect 32815 30212 32956 30240
rect 32815 30209 32827 30212
rect 32769 30203 32827 30209
rect 26602 30172 26608 30184
rect 26436 30144 26608 30172
rect 24949 30135 25007 30141
rect 22204 30076 23704 30104
rect 21821 30067 21879 30073
rect 22462 30036 22468 30048
rect 21284 30008 22468 30036
rect 22462 29996 22468 30008
rect 22520 30036 22526 30048
rect 23198 30036 23204 30048
rect 22520 30008 23204 30036
rect 22520 29996 22526 30008
rect 23198 29996 23204 30008
rect 23256 29996 23262 30048
rect 23676 30036 23704 30076
rect 24486 30036 24492 30048
rect 23676 30008 24492 30036
rect 24486 29996 24492 30008
rect 24544 29996 24550 30048
rect 24670 29996 24676 30048
rect 24728 30036 24734 30048
rect 24964 30036 24992 30135
rect 26602 30132 26608 30144
rect 26660 30132 26666 30184
rect 32692 30172 32720 30203
rect 32950 30200 32956 30212
rect 33008 30200 33014 30252
rect 33045 30243 33103 30249
rect 33045 30209 33057 30243
rect 33091 30240 33103 30243
rect 33134 30240 33140 30252
rect 33091 30212 33140 30240
rect 33091 30209 33103 30212
rect 33045 30203 33103 30209
rect 33134 30200 33140 30212
rect 33192 30200 33198 30252
rect 34330 30200 34336 30252
rect 34388 30240 34394 30252
rect 34977 30243 35035 30249
rect 34977 30240 34989 30243
rect 34388 30212 34989 30240
rect 34388 30200 34394 30212
rect 34977 30209 34989 30212
rect 35023 30209 35035 30243
rect 34977 30203 35035 30209
rect 35161 30243 35219 30249
rect 35161 30209 35173 30243
rect 35207 30209 35219 30243
rect 35161 30203 35219 30209
rect 33686 30172 33692 30184
rect 32692 30144 33692 30172
rect 33686 30132 33692 30144
rect 33744 30132 33750 30184
rect 34606 30132 34612 30184
rect 34664 30172 34670 30184
rect 35176 30172 35204 30203
rect 34664 30144 35204 30172
rect 34664 30132 34670 30144
rect 26050 30064 26056 30116
rect 26108 30104 26114 30116
rect 30466 30104 30472 30116
rect 26108 30076 30472 30104
rect 26108 30064 26114 30076
rect 30466 30064 30472 30076
rect 30524 30064 30530 30116
rect 33962 30064 33968 30116
rect 34020 30104 34026 30116
rect 35544 30104 35572 30280
rect 35723 30249 35751 30348
rect 36354 30336 36360 30348
rect 36412 30376 36418 30388
rect 37550 30376 37556 30388
rect 36412 30348 37556 30376
rect 36412 30336 36418 30348
rect 37550 30336 37556 30348
rect 37608 30336 37614 30388
rect 38194 30336 38200 30388
rect 38252 30336 38258 30388
rect 40034 30336 40040 30388
rect 40092 30376 40098 30388
rect 40129 30379 40187 30385
rect 40129 30376 40141 30379
rect 40092 30348 40141 30376
rect 40092 30336 40098 30348
rect 40129 30345 40141 30348
rect 40175 30345 40187 30379
rect 40129 30339 40187 30345
rect 40494 30336 40500 30388
rect 40552 30336 40558 30388
rect 40954 30336 40960 30388
rect 41012 30336 41018 30388
rect 41230 30336 41236 30388
rect 41288 30376 41294 30388
rect 41417 30379 41475 30385
rect 41417 30376 41429 30379
rect 41288 30348 41429 30376
rect 41288 30336 41294 30348
rect 41417 30345 41429 30348
rect 41463 30345 41475 30379
rect 41417 30339 41475 30345
rect 35805 30311 35863 30317
rect 35805 30277 35817 30311
rect 35851 30308 35863 30311
rect 36722 30308 36728 30320
rect 35851 30280 36728 30308
rect 35851 30277 35863 30280
rect 35805 30271 35863 30277
rect 36722 30268 36728 30280
rect 36780 30268 36786 30320
rect 37918 30308 37924 30320
rect 37476 30280 37924 30308
rect 35708 30243 35766 30249
rect 35708 30209 35720 30243
rect 35754 30209 35766 30243
rect 35897 30243 35955 30249
rect 35897 30240 35909 30243
rect 35708 30203 35766 30209
rect 35821 30212 35909 30240
rect 35821 30184 35849 30212
rect 35897 30209 35909 30212
rect 35943 30209 35955 30243
rect 35897 30203 35955 30209
rect 35986 30200 35992 30252
rect 36044 30249 36050 30252
rect 36044 30243 36083 30249
rect 36071 30209 36083 30243
rect 36044 30203 36083 30209
rect 36044 30200 36050 30203
rect 36170 30200 36176 30252
rect 36228 30200 36234 30252
rect 36262 30200 36268 30252
rect 36320 30200 36326 30252
rect 36446 30200 36452 30252
rect 36504 30200 36510 30252
rect 36538 30200 36544 30252
rect 36596 30200 36602 30252
rect 36630 30200 36636 30252
rect 36688 30200 36694 30252
rect 37277 30243 37335 30249
rect 37277 30240 37289 30243
rect 36832 30212 37289 30240
rect 35802 30132 35808 30184
rect 35860 30132 35866 30184
rect 36832 30113 36860 30212
rect 37277 30209 37289 30212
rect 37323 30209 37335 30243
rect 37277 30203 37335 30209
rect 37366 30200 37372 30252
rect 37424 30249 37430 30252
rect 37476 30249 37504 30280
rect 37918 30268 37924 30280
rect 37976 30268 37982 30320
rect 38654 30308 38660 30320
rect 38028 30280 38660 30308
rect 37424 30243 37504 30249
rect 37424 30209 37437 30243
rect 37471 30212 37504 30243
rect 37471 30209 37483 30212
rect 37424 30203 37483 30209
rect 37424 30200 37430 30203
rect 37550 30200 37556 30252
rect 37608 30200 37614 30252
rect 37826 30249 37832 30252
rect 37645 30243 37703 30249
rect 37645 30209 37657 30243
rect 37691 30209 37703 30243
rect 37645 30203 37703 30209
rect 37783 30243 37832 30249
rect 37783 30209 37795 30243
rect 37829 30209 37832 30243
rect 37783 30203 37832 30209
rect 37660 30172 37688 30203
rect 37826 30200 37832 30203
rect 37884 30200 37890 30252
rect 38028 30172 38056 30280
rect 38654 30268 38660 30280
rect 38712 30268 38718 30320
rect 38746 30268 38752 30320
rect 38804 30308 38810 30320
rect 39114 30308 39120 30320
rect 38804 30280 39120 30308
rect 38804 30268 38810 30280
rect 39114 30268 39120 30280
rect 39172 30268 39178 30320
rect 39942 30268 39948 30320
rect 40000 30308 40006 30320
rect 40589 30311 40647 30317
rect 40589 30308 40601 30311
rect 40000 30280 40601 30308
rect 40000 30268 40006 30280
rect 40589 30277 40601 30280
rect 40635 30277 40647 30311
rect 40589 30271 40647 30277
rect 38378 30200 38384 30252
rect 38436 30240 38442 30252
rect 38565 30243 38623 30249
rect 38565 30240 38577 30243
rect 38436 30212 38577 30240
rect 38436 30200 38442 30212
rect 38565 30209 38577 30212
rect 38611 30209 38623 30243
rect 38672 30240 38700 30268
rect 39758 30240 39764 30252
rect 38672 30212 39764 30240
rect 38565 30203 38623 30209
rect 39758 30200 39764 30212
rect 39816 30200 39822 30252
rect 41325 30243 41383 30249
rect 41325 30240 41337 30243
rect 39868 30212 41337 30240
rect 37660 30144 38056 30172
rect 38654 30132 38660 30184
rect 38712 30132 38718 30184
rect 38841 30175 38899 30181
rect 38841 30141 38853 30175
rect 38887 30172 38899 30175
rect 38930 30172 38936 30184
rect 38887 30144 38936 30172
rect 38887 30141 38899 30144
rect 38841 30135 38899 30141
rect 38930 30132 38936 30144
rect 38988 30132 38994 30184
rect 39022 30132 39028 30184
rect 39080 30172 39086 30184
rect 39868 30172 39896 30212
rect 41325 30209 41337 30212
rect 41371 30209 41383 30243
rect 41325 30203 41383 30209
rect 41782 30200 41788 30252
rect 41840 30200 41846 30252
rect 39080 30144 39896 30172
rect 39945 30175 40003 30181
rect 39080 30132 39086 30144
rect 39945 30141 39957 30175
rect 39991 30172 40003 30175
rect 40402 30172 40408 30184
rect 39991 30144 40408 30172
rect 39991 30141 40003 30144
rect 39945 30135 40003 30141
rect 40402 30132 40408 30144
rect 40460 30132 40466 30184
rect 40586 30132 40592 30184
rect 40644 30172 40650 30184
rect 40681 30175 40739 30181
rect 40681 30172 40693 30175
rect 40644 30144 40693 30172
rect 40644 30132 40650 30144
rect 40681 30141 40693 30144
rect 40727 30172 40739 30175
rect 41509 30175 41567 30181
rect 41509 30172 41521 30175
rect 40727 30144 41521 30172
rect 40727 30141 40739 30144
rect 40681 30135 40739 30141
rect 41509 30141 41521 30144
rect 41555 30141 41567 30175
rect 41509 30135 41567 30141
rect 36817 30107 36875 30113
rect 34020 30076 34928 30104
rect 35544 30076 36584 30104
rect 34020 30064 34026 30076
rect 24728 30008 24992 30036
rect 24728 29996 24734 30008
rect 26142 29996 26148 30048
rect 26200 30036 26206 30048
rect 26697 30039 26755 30045
rect 26697 30036 26709 30039
rect 26200 30008 26709 30036
rect 26200 29996 26206 30008
rect 26697 30005 26709 30008
rect 26743 30036 26755 30039
rect 32953 30039 33011 30045
rect 32953 30036 32965 30039
rect 26743 30008 32965 30036
rect 26743 30005 26755 30008
rect 26697 29999 26755 30005
rect 32953 30005 32965 30008
rect 32999 30005 33011 30039
rect 32953 29999 33011 30005
rect 34422 29996 34428 30048
rect 34480 30036 34486 30048
rect 34517 30039 34575 30045
rect 34517 30036 34529 30039
rect 34480 30008 34529 30036
rect 34480 29996 34486 30008
rect 34517 30005 34529 30008
rect 34563 30005 34575 30039
rect 34517 29999 34575 30005
rect 34701 30039 34759 30045
rect 34701 30005 34713 30039
rect 34747 30036 34759 30039
rect 34790 30036 34796 30048
rect 34747 30008 34796 30036
rect 34747 30005 34759 30008
rect 34701 29999 34759 30005
rect 34790 29996 34796 30008
rect 34848 29996 34854 30048
rect 34900 30036 34928 30076
rect 36556 30048 36584 30076
rect 36817 30073 36829 30107
rect 36863 30073 36875 30107
rect 39040 30104 39068 30132
rect 36817 30067 36875 30073
rect 36924 30076 39068 30104
rect 35618 30036 35624 30048
rect 34900 30008 35624 30036
rect 35618 29996 35624 30008
rect 35676 29996 35682 30048
rect 35894 29996 35900 30048
rect 35952 30036 35958 30048
rect 36262 30036 36268 30048
rect 35952 30008 36268 30036
rect 35952 29996 35958 30008
rect 36262 29996 36268 30008
rect 36320 29996 36326 30048
rect 36538 29996 36544 30048
rect 36596 30036 36602 30048
rect 36924 30036 36952 30076
rect 36596 30008 36952 30036
rect 37921 30039 37979 30045
rect 36596 29996 36602 30008
rect 37921 30005 37933 30039
rect 37967 30036 37979 30039
rect 40034 30036 40040 30048
rect 37967 30008 40040 30036
rect 37967 30005 37979 30008
rect 37921 29999 37979 30005
rect 40034 29996 40040 30008
rect 40092 29996 40098 30048
rect 41966 29996 41972 30048
rect 42024 29996 42030 30048
rect 1104 29946 42504 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 42504 29946
rect 1104 29872 42504 29894
rect 5353 29835 5411 29841
rect 3436 29804 4384 29832
rect 3436 29776 3464 29804
rect 3418 29724 3424 29776
rect 3476 29724 3482 29776
rect 3602 29724 3608 29776
rect 3660 29764 3666 29776
rect 3660 29736 4200 29764
rect 3660 29724 3666 29736
rect 3436 29696 3464 29724
rect 4172 29705 4200 29736
rect 4065 29699 4123 29705
rect 4065 29696 4077 29699
rect 3436 29668 4077 29696
rect 4065 29665 4077 29668
rect 4111 29665 4123 29699
rect 4065 29659 4123 29665
rect 4157 29699 4215 29705
rect 4157 29665 4169 29699
rect 4203 29665 4215 29699
rect 4157 29659 4215 29665
rect 4356 29640 4384 29804
rect 5353 29801 5365 29835
rect 5399 29832 5411 29835
rect 5626 29832 5632 29844
rect 5399 29804 5632 29832
rect 5399 29801 5411 29804
rect 5353 29795 5411 29801
rect 5626 29792 5632 29804
rect 5684 29792 5690 29844
rect 9030 29792 9036 29844
rect 9088 29832 9094 29844
rect 9585 29835 9643 29841
rect 9585 29832 9597 29835
rect 9088 29804 9597 29832
rect 9088 29792 9094 29804
rect 9585 29801 9597 29804
rect 9631 29801 9643 29835
rect 9585 29795 9643 29801
rect 13078 29792 13084 29844
rect 13136 29792 13142 29844
rect 16298 29792 16304 29844
rect 16356 29792 16362 29844
rect 17586 29832 17592 29844
rect 16500 29804 17592 29832
rect 5718 29764 5724 29776
rect 4908 29736 5724 29764
rect 4430 29656 4436 29708
rect 4488 29696 4494 29708
rect 4908 29696 4936 29736
rect 5718 29724 5724 29736
rect 5776 29724 5782 29776
rect 6086 29764 6092 29776
rect 5828 29736 6092 29764
rect 5828 29696 5856 29736
rect 6086 29724 6092 29736
rect 6144 29764 6150 29776
rect 6546 29764 6552 29776
rect 6144 29736 6552 29764
rect 6144 29724 6150 29736
rect 6546 29724 6552 29736
rect 6604 29724 6610 29776
rect 10962 29764 10968 29776
rect 8036 29736 10968 29764
rect 4488 29668 4936 29696
rect 4488 29656 4494 29668
rect 1762 29588 1768 29640
rect 1820 29628 1826 29640
rect 2777 29631 2835 29637
rect 2777 29628 2789 29631
rect 1820 29600 2789 29628
rect 1820 29588 1826 29600
rect 2777 29597 2789 29600
rect 2823 29628 2835 29631
rect 2866 29628 2872 29640
rect 2823 29600 2872 29628
rect 2823 29597 2835 29600
rect 2777 29591 2835 29597
rect 2866 29588 2872 29600
rect 2924 29588 2930 29640
rect 3050 29588 3056 29640
rect 3108 29588 3114 29640
rect 3421 29631 3479 29637
rect 3421 29597 3433 29631
rect 3467 29628 3479 29631
rect 3694 29628 3700 29640
rect 3467 29600 3700 29628
rect 3467 29597 3479 29600
rect 3421 29591 3479 29597
rect 3694 29588 3700 29600
rect 3752 29588 3758 29640
rect 3786 29588 3792 29640
rect 3844 29628 3850 29640
rect 3970 29628 3976 29640
rect 3844 29600 3976 29628
rect 3844 29588 3850 29600
rect 3970 29588 3976 29600
rect 4028 29588 4034 29640
rect 4249 29631 4307 29637
rect 4249 29597 4261 29631
rect 4295 29597 4307 29631
rect 4249 29591 4307 29597
rect 1946 29520 1952 29572
rect 2004 29560 2010 29572
rect 2593 29563 2651 29569
rect 2593 29560 2605 29563
rect 2004 29532 2605 29560
rect 2004 29520 2010 29532
rect 2593 29529 2605 29532
rect 2639 29560 2651 29563
rect 2639 29532 3096 29560
rect 2639 29529 2651 29532
rect 2593 29523 2651 29529
rect 2406 29452 2412 29504
rect 2464 29452 2470 29504
rect 2866 29452 2872 29504
rect 2924 29452 2930 29504
rect 3068 29492 3096 29532
rect 3142 29520 3148 29572
rect 3200 29520 3206 29572
rect 3237 29563 3295 29569
rect 3237 29529 3249 29563
rect 3283 29560 3295 29563
rect 3878 29560 3884 29572
rect 3283 29532 3884 29560
rect 3283 29529 3295 29532
rect 3237 29523 3295 29529
rect 3878 29520 3884 29532
rect 3936 29560 3942 29572
rect 4264 29560 4292 29591
rect 4338 29588 4344 29640
rect 4396 29628 4402 29640
rect 4908 29637 4936 29668
rect 5736 29668 5856 29696
rect 4709 29631 4767 29637
rect 4709 29628 4721 29631
rect 4396 29600 4721 29628
rect 4396 29588 4402 29600
rect 4709 29597 4721 29600
rect 4755 29597 4767 29631
rect 4709 29591 4767 29597
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29597 4951 29631
rect 4893 29591 4951 29597
rect 4985 29631 5043 29637
rect 4985 29597 4997 29631
rect 5031 29597 5043 29631
rect 4985 29591 5043 29597
rect 5077 29631 5135 29637
rect 5077 29597 5089 29631
rect 5123 29628 5135 29631
rect 5442 29628 5448 29640
rect 5123 29600 5448 29628
rect 5123 29597 5135 29600
rect 5077 29591 5135 29597
rect 3936 29532 4292 29560
rect 3936 29520 3942 29532
rect 4798 29520 4804 29572
rect 4856 29560 4862 29572
rect 5000 29560 5028 29591
rect 5442 29588 5448 29600
rect 5500 29588 5506 29640
rect 5626 29588 5632 29640
rect 5684 29588 5690 29640
rect 5736 29637 5764 29668
rect 5902 29656 5908 29708
rect 5960 29656 5966 29708
rect 6365 29699 6423 29705
rect 6365 29665 6377 29699
rect 6411 29696 6423 29699
rect 6454 29696 6460 29708
rect 6411 29668 6460 29696
rect 6411 29665 6423 29668
rect 6365 29659 6423 29665
rect 6454 29656 6460 29668
rect 6512 29656 6518 29708
rect 6638 29656 6644 29708
rect 6696 29656 6702 29708
rect 5721 29631 5779 29637
rect 5721 29597 5733 29631
rect 5767 29597 5779 29631
rect 5721 29591 5779 29597
rect 5810 29588 5816 29640
rect 5868 29628 5874 29640
rect 6273 29631 6331 29637
rect 6273 29628 6285 29631
rect 5868 29600 6285 29628
rect 5868 29588 5874 29600
rect 6273 29597 6285 29600
rect 6319 29597 6331 29631
rect 8036 29614 8064 29736
rect 10962 29724 10968 29736
rect 11020 29724 11026 29776
rect 12989 29767 13047 29773
rect 12989 29733 13001 29767
rect 13035 29764 13047 29767
rect 13538 29764 13544 29776
rect 13035 29736 13544 29764
rect 13035 29733 13047 29736
rect 12989 29727 13047 29733
rect 13538 29724 13544 29736
rect 13596 29724 13602 29776
rect 10226 29696 10232 29708
rect 9784 29668 10232 29696
rect 9784 29637 9812 29668
rect 10226 29656 10232 29668
rect 10284 29656 10290 29708
rect 11241 29699 11299 29705
rect 11241 29665 11253 29699
rect 11287 29696 11299 29699
rect 11606 29696 11612 29708
rect 11287 29668 11612 29696
rect 11287 29665 11299 29668
rect 11241 29659 11299 29665
rect 11606 29656 11612 29668
rect 11664 29656 11670 29708
rect 13998 29656 14004 29708
rect 14056 29696 14062 29708
rect 14645 29699 14703 29705
rect 14645 29696 14657 29699
rect 14056 29668 14657 29696
rect 14056 29656 14062 29668
rect 14645 29665 14657 29668
rect 14691 29696 14703 29699
rect 14829 29699 14887 29705
rect 14829 29696 14841 29699
rect 14691 29668 14841 29696
rect 14691 29665 14703 29668
rect 14645 29659 14703 29665
rect 14829 29665 14841 29668
rect 14875 29665 14887 29699
rect 14829 29659 14887 29665
rect 9769 29631 9827 29637
rect 6273 29591 6331 29597
rect 9769 29597 9781 29631
rect 9815 29597 9827 29631
rect 10045 29631 10103 29637
rect 10045 29628 10057 29631
rect 9769 29591 9827 29597
rect 9876 29600 10057 29628
rect 4856 29532 5028 29560
rect 6549 29563 6607 29569
rect 4856 29520 4862 29532
rect 6549 29529 6561 29563
rect 6595 29560 6607 29563
rect 6917 29563 6975 29569
rect 6917 29560 6929 29563
rect 6595 29532 6929 29560
rect 6595 29529 6607 29532
rect 6549 29523 6607 29529
rect 6917 29529 6929 29532
rect 6963 29529 6975 29563
rect 6917 29523 6975 29529
rect 3602 29492 3608 29504
rect 3068 29464 3608 29492
rect 3602 29452 3608 29464
rect 3660 29452 3666 29504
rect 3786 29452 3792 29504
rect 3844 29452 3850 29504
rect 3970 29452 3976 29504
rect 4028 29492 4034 29504
rect 5537 29495 5595 29501
rect 5537 29492 5549 29495
rect 4028 29464 5549 29492
rect 4028 29452 4034 29464
rect 5537 29461 5549 29464
rect 5583 29492 5595 29495
rect 5718 29492 5724 29504
rect 5583 29464 5724 29492
rect 5583 29461 5595 29464
rect 5537 29455 5595 29461
rect 5718 29452 5724 29464
rect 5776 29452 5782 29504
rect 8202 29452 8208 29504
rect 8260 29492 8266 29504
rect 8389 29495 8447 29501
rect 8389 29492 8401 29495
rect 8260 29464 8401 29492
rect 8260 29452 8266 29464
rect 8389 29461 8401 29464
rect 8435 29492 8447 29495
rect 9876 29492 9904 29600
rect 10045 29597 10057 29600
rect 10091 29597 10103 29631
rect 10045 29591 10103 29597
rect 13262 29588 13268 29640
rect 13320 29588 13326 29640
rect 13357 29631 13415 29637
rect 13357 29597 13369 29631
rect 13403 29628 13415 29631
rect 14093 29631 14151 29637
rect 14093 29628 14105 29631
rect 13403 29600 14105 29628
rect 13403 29597 13415 29600
rect 13357 29591 13415 29597
rect 14093 29597 14105 29600
rect 14139 29597 14151 29631
rect 14093 29591 14151 29597
rect 15194 29588 15200 29640
rect 15252 29588 15258 29640
rect 16500 29637 16528 29804
rect 17586 29792 17592 29804
rect 17644 29792 17650 29844
rect 19150 29792 19156 29844
rect 19208 29832 19214 29844
rect 19245 29835 19303 29841
rect 19245 29832 19257 29835
rect 19208 29804 19257 29832
rect 19208 29792 19214 29804
rect 19245 29801 19257 29804
rect 19291 29801 19303 29835
rect 19245 29795 19303 29801
rect 19702 29792 19708 29844
rect 19760 29792 19766 29844
rect 21174 29841 21180 29844
rect 19889 29835 19947 29841
rect 19889 29801 19901 29835
rect 19935 29801 19947 29835
rect 19889 29795 19947 29801
rect 21164 29835 21180 29841
rect 21164 29801 21176 29835
rect 21164 29795 21180 29801
rect 16577 29767 16635 29773
rect 16577 29733 16589 29767
rect 16623 29764 16635 29767
rect 18322 29764 18328 29776
rect 16623 29736 18328 29764
rect 16623 29733 16635 29736
rect 16577 29727 16635 29733
rect 18322 29724 18328 29736
rect 18380 29724 18386 29776
rect 19061 29767 19119 29773
rect 19061 29733 19073 29767
rect 19107 29764 19119 29767
rect 19904 29764 19932 29795
rect 21174 29792 21180 29795
rect 21232 29792 21238 29844
rect 21818 29792 21824 29844
rect 21876 29832 21882 29844
rect 21876 29804 22232 29832
rect 21876 29792 21882 29804
rect 19107 29736 19932 29764
rect 22204 29764 22232 29804
rect 22462 29792 22468 29844
rect 22520 29832 22526 29844
rect 22649 29835 22707 29841
rect 22649 29832 22661 29835
rect 22520 29804 22661 29832
rect 22520 29792 22526 29804
rect 22649 29801 22661 29804
rect 22695 29801 22707 29835
rect 22649 29795 22707 29801
rect 22756 29804 24532 29832
rect 22756 29764 22784 29804
rect 23842 29764 23848 29776
rect 22204 29736 22784 29764
rect 23400 29736 23848 29764
rect 19107 29733 19119 29736
rect 19061 29727 19119 29733
rect 16758 29656 16764 29708
rect 16816 29656 16822 29708
rect 16850 29656 16856 29708
rect 16908 29696 16914 29708
rect 17129 29699 17187 29705
rect 17129 29696 17141 29699
rect 16908 29668 17141 29696
rect 16908 29656 16914 29668
rect 17129 29665 17141 29668
rect 17175 29696 17187 29699
rect 18049 29699 18107 29705
rect 18049 29696 18061 29699
rect 17175 29668 18061 29696
rect 17175 29665 17187 29668
rect 17129 29659 17187 29665
rect 18049 29665 18061 29668
rect 18095 29665 18107 29699
rect 18049 29659 18107 29665
rect 18230 29656 18236 29708
rect 18288 29696 18294 29708
rect 19794 29696 19800 29708
rect 18288 29668 19800 29696
rect 18288 29656 18294 29668
rect 16485 29631 16543 29637
rect 16485 29597 16497 29631
rect 16531 29597 16543 29631
rect 16485 29591 16543 29597
rect 16669 29631 16727 29637
rect 16669 29597 16681 29631
rect 16715 29597 16727 29631
rect 16669 29591 16727 29597
rect 9953 29563 10011 29569
rect 9953 29529 9965 29563
rect 9999 29560 10011 29563
rect 10410 29560 10416 29572
rect 9999 29532 10416 29560
rect 9999 29529 10011 29532
rect 9953 29523 10011 29529
rect 10410 29520 10416 29532
rect 10468 29520 10474 29572
rect 11517 29563 11575 29569
rect 11517 29529 11529 29563
rect 11563 29560 11575 29563
rect 11790 29560 11796 29572
rect 11563 29532 11796 29560
rect 11563 29529 11575 29532
rect 11517 29523 11575 29529
rect 11790 29520 11796 29532
rect 11848 29520 11854 29572
rect 12986 29560 12992 29572
rect 12742 29532 12992 29560
rect 12986 29520 12992 29532
rect 13044 29560 13050 29572
rect 13044 29532 13860 29560
rect 13044 29520 13050 29532
rect 8435 29464 9904 29492
rect 8435 29461 8447 29464
rect 8389 29455 8447 29461
rect 13538 29452 13544 29504
rect 13596 29492 13602 29504
rect 13725 29495 13783 29501
rect 13725 29492 13737 29495
rect 13596 29464 13737 29492
rect 13596 29452 13602 29464
rect 13725 29461 13737 29464
rect 13771 29461 13783 29495
rect 13832 29492 13860 29532
rect 13906 29520 13912 29572
rect 13964 29560 13970 29572
rect 15105 29563 15163 29569
rect 15105 29560 15117 29563
rect 13964 29532 15117 29560
rect 13964 29520 13970 29532
rect 15105 29529 15117 29532
rect 15151 29529 15163 29563
rect 16684 29560 16712 29591
rect 16942 29588 16948 29640
rect 17000 29588 17006 29640
rect 17313 29631 17371 29637
rect 17313 29597 17325 29631
rect 17359 29628 17371 29631
rect 17402 29628 17408 29640
rect 17359 29600 17408 29628
rect 17359 29597 17371 29600
rect 17313 29591 17371 29597
rect 17402 29588 17408 29600
rect 17460 29628 17466 29640
rect 17862 29628 17868 29640
rect 17460 29600 17868 29628
rect 17460 29588 17466 29600
rect 17862 29588 17868 29600
rect 17920 29628 17926 29640
rect 18325 29631 18383 29637
rect 17920 29600 18092 29628
rect 17920 29588 17926 29600
rect 17954 29560 17960 29572
rect 16684 29532 17960 29560
rect 15105 29523 15163 29529
rect 17954 29520 17960 29532
rect 18012 29520 18018 29572
rect 14734 29492 14740 29504
rect 13832 29464 14740 29492
rect 13725 29455 13783 29461
rect 14734 29452 14740 29464
rect 14792 29492 14798 29504
rect 15013 29495 15071 29501
rect 15013 29492 15025 29495
rect 14792 29464 15025 29492
rect 14792 29452 14798 29464
rect 15013 29461 15025 29464
rect 15059 29461 15071 29495
rect 15013 29455 15071 29461
rect 15381 29495 15439 29501
rect 15381 29461 15393 29495
rect 15427 29492 15439 29495
rect 16206 29492 16212 29504
rect 15427 29464 16212 29492
rect 15427 29461 15439 29464
rect 15381 29455 15439 29461
rect 16206 29452 16212 29464
rect 16264 29452 16270 29504
rect 17218 29452 17224 29504
rect 17276 29492 17282 29504
rect 17405 29495 17463 29501
rect 17405 29492 17417 29495
rect 17276 29464 17417 29492
rect 17276 29452 17282 29464
rect 17405 29461 17417 29464
rect 17451 29492 17463 29495
rect 17586 29492 17592 29504
rect 17451 29464 17592 29492
rect 17451 29461 17463 29464
rect 17405 29455 17463 29461
rect 17586 29452 17592 29464
rect 17644 29452 17650 29504
rect 17770 29452 17776 29504
rect 17828 29452 17834 29504
rect 18064 29492 18092 29600
rect 18325 29597 18337 29631
rect 18371 29628 18383 29631
rect 18414 29628 18420 29640
rect 18371 29600 18420 29628
rect 18371 29597 18383 29600
rect 18325 29591 18383 29597
rect 18414 29588 18420 29600
rect 18472 29588 18478 29640
rect 18509 29631 18567 29637
rect 18509 29597 18521 29631
rect 18555 29628 18567 29631
rect 18598 29628 18604 29640
rect 18555 29600 18604 29628
rect 18555 29597 18567 29600
rect 18509 29591 18567 29597
rect 18598 29588 18604 29600
rect 18656 29588 18662 29640
rect 18892 29637 18920 29668
rect 19794 29656 19800 29668
rect 19852 29656 19858 29708
rect 20901 29699 20959 29705
rect 20901 29665 20913 29699
rect 20947 29696 20959 29699
rect 23400 29696 23428 29736
rect 23842 29724 23848 29736
rect 23900 29724 23906 29776
rect 23937 29767 23995 29773
rect 23937 29733 23949 29767
rect 23983 29733 23995 29767
rect 24504 29764 24532 29804
rect 24578 29792 24584 29844
rect 24636 29832 24642 29844
rect 24949 29835 25007 29841
rect 24949 29832 24961 29835
rect 24636 29804 24961 29832
rect 24636 29792 24642 29804
rect 24949 29801 24961 29804
rect 24995 29801 25007 29835
rect 26145 29835 26203 29841
rect 24949 29795 25007 29801
rect 25056 29804 26096 29832
rect 25056 29764 25084 29804
rect 24504 29736 25084 29764
rect 23937 29727 23995 29733
rect 20947 29668 23428 29696
rect 23952 29696 23980 29727
rect 25222 29724 25228 29776
rect 25280 29764 25286 29776
rect 26068 29764 26096 29804
rect 26145 29801 26157 29835
rect 26191 29832 26203 29835
rect 26510 29832 26516 29844
rect 26191 29804 26516 29832
rect 26191 29801 26203 29804
rect 26145 29795 26203 29801
rect 26510 29792 26516 29804
rect 26568 29792 26574 29844
rect 26602 29792 26608 29844
rect 26660 29832 26666 29844
rect 26789 29835 26847 29841
rect 26789 29832 26801 29835
rect 26660 29804 26801 29832
rect 26660 29792 26666 29804
rect 26789 29801 26801 29804
rect 26835 29801 26847 29835
rect 26789 29795 26847 29801
rect 29273 29835 29331 29841
rect 29273 29801 29285 29835
rect 29319 29832 29331 29835
rect 30009 29835 30067 29841
rect 30009 29832 30021 29835
rect 29319 29804 30021 29832
rect 29319 29801 29331 29804
rect 29273 29795 29331 29801
rect 30009 29801 30021 29804
rect 30055 29832 30067 29835
rect 32582 29832 32588 29844
rect 30055 29804 32588 29832
rect 30055 29801 30067 29804
rect 30009 29795 30067 29801
rect 32582 29792 32588 29804
rect 32640 29792 32646 29844
rect 32950 29792 32956 29844
rect 33008 29792 33014 29844
rect 33134 29832 33140 29844
rect 33051 29804 33140 29832
rect 31478 29764 31484 29776
rect 25280 29736 25912 29764
rect 26068 29736 31484 29764
rect 25280 29724 25286 29736
rect 23952 29668 24072 29696
rect 20947 29665 20959 29668
rect 20901 29659 20959 29665
rect 18877 29631 18935 29637
rect 18877 29597 18889 29631
rect 18923 29597 18935 29631
rect 18877 29591 18935 29597
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29628 19487 29631
rect 19518 29628 19524 29640
rect 19475 29600 19524 29628
rect 19475 29597 19487 29600
rect 19429 29591 19487 29597
rect 19518 29588 19524 29600
rect 19576 29588 19582 29640
rect 19613 29631 19671 29637
rect 19613 29597 19625 29631
rect 19659 29628 19671 29631
rect 20070 29628 20076 29640
rect 19659 29600 20076 29628
rect 19659 29597 19671 29600
rect 19613 29591 19671 29597
rect 20070 29588 20076 29600
rect 20128 29628 20134 29640
rect 20128 29600 20208 29628
rect 20128 29588 20134 29600
rect 18690 29520 18696 29572
rect 18748 29520 18754 29572
rect 18785 29563 18843 29569
rect 18785 29529 18797 29563
rect 18831 29529 18843 29563
rect 20180 29560 20208 29600
rect 20254 29588 20260 29640
rect 20312 29588 20318 29640
rect 20625 29631 20683 29637
rect 20625 29597 20637 29631
rect 20671 29628 20683 29631
rect 20714 29628 20720 29640
rect 20671 29600 20720 29628
rect 20671 29597 20683 29600
rect 20625 29591 20683 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 23014 29628 23020 29640
rect 22310 29600 23020 29628
rect 23014 29588 23020 29600
rect 23072 29588 23078 29640
rect 23198 29588 23204 29640
rect 23256 29628 23262 29640
rect 23474 29637 23480 29640
rect 23293 29631 23351 29637
rect 23293 29628 23305 29631
rect 23256 29600 23305 29628
rect 23256 29588 23262 29600
rect 23293 29597 23305 29600
rect 23339 29597 23351 29631
rect 23293 29591 23351 29597
rect 23441 29631 23480 29637
rect 23441 29597 23453 29631
rect 23441 29591 23480 29597
rect 23474 29588 23480 29591
rect 23532 29588 23538 29640
rect 23658 29588 23664 29640
rect 23716 29588 23722 29640
rect 23750 29588 23756 29640
rect 23808 29637 23814 29640
rect 23808 29628 23816 29637
rect 23808 29600 23853 29628
rect 23808 29591 23816 29600
rect 23808 29588 23814 29591
rect 23569 29563 23627 29569
rect 20180 29532 21496 29560
rect 18785 29523 18843 29529
rect 18800 29492 18828 29523
rect 19610 29492 19616 29504
rect 18064 29464 19616 29492
rect 19610 29452 19616 29464
rect 19668 29452 19674 29504
rect 19889 29495 19947 29501
rect 19889 29461 19901 29495
rect 19935 29492 19947 29495
rect 20441 29495 20499 29501
rect 20441 29492 20453 29495
rect 19935 29464 20453 29492
rect 19935 29461 19947 29464
rect 19889 29455 19947 29461
rect 20441 29461 20453 29464
rect 20487 29492 20499 29495
rect 21358 29492 21364 29504
rect 20487 29464 21364 29492
rect 20487 29461 20499 29464
rect 20441 29455 20499 29461
rect 21358 29452 21364 29464
rect 21416 29452 21422 29504
rect 21468 29492 21496 29532
rect 23569 29529 23581 29563
rect 23615 29529 23627 29563
rect 24044 29560 24072 29668
rect 24486 29656 24492 29708
rect 24544 29656 24550 29708
rect 24578 29656 24584 29708
rect 24636 29696 24642 29708
rect 25884 29705 25912 29736
rect 31478 29724 31484 29736
rect 31536 29724 31542 29776
rect 31662 29724 31668 29776
rect 31720 29764 31726 29776
rect 31754 29764 31760 29776
rect 31720 29736 31760 29764
rect 31720 29724 31726 29736
rect 31754 29724 31760 29736
rect 31812 29764 31818 29776
rect 33051 29764 33079 29804
rect 33134 29792 33140 29804
rect 33192 29792 33198 29844
rect 33686 29792 33692 29844
rect 33744 29792 33750 29844
rect 33873 29835 33931 29841
rect 33873 29801 33885 29835
rect 33919 29832 33931 29835
rect 34146 29832 34152 29844
rect 33919 29804 34152 29832
rect 33919 29801 33931 29804
rect 33873 29795 33931 29801
rect 34146 29792 34152 29804
rect 34204 29792 34210 29844
rect 34606 29792 34612 29844
rect 34664 29832 34670 29844
rect 34885 29835 34943 29841
rect 34885 29832 34897 29835
rect 34664 29804 34897 29832
rect 34664 29792 34670 29804
rect 34885 29801 34897 29804
rect 34931 29801 34943 29835
rect 35986 29832 35992 29844
rect 34885 29795 34943 29801
rect 35084 29804 35992 29832
rect 31812 29736 31892 29764
rect 31812 29724 31818 29736
rect 25685 29699 25743 29705
rect 25685 29696 25697 29699
rect 24636 29668 25697 29696
rect 24636 29656 24642 29668
rect 25685 29665 25697 29668
rect 25731 29665 25743 29699
rect 25685 29659 25743 29665
rect 25869 29699 25927 29705
rect 25869 29665 25881 29699
rect 25915 29665 25927 29699
rect 25869 29659 25927 29665
rect 26602 29656 26608 29708
rect 26660 29656 26666 29708
rect 27890 29696 27896 29708
rect 27080 29668 27896 29696
rect 24118 29588 24124 29640
rect 24176 29628 24182 29640
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 24176 29600 24409 29628
rect 24176 29588 24182 29600
rect 24397 29597 24409 29600
rect 24443 29597 24455 29631
rect 24397 29591 24455 29597
rect 24673 29631 24731 29637
rect 24673 29597 24685 29631
rect 24719 29597 24731 29631
rect 24673 29591 24731 29597
rect 24688 29560 24716 29591
rect 24762 29588 24768 29640
rect 24820 29588 24826 29640
rect 25590 29588 25596 29640
rect 25648 29588 25654 29640
rect 25774 29588 25780 29640
rect 25832 29628 25838 29640
rect 26329 29631 26387 29637
rect 26329 29628 26341 29631
rect 25832 29600 26341 29628
rect 25832 29588 25838 29600
rect 26329 29597 26341 29600
rect 26375 29597 26387 29631
rect 26329 29591 26387 29597
rect 26421 29631 26479 29637
rect 26421 29597 26433 29631
rect 26467 29628 26479 29631
rect 26510 29628 26516 29640
rect 26467 29600 26516 29628
rect 26467 29597 26479 29600
rect 26421 29591 26479 29597
rect 26510 29588 26516 29600
rect 26568 29588 26574 29640
rect 26697 29631 26755 29637
rect 26697 29597 26709 29631
rect 26743 29628 26755 29631
rect 26786 29628 26792 29640
rect 26743 29600 26792 29628
rect 26743 29597 26755 29600
rect 26697 29591 26755 29597
rect 26786 29588 26792 29600
rect 26844 29588 26850 29640
rect 27080 29637 27108 29668
rect 27890 29656 27896 29668
rect 27948 29656 27954 29708
rect 30466 29656 30472 29708
rect 30524 29656 30530 29708
rect 31864 29705 31892 29736
rect 32600 29736 33079 29764
rect 32600 29705 32628 29736
rect 34238 29724 34244 29776
rect 34296 29724 34302 29776
rect 31849 29699 31907 29705
rect 31849 29665 31861 29699
rect 31895 29665 31907 29699
rect 31849 29659 31907 29665
rect 32585 29699 32643 29705
rect 32585 29665 32597 29699
rect 32631 29665 32643 29699
rect 32585 29659 32643 29665
rect 32766 29656 32772 29708
rect 32824 29656 32830 29708
rect 32876 29668 33364 29696
rect 26973 29631 27031 29637
rect 26973 29597 26985 29631
rect 27019 29597 27031 29631
rect 26973 29591 27031 29597
rect 27065 29631 27123 29637
rect 27065 29597 27077 29631
rect 27111 29597 27123 29631
rect 27065 29591 27123 29597
rect 24044 29532 24716 29560
rect 23569 29523 23627 29529
rect 21818 29492 21824 29504
rect 21468 29464 21824 29492
rect 21818 29452 21824 29464
rect 21876 29452 21882 29504
rect 22094 29452 22100 29504
rect 22152 29492 22158 29504
rect 23584 29492 23612 29523
rect 25314 29520 25320 29572
rect 25372 29560 25378 29572
rect 26988 29560 27016 29591
rect 27338 29588 27344 29640
rect 27396 29588 27402 29640
rect 27430 29588 27436 29640
rect 27488 29588 27494 29640
rect 27614 29588 27620 29640
rect 27672 29588 27678 29640
rect 28534 29588 28540 29640
rect 28592 29628 28598 29640
rect 29549 29631 29607 29637
rect 29549 29628 29561 29631
rect 28592 29600 29561 29628
rect 28592 29588 28598 29600
rect 29549 29597 29561 29600
rect 29595 29597 29607 29631
rect 29549 29591 29607 29597
rect 29730 29588 29736 29640
rect 29788 29588 29794 29640
rect 29822 29588 29828 29640
rect 29880 29588 29886 29640
rect 30098 29588 30104 29640
rect 30156 29628 30162 29640
rect 30193 29631 30251 29637
rect 30193 29628 30205 29631
rect 30156 29600 30205 29628
rect 30156 29588 30162 29600
rect 30193 29597 30205 29600
rect 30239 29597 30251 29631
rect 30193 29591 30251 29597
rect 30285 29631 30343 29637
rect 30285 29597 30297 29631
rect 30331 29628 30343 29631
rect 30374 29628 30380 29640
rect 30331 29600 30380 29628
rect 30331 29597 30343 29600
rect 30285 29591 30343 29597
rect 30374 29588 30380 29600
rect 30432 29628 30438 29640
rect 31018 29628 31024 29640
rect 30432 29600 31024 29628
rect 30432 29588 30438 29600
rect 31018 29588 31024 29600
rect 31076 29588 31082 29640
rect 31110 29588 31116 29640
rect 31168 29588 31174 29640
rect 25372 29532 27016 29560
rect 27157 29563 27215 29569
rect 25372 29520 25378 29532
rect 27157 29529 27169 29563
rect 27203 29560 27215 29563
rect 27246 29560 27252 29572
rect 27203 29532 27252 29560
rect 27203 29529 27215 29532
rect 27157 29523 27215 29529
rect 27246 29520 27252 29532
rect 27304 29560 27310 29572
rect 27304 29532 27844 29560
rect 27304 29520 27310 29532
rect 25498 29492 25504 29504
rect 22152 29464 25504 29492
rect 22152 29452 22158 29464
rect 25498 29452 25504 29464
rect 25556 29452 25562 29504
rect 25866 29452 25872 29504
rect 25924 29452 25930 29504
rect 26510 29452 26516 29504
rect 26568 29492 26574 29504
rect 27525 29495 27583 29501
rect 27525 29492 27537 29495
rect 26568 29464 27537 29492
rect 26568 29452 26574 29464
rect 27525 29461 27537 29464
rect 27571 29461 27583 29495
rect 27816 29492 27844 29532
rect 28994 29520 29000 29572
rect 29052 29560 29058 29572
rect 29181 29563 29239 29569
rect 29181 29560 29193 29563
rect 29052 29532 29193 29560
rect 29052 29520 29058 29532
rect 29181 29529 29193 29532
rect 29227 29529 29239 29563
rect 32876 29560 32904 29668
rect 33336 29637 33364 29668
rect 34422 29656 34428 29708
rect 34480 29696 34486 29708
rect 34793 29699 34851 29705
rect 34793 29696 34805 29699
rect 34480 29668 34805 29696
rect 34480 29656 34486 29668
rect 34793 29665 34805 29668
rect 34839 29665 34851 29699
rect 34793 29659 34851 29665
rect 34974 29656 34980 29708
rect 35032 29656 35038 29708
rect 33132 29631 33190 29637
rect 33132 29597 33144 29631
rect 33178 29597 33190 29631
rect 33132 29591 33190 29597
rect 33229 29631 33287 29637
rect 33229 29597 33241 29631
rect 33275 29597 33287 29631
rect 33229 29591 33287 29597
rect 33321 29631 33379 29637
rect 33321 29597 33333 29631
rect 33367 29597 33379 29631
rect 33321 29591 33379 29597
rect 29181 29523 29239 29529
rect 30392 29532 32904 29560
rect 30392 29492 30420 29532
rect 33042 29520 33048 29572
rect 33100 29560 33106 29572
rect 33152 29560 33180 29591
rect 33100 29532 33180 29560
rect 33100 29520 33106 29532
rect 27816 29464 30420 29492
rect 30469 29495 30527 29501
rect 27525 29455 27583 29461
rect 30469 29461 30481 29495
rect 30515 29492 30527 29495
rect 30558 29492 30564 29504
rect 30515 29464 30564 29492
rect 30515 29461 30527 29464
rect 30469 29455 30527 29461
rect 30558 29452 30564 29464
rect 30616 29452 30622 29504
rect 31294 29452 31300 29504
rect 31352 29492 31358 29504
rect 32125 29495 32183 29501
rect 32125 29492 32137 29495
rect 31352 29464 32137 29492
rect 31352 29452 31358 29464
rect 32125 29461 32137 29464
rect 32171 29461 32183 29495
rect 32125 29455 32183 29461
rect 32398 29452 32404 29504
rect 32456 29492 32462 29504
rect 32493 29495 32551 29501
rect 32493 29492 32505 29495
rect 32456 29464 32505 29492
rect 32456 29452 32462 29464
rect 32493 29461 32505 29464
rect 32539 29461 32551 29495
rect 32493 29455 32551 29461
rect 32858 29452 32864 29504
rect 32916 29492 32922 29504
rect 33247 29492 33275 29591
rect 33410 29588 33416 29640
rect 33468 29637 33474 29640
rect 33468 29631 33507 29637
rect 33495 29597 33507 29631
rect 33468 29591 33507 29597
rect 33468 29588 33474 29591
rect 33594 29588 33600 29640
rect 33652 29588 33658 29640
rect 35084 29637 35112 29804
rect 35986 29792 35992 29804
rect 36044 29792 36050 29844
rect 36078 29792 36084 29844
rect 36136 29832 36142 29844
rect 36136 29804 36952 29832
rect 36136 29792 36142 29804
rect 35526 29764 35532 29776
rect 35360 29736 35532 29764
rect 35360 29637 35388 29736
rect 35526 29724 35532 29736
rect 35584 29724 35590 29776
rect 35621 29767 35679 29773
rect 35621 29733 35633 29767
rect 35667 29733 35679 29767
rect 35621 29727 35679 29733
rect 36357 29767 36415 29773
rect 36357 29733 36369 29767
rect 36403 29764 36415 29767
rect 36403 29736 36676 29764
rect 36403 29733 36415 29736
rect 36357 29727 36415 29733
rect 35636 29696 35664 29727
rect 36648 29696 36676 29736
rect 36814 29696 36820 29708
rect 35636 29668 36492 29696
rect 36648 29668 36820 29696
rect 34701 29631 34759 29637
rect 34701 29597 34713 29631
rect 34747 29597 34759 29631
rect 34701 29591 34759 29597
rect 35069 29631 35127 29637
rect 35069 29597 35081 29631
rect 35115 29597 35127 29631
rect 35253 29631 35311 29637
rect 35253 29606 35265 29631
rect 35069 29591 35127 29597
rect 35176 29597 35265 29606
rect 35299 29597 35311 29631
rect 35176 29591 35311 29597
rect 35345 29631 35403 29637
rect 35345 29597 35357 29631
rect 35391 29597 35403 29631
rect 35345 29591 35403 29597
rect 33870 29520 33876 29572
rect 33928 29520 33934 29572
rect 34054 29520 34060 29572
rect 34112 29560 34118 29572
rect 34717 29560 34745 29591
rect 35176 29578 35296 29591
rect 35434 29588 35440 29640
rect 35492 29588 35498 29640
rect 35618 29588 35624 29640
rect 35676 29628 35682 29640
rect 35713 29631 35771 29637
rect 35713 29628 35725 29631
rect 35676 29600 35725 29628
rect 35676 29588 35682 29600
rect 35713 29597 35725 29600
rect 35759 29597 35771 29631
rect 35713 29591 35771 29597
rect 35806 29631 35864 29637
rect 35806 29597 35818 29631
rect 35852 29628 35864 29631
rect 35894 29628 35900 29640
rect 35852 29600 35900 29628
rect 35852 29597 35864 29600
rect 35806 29591 35864 29597
rect 34790 29560 34796 29572
rect 34112 29532 34796 29560
rect 34112 29520 34118 29532
rect 34790 29520 34796 29532
rect 34848 29520 34854 29572
rect 32916 29464 33275 29492
rect 32916 29452 32922 29464
rect 33410 29452 33416 29504
rect 33468 29492 33474 29504
rect 35176 29492 35204 29578
rect 35821 29560 35849 29591
rect 35894 29588 35900 29600
rect 35952 29588 35958 29640
rect 36219 29631 36277 29637
rect 36219 29597 36231 29631
rect 36265 29628 36277 29631
rect 36354 29628 36360 29640
rect 36265 29600 36360 29628
rect 36265 29597 36277 29600
rect 36219 29591 36277 29597
rect 36354 29588 36360 29600
rect 36412 29588 36418 29640
rect 36464 29628 36492 29668
rect 36814 29656 36820 29668
rect 36872 29656 36878 29708
rect 36633 29631 36691 29637
rect 36633 29628 36645 29631
rect 36464 29600 36645 29628
rect 36633 29597 36645 29600
rect 36679 29597 36691 29631
rect 36633 29591 36691 29597
rect 36722 29588 36728 29640
rect 36780 29628 36786 29640
rect 36924 29637 36952 29804
rect 38654 29792 38660 29844
rect 38712 29832 38718 29844
rect 38933 29835 38991 29841
rect 38933 29832 38945 29835
rect 38712 29804 38945 29832
rect 38712 29792 38718 29804
rect 38933 29801 38945 29804
rect 38979 29801 38991 29835
rect 38933 29795 38991 29801
rect 40313 29835 40371 29841
rect 40313 29801 40325 29835
rect 40359 29832 40371 29835
rect 40678 29832 40684 29844
rect 40359 29804 40684 29832
rect 40359 29801 40371 29804
rect 40313 29795 40371 29801
rect 40678 29792 40684 29804
rect 40736 29792 40742 29844
rect 42150 29792 42156 29844
rect 42208 29792 42214 29844
rect 37277 29767 37335 29773
rect 37277 29733 37289 29767
rect 37323 29764 37335 29767
rect 40126 29764 40132 29776
rect 37323 29736 40132 29764
rect 37323 29733 37335 29736
rect 37277 29727 37335 29733
rect 40126 29724 40132 29736
rect 40184 29724 40190 29776
rect 38010 29696 38016 29708
rect 37016 29668 38016 29696
rect 37016 29637 37044 29668
rect 38010 29656 38016 29668
rect 38068 29696 38074 29708
rect 38470 29696 38476 29708
rect 38068 29668 38476 29696
rect 38068 29656 38074 29668
rect 38470 29656 38476 29668
rect 38528 29656 38534 29708
rect 39482 29656 39488 29708
rect 39540 29656 39546 29708
rect 40310 29656 40316 29708
rect 40368 29696 40374 29708
rect 40681 29699 40739 29705
rect 40681 29696 40693 29699
rect 40368 29668 40693 29696
rect 40368 29656 40374 29668
rect 40681 29665 40693 29668
rect 40727 29665 40739 29699
rect 40681 29659 40739 29665
rect 36909 29631 36967 29637
rect 36780 29600 36825 29628
rect 36780 29588 36786 29600
rect 36909 29597 36921 29631
rect 36955 29597 36967 29631
rect 36909 29591 36967 29597
rect 37001 29631 37059 29637
rect 37001 29597 37013 29631
rect 37047 29597 37059 29631
rect 37001 29591 37059 29597
rect 37090 29588 37096 29640
rect 37148 29637 37154 29640
rect 37148 29631 37197 29637
rect 37148 29597 37151 29631
rect 37185 29628 37197 29631
rect 37826 29628 37832 29640
rect 37185 29600 37832 29628
rect 37185 29597 37197 29600
rect 37148 29591 37197 29597
rect 37148 29588 37154 29591
rect 37826 29588 37832 29600
rect 37884 29588 37890 29640
rect 39850 29588 39856 29640
rect 39908 29588 39914 29640
rect 40034 29588 40040 29640
rect 40092 29628 40098 29640
rect 40129 29631 40187 29637
rect 40129 29628 40141 29631
rect 40092 29600 40141 29628
rect 40092 29588 40098 29600
rect 40129 29597 40141 29600
rect 40175 29597 40187 29631
rect 40129 29591 40187 29597
rect 40402 29588 40408 29640
rect 40460 29588 40466 29640
rect 35544 29532 35849 29560
rect 35989 29563 36047 29569
rect 35544 29504 35572 29532
rect 35989 29529 36001 29563
rect 36035 29529 36047 29563
rect 35989 29523 36047 29529
rect 36081 29563 36139 29569
rect 36081 29529 36093 29563
rect 36127 29560 36139 29563
rect 37366 29560 37372 29572
rect 36127 29532 36860 29560
rect 36127 29529 36139 29532
rect 36081 29523 36139 29529
rect 33468 29464 35204 29492
rect 33468 29452 33474 29464
rect 35526 29452 35532 29504
rect 35584 29452 35590 29504
rect 35710 29452 35716 29504
rect 35768 29492 35774 29504
rect 36004 29492 36032 29523
rect 36170 29492 36176 29504
rect 35768 29464 36176 29492
rect 35768 29452 35774 29464
rect 36170 29452 36176 29464
rect 36228 29452 36234 29504
rect 36832 29492 36860 29532
rect 37108 29532 37372 29560
rect 37108 29492 37136 29532
rect 37366 29520 37372 29532
rect 37424 29520 37430 29572
rect 39945 29563 40003 29569
rect 39945 29529 39957 29563
rect 39991 29560 40003 29563
rect 40770 29560 40776 29572
rect 39991 29532 40776 29560
rect 39991 29529 40003 29532
rect 39945 29523 40003 29529
rect 40770 29520 40776 29532
rect 40828 29520 40834 29572
rect 41690 29520 41696 29572
rect 41748 29520 41754 29572
rect 36832 29464 37136 29492
rect 38562 29452 38568 29504
rect 38620 29492 38626 29504
rect 40494 29492 40500 29504
rect 38620 29464 40500 29492
rect 38620 29452 38626 29464
rect 40494 29452 40500 29464
rect 40552 29452 40558 29504
rect 1104 29402 42504 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 42504 29402
rect 1104 29328 42504 29350
rect 3786 29288 3792 29300
rect 2240 29260 3792 29288
rect 1762 29112 1768 29164
rect 1820 29112 1826 29164
rect 1946 29112 1952 29164
rect 2004 29112 2010 29164
rect 2240 29161 2268 29260
rect 3786 29248 3792 29260
rect 3844 29248 3850 29300
rect 4706 29248 4712 29300
rect 4764 29288 4770 29300
rect 4801 29291 4859 29297
rect 4801 29288 4813 29291
rect 4764 29260 4813 29288
rect 4764 29248 4770 29260
rect 4801 29257 4813 29260
rect 4847 29257 4859 29291
rect 4801 29251 4859 29257
rect 5534 29248 5540 29300
rect 5592 29248 5598 29300
rect 5718 29248 5724 29300
rect 5776 29288 5782 29300
rect 6365 29291 6423 29297
rect 5776 29260 6132 29288
rect 5776 29248 5782 29260
rect 2406 29180 2412 29232
rect 2464 29180 2470 29232
rect 2547 29223 2605 29229
rect 2547 29189 2559 29223
rect 2593 29220 2605 29223
rect 3050 29220 3056 29232
rect 2593 29192 3056 29220
rect 2593 29189 2605 29192
rect 2547 29183 2605 29189
rect 3050 29180 3056 29192
rect 3108 29180 3114 29232
rect 3142 29180 3148 29232
rect 3200 29220 3206 29232
rect 3513 29223 3571 29229
rect 3513 29220 3525 29223
rect 3200 29192 3525 29220
rect 3200 29180 3206 29192
rect 3513 29189 3525 29192
rect 3559 29189 3571 29223
rect 3513 29183 3571 29189
rect 4430 29180 4436 29232
rect 4488 29180 4494 29232
rect 5905 29223 5963 29229
rect 5905 29220 5917 29223
rect 4540 29192 5917 29220
rect 2225 29155 2283 29161
rect 2225 29121 2237 29155
rect 2271 29121 2283 29155
rect 2225 29115 2283 29121
rect 2317 29155 2375 29161
rect 2317 29121 2329 29155
rect 2363 29121 2375 29155
rect 2317 29115 2375 29121
rect 3421 29155 3479 29161
rect 3421 29121 3433 29155
rect 3467 29152 3479 29155
rect 3602 29152 3608 29164
rect 3467 29124 3608 29152
rect 3467 29121 3479 29124
rect 3421 29115 3479 29121
rect 1857 29087 1915 29093
rect 1857 29053 1869 29087
rect 1903 29084 1915 29087
rect 2332 29084 2360 29115
rect 3602 29112 3608 29124
rect 3660 29112 3666 29164
rect 4154 29112 4160 29164
rect 4212 29112 4218 29164
rect 4249 29155 4307 29161
rect 4249 29121 4261 29155
rect 4295 29121 4307 29155
rect 4249 29115 4307 29121
rect 1903 29056 2360 29084
rect 1903 29053 1915 29056
rect 1857 29047 1915 29053
rect 2332 29016 2360 29056
rect 2685 29087 2743 29093
rect 2685 29053 2697 29087
rect 2731 29084 2743 29087
rect 2777 29087 2835 29093
rect 2777 29084 2789 29087
rect 2731 29056 2789 29084
rect 2731 29053 2743 29056
rect 2685 29047 2743 29053
rect 2777 29053 2789 29056
rect 2823 29053 2835 29087
rect 4264 29084 4292 29115
rect 4540 29084 4568 29192
rect 5905 29189 5917 29192
rect 5951 29189 5963 29223
rect 5905 29183 5963 29189
rect 4617 29155 4675 29161
rect 4617 29121 4629 29155
rect 4663 29152 4675 29155
rect 4985 29155 5043 29161
rect 4985 29152 4997 29155
rect 4663 29124 4997 29152
rect 4663 29121 4675 29124
rect 4617 29115 4675 29121
rect 4985 29121 4997 29124
rect 5031 29121 5043 29155
rect 4985 29115 5043 29121
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29121 5135 29155
rect 5077 29115 5135 29121
rect 4706 29084 4712 29096
rect 4264 29056 4712 29084
rect 2777 29047 2835 29053
rect 4706 29044 4712 29056
rect 4764 29044 4770 29096
rect 3418 29016 3424 29028
rect 2332 28988 3424 29016
rect 3418 28976 3424 28988
rect 3476 28976 3482 29028
rect 3970 28976 3976 29028
rect 4028 29016 4034 29028
rect 5092 29016 5120 29115
rect 5166 29112 5172 29164
rect 5224 29112 5230 29164
rect 5287 29155 5345 29161
rect 5287 29121 5299 29155
rect 5333 29152 5345 29155
rect 5333 29124 5672 29152
rect 5333 29121 5350 29124
rect 5287 29115 5350 29121
rect 4028 28988 5120 29016
rect 4028 28976 4034 28988
rect 5166 28976 5172 29028
rect 5224 29016 5230 29028
rect 5322 29016 5350 29115
rect 5445 29087 5503 29093
rect 5445 29053 5457 29087
rect 5491 29053 5503 29087
rect 5644 29084 5672 29124
rect 5718 29112 5724 29164
rect 5776 29112 5782 29164
rect 5810 29112 5816 29164
rect 5868 29112 5874 29164
rect 6104 29161 6132 29260
rect 6365 29257 6377 29291
rect 6411 29288 6423 29291
rect 6454 29288 6460 29300
rect 6411 29260 6460 29288
rect 6411 29257 6423 29260
rect 6365 29251 6423 29257
rect 6454 29248 6460 29260
rect 6512 29248 6518 29300
rect 11790 29248 11796 29300
rect 11848 29288 11854 29300
rect 12069 29291 12127 29297
rect 12069 29288 12081 29291
rect 11848 29260 12081 29288
rect 11848 29248 11854 29260
rect 12069 29257 12081 29260
rect 12115 29257 12127 29291
rect 12069 29251 12127 29257
rect 13354 29248 13360 29300
rect 13412 29288 13418 29300
rect 13633 29291 13691 29297
rect 13633 29288 13645 29291
rect 13412 29260 13645 29288
rect 13412 29248 13418 29260
rect 13633 29257 13645 29260
rect 13679 29257 13691 29291
rect 13633 29251 13691 29257
rect 16482 29248 16488 29300
rect 16540 29288 16546 29300
rect 17037 29291 17095 29297
rect 17037 29288 17049 29291
rect 16540 29260 17049 29288
rect 16540 29248 16546 29260
rect 17037 29257 17049 29260
rect 17083 29257 17095 29291
rect 17037 29251 17095 29257
rect 17402 29248 17408 29300
rect 17460 29248 17466 29300
rect 17586 29248 17592 29300
rect 17644 29288 17650 29300
rect 18230 29288 18236 29300
rect 17644 29260 18236 29288
rect 17644 29248 17650 29260
rect 18230 29248 18236 29260
rect 18288 29248 18294 29300
rect 18325 29291 18383 29297
rect 18325 29257 18337 29291
rect 18371 29288 18383 29291
rect 18966 29288 18972 29300
rect 18371 29260 18972 29288
rect 18371 29257 18383 29260
rect 18325 29251 18383 29257
rect 18966 29248 18972 29260
rect 19024 29248 19030 29300
rect 19243 29248 19249 29300
rect 19301 29288 19307 29300
rect 19981 29291 20039 29297
rect 19981 29288 19993 29291
rect 19301 29260 19993 29288
rect 19301 29248 19307 29260
rect 19981 29257 19993 29260
rect 20027 29257 20039 29291
rect 19981 29251 20039 29257
rect 21358 29248 21364 29300
rect 21416 29288 21422 29300
rect 24029 29291 24087 29297
rect 21416 29260 23612 29288
rect 21416 29248 21422 29260
rect 23584 29232 23612 29260
rect 24029 29257 24041 29291
rect 24075 29288 24087 29291
rect 24762 29288 24768 29300
rect 24075 29260 24768 29288
rect 24075 29257 24087 29260
rect 24029 29251 24087 29257
rect 24762 29248 24768 29260
rect 24820 29248 24826 29300
rect 25222 29248 25228 29300
rect 25280 29288 25286 29300
rect 25961 29291 26019 29297
rect 25961 29288 25973 29291
rect 25280 29260 25973 29288
rect 25280 29248 25286 29260
rect 25961 29257 25973 29260
rect 26007 29257 26019 29291
rect 25961 29251 26019 29257
rect 26139 29291 26197 29297
rect 26139 29257 26151 29291
rect 26185 29288 26197 29291
rect 26185 29260 26740 29288
rect 26185 29257 26197 29260
rect 26139 29251 26197 29257
rect 17126 29220 17132 29232
rect 12268 29192 17132 29220
rect 6089 29155 6147 29161
rect 6089 29121 6101 29155
rect 6135 29121 6147 29155
rect 6089 29115 6147 29121
rect 6270 29112 6276 29164
rect 6328 29152 6334 29164
rect 6733 29155 6791 29161
rect 6733 29152 6745 29155
rect 6328 29124 6745 29152
rect 6328 29112 6334 29124
rect 6733 29121 6745 29124
rect 6779 29152 6791 29155
rect 7377 29155 7435 29161
rect 7377 29152 7389 29155
rect 6779 29124 7389 29152
rect 6779 29121 6791 29124
rect 6733 29115 6791 29121
rect 7377 29121 7389 29124
rect 7423 29121 7435 29155
rect 7377 29115 7435 29121
rect 7469 29155 7527 29161
rect 7469 29121 7481 29155
rect 7515 29152 7527 29155
rect 8202 29152 8208 29164
rect 7515 29124 8208 29152
rect 7515 29121 7527 29124
rect 7469 29115 7527 29121
rect 8202 29112 8208 29124
rect 8260 29112 8266 29164
rect 12268 29152 12296 29192
rect 17126 29180 17132 29192
rect 17184 29180 17190 29232
rect 17221 29223 17279 29229
rect 17221 29189 17233 29223
rect 17267 29220 17279 29223
rect 17267 29192 17632 29220
rect 17267 29189 17279 29192
rect 17221 29183 17279 29189
rect 10902 29124 11008 29152
rect 5828 29084 5856 29112
rect 10980 29096 11008 29124
rect 11256 29124 12296 29152
rect 12345 29155 12403 29161
rect 5644 29056 5856 29084
rect 5445 29047 5503 29053
rect 5224 28988 5350 29016
rect 5460 29016 5488 29047
rect 6546 29044 6552 29096
rect 6604 29084 6610 29096
rect 6641 29087 6699 29093
rect 6641 29084 6653 29087
rect 6604 29056 6653 29084
rect 6604 29044 6610 29056
rect 6641 29053 6653 29056
rect 6687 29053 6699 29087
rect 6641 29047 6699 29053
rect 9490 29044 9496 29096
rect 9548 29044 9554 29096
rect 9766 29044 9772 29096
rect 9824 29044 9830 29096
rect 10962 29044 10968 29096
rect 11020 29044 11026 29096
rect 5718 29016 5724 29028
rect 5460 28988 5724 29016
rect 5224 28976 5230 28988
rect 5718 28976 5724 28988
rect 5776 29016 5782 29028
rect 6564 29016 6592 29044
rect 11256 29028 11284 29124
rect 12345 29121 12357 29155
rect 12391 29152 12403 29155
rect 12805 29155 12863 29161
rect 12805 29152 12817 29155
rect 12391 29124 12817 29152
rect 12391 29121 12403 29124
rect 12345 29115 12403 29121
rect 12805 29121 12817 29124
rect 12851 29121 12863 29155
rect 12805 29115 12863 29121
rect 13446 29112 13452 29164
rect 13504 29112 13510 29164
rect 13538 29112 13544 29164
rect 13596 29112 13602 29164
rect 13725 29155 13783 29161
rect 13725 29121 13737 29155
rect 13771 29121 13783 29155
rect 13725 29115 13783 29121
rect 16945 29155 17003 29161
rect 16945 29121 16957 29155
rect 16991 29152 17003 29155
rect 17034 29152 17040 29164
rect 16991 29124 17040 29152
rect 16991 29121 17003 29124
rect 16945 29115 17003 29121
rect 12253 29087 12311 29093
rect 12253 29053 12265 29087
rect 12299 29084 12311 29087
rect 12299 29056 12434 29084
rect 12299 29053 12311 29056
rect 12253 29047 12311 29053
rect 5776 28988 6592 29016
rect 5776 28976 5782 28988
rect 11238 28976 11244 29028
rect 11296 28976 11302 29028
rect 12406 29016 12434 29056
rect 12526 29044 12532 29096
rect 12584 29084 12590 29096
rect 12713 29087 12771 29093
rect 12713 29084 12725 29087
rect 12584 29056 12725 29084
rect 12584 29044 12590 29056
rect 12713 29053 12725 29056
rect 12759 29084 12771 29087
rect 13262 29084 13268 29096
rect 12759 29056 13268 29084
rect 12759 29053 12771 29056
rect 12713 29047 12771 29053
rect 13262 29044 13268 29056
rect 13320 29084 13326 29096
rect 13740 29084 13768 29115
rect 17034 29112 17040 29124
rect 17092 29112 17098 29164
rect 17144 29152 17172 29180
rect 17604 29161 17632 29192
rect 17770 29180 17776 29232
rect 17828 29220 17834 29232
rect 18509 29223 18567 29229
rect 17828 29192 18460 29220
rect 17828 29180 17834 29192
rect 17313 29155 17371 29161
rect 17313 29152 17325 29155
rect 17144 29124 17325 29152
rect 17313 29121 17325 29124
rect 17359 29121 17371 29155
rect 17313 29115 17371 29121
rect 17589 29155 17647 29161
rect 17589 29121 17601 29155
rect 17635 29152 17647 29155
rect 17635 29124 17825 29152
rect 17635 29121 17647 29124
rect 17589 29115 17647 29121
rect 13320 29056 13768 29084
rect 13320 29044 13326 29056
rect 16850 29044 16856 29096
rect 16908 29084 16914 29096
rect 17126 29084 17132 29096
rect 16908 29056 17132 29084
rect 16908 29044 16914 29056
rect 17126 29044 17132 29056
rect 17184 29044 17190 29096
rect 13538 29016 13544 29028
rect 12406 28988 13544 29016
rect 13538 28976 13544 28988
rect 13596 28976 13602 29028
rect 17221 29019 17279 29025
rect 17221 28985 17233 29019
rect 17267 29016 17279 29019
rect 17310 29016 17316 29028
rect 17267 28988 17316 29016
rect 17267 28985 17279 28988
rect 17221 28979 17279 28985
rect 17310 28976 17316 28988
rect 17368 28976 17374 29028
rect 17589 29019 17647 29025
rect 17589 28985 17601 29019
rect 17635 29016 17647 29019
rect 17678 29016 17684 29028
rect 17635 28988 17684 29016
rect 17635 28985 17647 28988
rect 17589 28979 17647 28985
rect 17678 28976 17684 28988
rect 17736 28976 17742 29028
rect 17797 29016 17825 29124
rect 17954 29112 17960 29164
rect 18012 29152 18018 29164
rect 18432 29161 18460 29192
rect 18509 29189 18521 29223
rect 18555 29220 18567 29223
rect 18690 29220 18696 29232
rect 18555 29192 18696 29220
rect 18555 29189 18567 29192
rect 18509 29183 18567 29189
rect 18690 29180 18696 29192
rect 18748 29220 18754 29232
rect 19889 29223 19947 29229
rect 19889 29220 19901 29223
rect 18748 29192 19901 29220
rect 18748 29180 18754 29192
rect 19889 29189 19901 29192
rect 19935 29220 19947 29223
rect 20809 29223 20867 29229
rect 19935 29192 20760 29220
rect 19935 29189 19947 29192
rect 19889 29183 19947 29189
rect 18141 29155 18199 29161
rect 18141 29152 18153 29155
rect 18012 29124 18153 29152
rect 18012 29112 18018 29124
rect 18141 29121 18153 29124
rect 18187 29121 18199 29155
rect 18141 29115 18199 29121
rect 18417 29155 18475 29161
rect 18417 29121 18429 29155
rect 18463 29121 18475 29155
rect 18417 29115 18475 29121
rect 18601 29155 18659 29161
rect 18601 29121 18613 29155
rect 18647 29152 18659 29155
rect 18836 29152 19334 29162
rect 19426 29152 19432 29164
rect 18647 29134 19432 29152
rect 18647 29124 18864 29134
rect 19306 29124 19432 29134
rect 18647 29121 18659 29124
rect 18601 29115 18659 29121
rect 17862 29044 17868 29096
rect 17920 29044 17926 29096
rect 18432 29084 18460 29115
rect 19426 29112 19432 29124
rect 19484 29112 19490 29164
rect 19610 29112 19616 29164
rect 19668 29112 19674 29164
rect 19794 29112 19800 29164
rect 19852 29112 19858 29164
rect 20732 29161 20760 29192
rect 20809 29189 20821 29223
rect 20855 29220 20867 29223
rect 20855 29192 22232 29220
rect 20855 29189 20867 29192
rect 20809 29183 20867 29189
rect 20717 29155 20775 29161
rect 20717 29121 20729 29155
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 20990 29112 20996 29164
rect 21048 29152 21054 29164
rect 21192 29161 21220 29192
rect 21085 29155 21143 29161
rect 21085 29152 21097 29155
rect 21048 29124 21097 29152
rect 21048 29112 21054 29124
rect 21085 29121 21097 29124
rect 21131 29121 21143 29155
rect 21085 29115 21143 29121
rect 21177 29155 21235 29161
rect 21177 29121 21189 29155
rect 21223 29121 21235 29155
rect 21177 29115 21235 29121
rect 21361 29155 21419 29161
rect 21361 29121 21373 29155
rect 21407 29121 21419 29155
rect 21361 29115 21419 29121
rect 21453 29155 21511 29161
rect 21453 29121 21465 29155
rect 21499 29152 21511 29155
rect 21818 29152 21824 29164
rect 21499 29124 21824 29152
rect 21499 29121 21511 29124
rect 21453 29115 21511 29121
rect 18432 29056 18828 29084
rect 18690 29016 18696 29028
rect 17797 28988 18696 29016
rect 18690 28976 18696 28988
rect 18748 28976 18754 29028
rect 18800 29016 18828 29056
rect 19058 29044 19064 29096
rect 19116 29084 19122 29096
rect 19199 29087 19257 29093
rect 19199 29084 19211 29087
rect 19116 29056 19211 29084
rect 19116 29044 19122 29056
rect 19199 29053 19211 29056
rect 19245 29053 19257 29087
rect 19199 29047 19257 29053
rect 19518 29044 19524 29096
rect 19576 29044 19582 29096
rect 20165 29087 20223 29093
rect 20165 29053 20177 29087
rect 20211 29084 20223 29087
rect 20254 29084 20260 29096
rect 20211 29056 20260 29084
rect 20211 29053 20223 29056
rect 20165 29047 20223 29053
rect 20254 29044 20260 29056
rect 20312 29084 20318 29096
rect 21008 29084 21036 29112
rect 20312 29056 21036 29084
rect 21376 29084 21404 29115
rect 21818 29112 21824 29124
rect 21876 29112 21882 29164
rect 22002 29161 22008 29164
rect 21984 29155 22008 29161
rect 21984 29152 21996 29155
rect 21928 29124 21996 29152
rect 21928 29084 21956 29124
rect 21984 29121 21996 29124
rect 21984 29115 22008 29121
rect 22002 29112 22008 29115
rect 22060 29112 22066 29164
rect 22094 29112 22100 29164
rect 22152 29112 22158 29164
rect 22204 29161 22232 29192
rect 22462 29180 22468 29232
rect 22520 29220 22526 29232
rect 22738 29220 22744 29232
rect 22520 29192 22744 29220
rect 22520 29180 22526 29192
rect 22738 29180 22744 29192
rect 22796 29180 22802 29232
rect 23382 29220 23388 29232
rect 22940 29192 23388 29220
rect 22940 29161 22968 29192
rect 23382 29180 23388 29192
rect 23440 29180 23446 29232
rect 23566 29180 23572 29232
rect 23624 29220 23630 29232
rect 23845 29223 23903 29229
rect 23845 29220 23857 29223
rect 23624 29192 23857 29220
rect 23624 29180 23630 29192
rect 23845 29189 23857 29192
rect 23891 29220 23903 29223
rect 24394 29220 24400 29232
rect 23891 29192 24400 29220
rect 23891 29189 23903 29192
rect 23845 29183 23903 29189
rect 24394 29180 24400 29192
rect 24452 29180 24458 29232
rect 25866 29180 25872 29232
rect 25924 29220 25930 29232
rect 25924 29192 26556 29220
rect 25924 29180 25930 29192
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29121 22247 29155
rect 22833 29155 22891 29161
rect 22833 29152 22845 29155
rect 22189 29115 22247 29121
rect 22480 29124 22845 29152
rect 21376 29056 21956 29084
rect 20312 29044 20318 29056
rect 19610 29016 19616 29028
rect 18800 28988 19616 29016
rect 19610 28976 19616 28988
rect 19668 28976 19674 29028
rect 2038 28908 2044 28960
rect 2096 28908 2102 28960
rect 4338 28908 4344 28960
rect 4396 28948 4402 28960
rect 5074 28948 5080 28960
rect 4396 28920 5080 28948
rect 4396 28908 4402 28920
rect 5074 28908 5080 28920
rect 5132 28908 5138 28960
rect 5626 28908 5632 28960
rect 5684 28948 5690 28960
rect 12894 28948 12900 28960
rect 5684 28920 12900 28948
rect 5684 28908 5690 28920
rect 12894 28908 12900 28920
rect 12952 28908 12958 28960
rect 12986 28908 12992 28960
rect 13044 28948 13050 28960
rect 17770 28948 17776 28960
rect 13044 28920 17776 28948
rect 13044 28908 13050 28920
rect 17770 28908 17776 28920
rect 17828 28908 17834 28960
rect 17957 28951 18015 28957
rect 17957 28917 17969 28951
rect 18003 28948 18015 28951
rect 18322 28948 18328 28960
rect 18003 28920 18328 28948
rect 18003 28917 18015 28920
rect 17957 28911 18015 28917
rect 18322 28908 18328 28920
rect 18380 28908 18386 28960
rect 21450 28908 21456 28960
rect 21508 28948 21514 28960
rect 21637 28951 21695 28957
rect 21637 28948 21649 28951
rect 21508 28920 21649 28948
rect 21508 28908 21514 28920
rect 21637 28917 21649 28920
rect 21683 28917 21695 28951
rect 21637 28911 21695 28917
rect 22370 28908 22376 28960
rect 22428 28948 22434 28960
rect 22480 28957 22508 29124
rect 22833 29121 22845 29124
rect 22879 29121 22891 29155
rect 22833 29115 22891 29121
rect 22925 29155 22983 29161
rect 22925 29121 22937 29155
rect 22971 29121 22983 29155
rect 22925 29115 22983 29121
rect 22554 29044 22560 29096
rect 22612 29084 22618 29096
rect 22940 29084 22968 29115
rect 23106 29112 23112 29164
rect 23164 29112 23170 29164
rect 23201 29155 23259 29161
rect 23201 29121 23213 29155
rect 23247 29121 23259 29155
rect 23201 29115 23259 29121
rect 22612 29056 22968 29084
rect 22612 29044 22618 29056
rect 23014 29044 23020 29096
rect 23072 29084 23078 29096
rect 23216 29084 23244 29115
rect 23290 29112 23296 29164
rect 23348 29152 23354 29164
rect 24118 29152 24124 29164
rect 23348 29124 24124 29152
rect 23348 29112 23354 29124
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 24302 29112 24308 29164
rect 24360 29112 24366 29164
rect 25222 29112 25228 29164
rect 25280 29112 25286 29164
rect 25501 29155 25559 29161
rect 25501 29121 25513 29155
rect 25547 29152 25559 29155
rect 25774 29152 25780 29164
rect 25547 29124 25780 29152
rect 25547 29121 25559 29124
rect 25501 29115 25559 29121
rect 25774 29112 25780 29124
rect 25832 29112 25838 29164
rect 26528 29161 26556 29192
rect 26602 29180 26608 29232
rect 26660 29180 26666 29232
rect 26712 29220 26740 29260
rect 26786 29248 26792 29300
rect 26844 29288 26850 29300
rect 27065 29291 27123 29297
rect 27065 29288 27077 29291
rect 26844 29260 27077 29288
rect 26844 29248 26850 29260
rect 27065 29257 27077 29260
rect 27111 29288 27123 29291
rect 27430 29288 27436 29300
rect 27111 29260 27436 29288
rect 27111 29257 27123 29260
rect 27065 29251 27123 29257
rect 27430 29248 27436 29260
rect 27488 29248 27494 29300
rect 29178 29288 29184 29300
rect 28276 29260 29184 29288
rect 27154 29220 27160 29232
rect 26712 29192 27160 29220
rect 27154 29180 27160 29192
rect 27212 29220 27218 29232
rect 27249 29223 27307 29229
rect 27249 29220 27261 29223
rect 27212 29192 27261 29220
rect 27212 29180 27218 29192
rect 27249 29189 27261 29192
rect 27295 29189 27307 29223
rect 27249 29183 27307 29189
rect 27798 29180 27804 29232
rect 27856 29180 27862 29232
rect 27890 29180 27896 29232
rect 27948 29180 27954 29232
rect 26053 29155 26111 29161
rect 26053 29121 26065 29155
rect 26099 29121 26111 29155
rect 26053 29115 26111 29121
rect 26513 29155 26571 29161
rect 26513 29121 26525 29155
rect 26559 29121 26571 29155
rect 26620 29152 26648 29180
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26620 29124 26985 29152
rect 26513 29115 26571 29121
rect 26973 29121 26985 29124
rect 27019 29121 27031 29155
rect 26973 29115 27031 29121
rect 23072 29056 23244 29084
rect 24489 29087 24547 29093
rect 23072 29044 23078 29056
rect 24489 29053 24501 29087
rect 24535 29084 24547 29087
rect 25317 29087 25375 29093
rect 25317 29084 25329 29087
rect 24535 29056 25329 29084
rect 24535 29053 24547 29056
rect 24489 29047 24547 29053
rect 25317 29053 25329 29056
rect 25363 29084 25375 29087
rect 25590 29084 25596 29096
rect 25363 29056 25596 29084
rect 25363 29053 25375 29056
rect 25317 29047 25375 29053
rect 25590 29044 25596 29056
rect 25648 29084 25654 29096
rect 25685 29087 25743 29093
rect 25685 29084 25697 29087
rect 25648 29056 25697 29084
rect 25648 29044 25654 29056
rect 25685 29053 25697 29056
rect 25731 29053 25743 29087
rect 26068 29084 26096 29115
rect 27338 29112 27344 29164
rect 27396 29152 27402 29164
rect 27617 29155 27675 29161
rect 27617 29152 27629 29155
rect 27396 29124 27629 29152
rect 27396 29112 27402 29124
rect 27617 29121 27629 29124
rect 27663 29121 27675 29155
rect 27617 29115 27675 29121
rect 27985 29155 28043 29161
rect 27985 29121 27997 29155
rect 28031 29152 28043 29155
rect 28074 29152 28080 29164
rect 28031 29124 28080 29152
rect 28031 29121 28043 29124
rect 27985 29115 28043 29121
rect 28074 29112 28080 29124
rect 28132 29112 28138 29164
rect 28276 29161 28304 29260
rect 29178 29248 29184 29260
rect 29236 29248 29242 29300
rect 31018 29248 31024 29300
rect 31076 29288 31082 29300
rect 31205 29291 31263 29297
rect 31205 29288 31217 29291
rect 31076 29260 31217 29288
rect 31076 29248 31082 29260
rect 31205 29257 31217 29260
rect 31251 29257 31263 29291
rect 31205 29251 31263 29257
rect 31389 29291 31447 29297
rect 31389 29257 31401 29291
rect 31435 29288 31447 29291
rect 32030 29288 32036 29300
rect 31435 29260 32036 29288
rect 31435 29257 31447 29260
rect 31389 29251 31447 29257
rect 32030 29248 32036 29260
rect 32088 29248 32094 29300
rect 32858 29288 32864 29300
rect 32508 29260 32864 29288
rect 28534 29180 28540 29232
rect 28592 29180 28598 29232
rect 28626 29180 28632 29232
rect 28684 29220 28690 29232
rect 30374 29220 30380 29232
rect 28684 29192 29026 29220
rect 30024 29192 30380 29220
rect 28684 29180 28690 29192
rect 28261 29155 28319 29161
rect 28261 29121 28273 29155
rect 28307 29121 28319 29155
rect 30024 29152 30052 29192
rect 28261 29115 28319 29121
rect 29748 29124 30052 29152
rect 26602 29084 26608 29096
rect 26068 29056 26608 29084
rect 25685 29047 25743 29053
rect 26602 29044 26608 29056
rect 26660 29084 26666 29096
rect 26786 29084 26792 29096
rect 26660 29056 26792 29084
rect 26660 29044 26666 29056
rect 26786 29044 26792 29056
rect 26844 29044 26850 29096
rect 29748 29084 29776 29124
rect 30098 29112 30104 29164
rect 30156 29112 30162 29164
rect 30300 29161 30328 29192
rect 30374 29180 30380 29192
rect 30432 29180 30438 29232
rect 30469 29223 30527 29229
rect 30469 29189 30481 29223
rect 30515 29220 30527 29223
rect 30650 29220 30656 29232
rect 30515 29192 30656 29220
rect 30515 29189 30527 29192
rect 30469 29183 30527 29189
rect 30650 29180 30656 29192
rect 30708 29220 30714 29232
rect 32508 29229 32536 29260
rect 32858 29248 32864 29260
rect 32916 29248 32922 29300
rect 33042 29248 33048 29300
rect 33100 29288 33106 29300
rect 33226 29288 33232 29300
rect 33100 29260 33232 29288
rect 33100 29248 33106 29260
rect 33226 29248 33232 29260
rect 33284 29288 33290 29300
rect 36354 29288 36360 29300
rect 33284 29260 36360 29288
rect 33284 29248 33290 29260
rect 36354 29248 36360 29260
rect 36412 29248 36418 29300
rect 36906 29248 36912 29300
rect 36964 29288 36970 29300
rect 41325 29291 41383 29297
rect 41325 29288 41337 29291
rect 36964 29260 41337 29288
rect 36964 29248 36970 29260
rect 41325 29257 41337 29260
rect 41371 29257 41383 29291
rect 41325 29251 41383 29257
rect 32493 29223 32551 29229
rect 30708 29192 30788 29220
rect 30708 29180 30714 29192
rect 30285 29155 30343 29161
rect 30285 29121 30297 29155
rect 30331 29121 30343 29155
rect 30285 29115 30343 29121
rect 30558 29112 30564 29164
rect 30616 29112 30622 29164
rect 30760 29161 30788 29192
rect 32493 29189 32505 29223
rect 32539 29189 32551 29223
rect 33060 29220 33088 29248
rect 34054 29220 34060 29232
rect 32493 29183 32551 29189
rect 32646 29192 33088 29220
rect 33796 29192 34060 29220
rect 30745 29155 30803 29161
rect 30745 29121 30757 29155
rect 30791 29121 30803 29155
rect 30745 29115 30803 29121
rect 31018 29112 31024 29164
rect 31076 29112 31082 29164
rect 31110 29112 31116 29164
rect 31168 29112 31174 29164
rect 31294 29112 31300 29164
rect 31352 29152 31358 29164
rect 31665 29155 31723 29161
rect 31665 29152 31677 29155
rect 31352 29124 31677 29152
rect 31352 29112 31358 29124
rect 31665 29121 31677 29124
rect 31711 29121 31723 29155
rect 31665 29115 31723 29121
rect 31849 29155 31907 29161
rect 31849 29121 31861 29155
rect 31895 29152 31907 29155
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 31895 29124 32137 29152
rect 31895 29121 31907 29124
rect 31849 29115 31907 29121
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 32214 29112 32220 29164
rect 32272 29152 32278 29164
rect 32646 29161 32674 29192
rect 32401 29155 32459 29161
rect 32272 29124 32317 29152
rect 32272 29112 32278 29124
rect 32401 29121 32413 29155
rect 32447 29121 32459 29155
rect 32401 29115 32459 29121
rect 32631 29155 32689 29161
rect 32631 29121 32643 29155
rect 32677 29121 32689 29155
rect 32631 29115 32689 29121
rect 32861 29155 32919 29161
rect 32861 29121 32873 29155
rect 32907 29152 32919 29155
rect 33042 29152 33048 29164
rect 32907 29124 33048 29152
rect 32907 29121 32919 29124
rect 32861 29115 32919 29121
rect 28092 29056 29776 29084
rect 30009 29087 30067 29093
rect 23477 29019 23535 29025
rect 23477 28985 23489 29019
rect 23523 29016 23535 29019
rect 23658 29016 23664 29028
rect 23523 28988 23664 29016
rect 23523 28985 23535 28988
rect 23477 28979 23535 28985
rect 23658 28976 23664 28988
rect 23716 29016 23722 29028
rect 24578 29016 24584 29028
rect 23716 28988 24584 29016
rect 23716 28976 23722 28988
rect 24578 28976 24584 28988
rect 24636 29016 24642 29028
rect 25409 29019 25467 29025
rect 25409 29016 25421 29019
rect 24636 28988 25421 29016
rect 24636 28976 24642 28988
rect 25409 28985 25421 28988
rect 25455 29016 25467 29019
rect 25777 29019 25835 29025
rect 25777 29016 25789 29019
rect 25455 28988 25789 29016
rect 25455 28985 25467 28988
rect 25409 28979 25467 28985
rect 25777 28985 25789 28988
rect 25823 28985 25835 29019
rect 28092 29016 28120 29056
rect 30009 29053 30021 29087
rect 30055 29084 30067 29087
rect 30116 29084 30144 29112
rect 30837 29087 30895 29093
rect 30837 29084 30849 29087
rect 30055 29056 30849 29084
rect 30055 29053 30067 29056
rect 30009 29047 30067 29053
rect 30837 29053 30849 29056
rect 30883 29053 30895 29087
rect 30837 29047 30895 29053
rect 31478 29044 31484 29096
rect 31536 29044 31542 29096
rect 32416 29084 32444 29115
rect 33042 29112 33048 29124
rect 33100 29112 33106 29164
rect 33134 29112 33140 29164
rect 33192 29152 33198 29164
rect 33796 29161 33824 29192
rect 34054 29180 34060 29192
rect 34112 29180 34118 29232
rect 34330 29180 34336 29232
rect 34388 29229 34394 29232
rect 34388 29223 34451 29229
rect 34388 29189 34405 29223
rect 34439 29189 34451 29223
rect 34388 29183 34451 29189
rect 34609 29223 34667 29229
rect 34609 29189 34621 29223
rect 34655 29189 34667 29223
rect 34609 29183 34667 29189
rect 35345 29223 35403 29229
rect 35345 29189 35357 29223
rect 35391 29220 35403 29223
rect 36814 29220 36820 29232
rect 35391 29192 35848 29220
rect 35391 29189 35403 29192
rect 35345 29183 35403 29189
rect 34388 29180 34394 29183
rect 33689 29155 33747 29161
rect 33689 29152 33701 29155
rect 33192 29124 33701 29152
rect 33192 29112 33198 29124
rect 33689 29121 33701 29124
rect 33735 29121 33747 29155
rect 33689 29115 33747 29121
rect 33781 29155 33839 29161
rect 33781 29121 33793 29155
rect 33827 29121 33839 29155
rect 33781 29115 33839 29121
rect 33410 29084 33416 29096
rect 31726 29056 33416 29084
rect 25777 28979 25835 28985
rect 26436 28988 28120 29016
rect 26436 28960 26464 28988
rect 28166 28976 28172 29028
rect 28224 28976 28230 29028
rect 29730 28976 29736 29028
rect 29788 29016 29794 29028
rect 30561 29019 30619 29025
rect 30561 29016 30573 29019
rect 29788 28988 30573 29016
rect 29788 28976 29794 28988
rect 30561 28985 30573 28988
rect 30607 28985 30619 29019
rect 30561 28979 30619 28985
rect 22465 28951 22523 28957
rect 22465 28948 22477 28951
rect 22428 28920 22477 28948
rect 22428 28908 22434 28920
rect 22465 28917 22477 28920
rect 22511 28948 22523 28951
rect 23290 28948 23296 28960
rect 22511 28920 23296 28948
rect 22511 28917 22523 28920
rect 22465 28911 22523 28917
rect 23290 28908 23296 28920
rect 23348 28908 23354 28960
rect 23385 28951 23443 28957
rect 23385 28917 23397 28951
rect 23431 28948 23443 28951
rect 23845 28951 23903 28957
rect 23845 28948 23857 28951
rect 23431 28920 23857 28948
rect 23431 28917 23443 28920
rect 23385 28911 23443 28917
rect 23845 28917 23857 28920
rect 23891 28917 23903 28951
rect 23845 28911 23903 28917
rect 25038 28908 25044 28960
rect 25096 28908 25102 28960
rect 26418 28908 26424 28960
rect 26476 28908 26482 28960
rect 27062 28908 27068 28960
rect 27120 28948 27126 28960
rect 27249 28951 27307 28957
rect 27249 28948 27261 28951
rect 27120 28920 27261 28948
rect 27120 28908 27126 28920
rect 27249 28917 27261 28920
rect 27295 28917 27307 28951
rect 27249 28911 27307 28917
rect 30374 28908 30380 28960
rect 30432 28948 30438 28960
rect 31726 28948 31754 29056
rect 33410 29044 33416 29056
rect 33468 29044 33474 29096
rect 33594 29016 33600 29028
rect 32968 28988 33600 29016
rect 30432 28920 31754 28948
rect 32769 28951 32827 28957
rect 30432 28908 30438 28920
rect 32769 28917 32781 28951
rect 32815 28948 32827 28951
rect 32968 28948 32996 28988
rect 33594 28976 33600 28988
rect 33652 28976 33658 29028
rect 32815 28920 32996 28948
rect 33704 28948 33732 29115
rect 33870 29112 33876 29164
rect 33928 29152 33934 29164
rect 34624 29152 34652 29183
rect 33928 29124 34652 29152
rect 33928 29112 33934 29124
rect 34882 29112 34888 29164
rect 34940 29152 34946 29164
rect 35161 29155 35219 29161
rect 35161 29152 35173 29155
rect 34940 29124 35173 29152
rect 34940 29112 34946 29124
rect 35161 29121 35173 29124
rect 35207 29121 35219 29155
rect 35161 29115 35219 29121
rect 35437 29155 35495 29161
rect 35437 29121 35449 29155
rect 35483 29152 35495 29155
rect 35526 29152 35532 29164
rect 35483 29124 35532 29152
rect 35483 29121 35495 29124
rect 35437 29115 35495 29121
rect 33965 29087 34023 29093
rect 33965 29053 33977 29087
rect 34011 29084 34023 29087
rect 34422 29084 34428 29096
rect 34011 29056 34428 29084
rect 34011 29053 34023 29056
rect 33965 29047 34023 29053
rect 34422 29044 34428 29056
rect 34480 29044 34486 29096
rect 35176 29084 35204 29115
rect 35526 29112 35532 29124
rect 35584 29112 35590 29164
rect 35820 29161 35848 29192
rect 36096 29192 36820 29220
rect 35805 29155 35863 29161
rect 35805 29121 35817 29155
rect 35851 29152 35863 29155
rect 35894 29152 35900 29164
rect 35851 29124 35900 29152
rect 35851 29121 35863 29124
rect 35805 29115 35863 29121
rect 35894 29112 35900 29124
rect 35952 29112 35958 29164
rect 36096 29161 36124 29192
rect 36814 29180 36820 29192
rect 36872 29180 36878 29232
rect 37553 29223 37611 29229
rect 37553 29220 37565 29223
rect 37292 29192 37565 29220
rect 36081 29155 36139 29161
rect 36081 29121 36093 29155
rect 36127 29121 36139 29155
rect 36081 29115 36139 29121
rect 36170 29112 36176 29164
rect 36228 29112 36234 29164
rect 37292 29152 37320 29192
rect 37553 29189 37565 29192
rect 37599 29189 37611 29223
rect 39942 29220 39948 29232
rect 38778 29192 39948 29220
rect 37553 29183 37611 29189
rect 39942 29180 39948 29192
rect 40000 29180 40006 29232
rect 40328 29192 41414 29220
rect 40328 29161 40356 29192
rect 36372 29124 37320 29152
rect 39669 29155 39727 29161
rect 35618 29084 35624 29096
rect 35176 29056 35624 29084
rect 35618 29044 35624 29056
rect 35676 29044 35682 29096
rect 36372 29093 36400 29124
rect 39669 29121 39681 29155
rect 39715 29121 39727 29155
rect 39669 29115 39727 29121
rect 40313 29155 40371 29161
rect 40313 29121 40325 29155
rect 40359 29121 40371 29155
rect 41386 29152 41414 29192
rect 41874 29152 41880 29164
rect 41386 29124 41880 29152
rect 40313 29115 40371 29121
rect 36357 29087 36415 29093
rect 36357 29053 36369 29087
rect 36403 29053 36415 29087
rect 36357 29047 36415 29053
rect 36446 29044 36452 29096
rect 36504 29084 36510 29096
rect 36814 29084 36820 29096
rect 36504 29056 36820 29084
rect 36504 29044 36510 29056
rect 36814 29044 36820 29056
rect 36872 29044 36878 29096
rect 37277 29087 37335 29093
rect 37277 29053 37289 29087
rect 37323 29084 37335 29087
rect 37918 29084 37924 29096
rect 37323 29056 37924 29084
rect 37323 29053 37335 29056
rect 37277 29047 37335 29053
rect 37918 29044 37924 29056
rect 37976 29084 37982 29096
rect 39684 29084 39712 29115
rect 41874 29112 41880 29124
rect 41932 29112 41938 29164
rect 40126 29084 40132 29096
rect 37976 29056 40132 29084
rect 37976 29044 37982 29056
rect 40126 29044 40132 29056
rect 40184 29084 40190 29096
rect 40402 29084 40408 29096
rect 40184 29056 40408 29084
rect 40184 29044 40190 29056
rect 40402 29044 40408 29056
rect 40460 29044 40466 29096
rect 40865 29087 40923 29093
rect 40865 29053 40877 29087
rect 40911 29084 40923 29087
rect 41417 29087 41475 29093
rect 41417 29084 41429 29087
rect 40911 29056 41429 29084
rect 40911 29053 40923 29056
rect 40865 29047 40923 29053
rect 41417 29053 41429 29056
rect 41463 29053 41475 29087
rect 41417 29047 41475 29053
rect 41509 29087 41567 29093
rect 41509 29053 41521 29087
rect 41555 29053 41567 29087
rect 41509 29047 41567 29053
rect 34146 28976 34152 29028
rect 34204 28976 34210 29028
rect 34238 28976 34244 29028
rect 34296 28976 34302 29028
rect 35250 28976 35256 29028
rect 35308 29016 35314 29028
rect 35802 29016 35808 29028
rect 35308 28988 35808 29016
rect 35308 28976 35314 28988
rect 35802 28976 35808 28988
rect 35860 29016 35866 29028
rect 35897 29019 35955 29025
rect 35897 29016 35909 29019
rect 35860 28988 35909 29016
rect 35860 28976 35866 28988
rect 35897 28985 35909 28988
rect 35943 28985 35955 29019
rect 35897 28979 35955 28985
rect 35986 28976 35992 29028
rect 36044 29016 36050 29028
rect 36906 29016 36912 29028
rect 36044 28988 36912 29016
rect 36044 28976 36050 28988
rect 36906 28976 36912 28988
rect 36964 28976 36970 29028
rect 39022 28976 39028 29028
rect 39080 28976 39086 29028
rect 39850 28976 39856 29028
rect 39908 29016 39914 29028
rect 39908 28988 40632 29016
rect 39908 28976 39914 28988
rect 34425 28951 34483 28957
rect 34425 28948 34437 28951
rect 33704 28920 34437 28948
rect 32815 28917 32827 28920
rect 32769 28911 32827 28917
rect 34425 28917 34437 28920
rect 34471 28917 34483 28951
rect 34425 28911 34483 28917
rect 34790 28908 34796 28960
rect 34848 28948 34854 28960
rect 34977 28951 35035 28957
rect 34977 28948 34989 28951
rect 34848 28920 34989 28948
rect 34848 28908 34854 28920
rect 34977 28917 34989 28920
rect 35023 28917 35035 28951
rect 40604 28948 40632 28988
rect 40678 28976 40684 29028
rect 40736 29016 40742 29028
rect 40957 29019 41015 29025
rect 40957 29016 40969 29019
rect 40736 28988 40969 29016
rect 40736 28976 40742 28988
rect 40957 28985 40969 28988
rect 41003 28985 41015 29019
rect 41524 29016 41552 29047
rect 40957 28979 41015 28985
rect 41064 28988 41552 29016
rect 41064 28948 41092 28988
rect 42058 28976 42064 29028
rect 42116 28976 42122 29028
rect 40604 28920 41092 28948
rect 34977 28911 35035 28917
rect 1104 28858 42504 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 42504 28858
rect 1104 28784 42504 28806
rect 3145 28747 3203 28753
rect 3145 28713 3157 28747
rect 3191 28744 3203 28747
rect 3602 28744 3608 28756
rect 3191 28716 3608 28744
rect 3191 28713 3203 28716
rect 3145 28707 3203 28713
rect 3602 28704 3608 28716
rect 3660 28704 3666 28756
rect 4709 28747 4767 28753
rect 4709 28713 4721 28747
rect 4755 28744 4767 28747
rect 4798 28744 4804 28756
rect 4755 28716 4804 28744
rect 4755 28713 4767 28716
rect 4709 28707 4767 28713
rect 4798 28704 4804 28716
rect 4856 28704 4862 28756
rect 4893 28747 4951 28753
rect 4893 28713 4905 28747
rect 4939 28744 4951 28747
rect 5350 28744 5356 28756
rect 4939 28716 5356 28744
rect 4939 28713 4951 28716
rect 4893 28707 4951 28713
rect 3050 28636 3056 28688
rect 3108 28676 3114 28688
rect 3329 28679 3387 28685
rect 3329 28676 3341 28679
rect 3108 28648 3341 28676
rect 3108 28636 3114 28648
rect 3329 28645 3341 28648
rect 3375 28645 3387 28679
rect 3329 28639 3387 28645
rect 3694 28636 3700 28688
rect 3752 28676 3758 28688
rect 3789 28679 3847 28685
rect 3789 28676 3801 28679
rect 3752 28648 3801 28676
rect 3752 28636 3758 28648
rect 3789 28645 3801 28648
rect 3835 28645 3847 28679
rect 4908 28676 4936 28707
rect 5350 28704 5356 28716
rect 5408 28704 5414 28756
rect 5994 28704 6000 28756
rect 6052 28744 6058 28756
rect 6089 28747 6147 28753
rect 6089 28744 6101 28747
rect 6052 28716 6101 28744
rect 6052 28704 6058 28716
rect 6089 28713 6101 28716
rect 6135 28713 6147 28747
rect 6089 28707 6147 28713
rect 6457 28747 6515 28753
rect 6457 28713 6469 28747
rect 6503 28744 6515 28747
rect 6822 28744 6828 28756
rect 6503 28716 6828 28744
rect 6503 28713 6515 28716
rect 6457 28707 6515 28713
rect 6822 28704 6828 28716
rect 6880 28704 6886 28756
rect 7466 28704 7472 28756
rect 7524 28744 7530 28756
rect 8205 28747 8263 28753
rect 8205 28744 8217 28747
rect 7524 28716 8217 28744
rect 7524 28704 7530 28716
rect 8205 28713 8217 28716
rect 8251 28744 8263 28747
rect 10870 28744 10876 28756
rect 8251 28716 10876 28744
rect 8251 28713 8263 28716
rect 8205 28707 8263 28713
rect 10870 28704 10876 28716
rect 10928 28704 10934 28756
rect 13173 28747 13231 28753
rect 13173 28713 13185 28747
rect 13219 28744 13231 28747
rect 13538 28744 13544 28756
rect 13219 28716 13544 28744
rect 13219 28713 13231 28716
rect 13173 28707 13231 28713
rect 13538 28704 13544 28716
rect 13596 28704 13602 28756
rect 13906 28704 13912 28756
rect 13964 28704 13970 28756
rect 17954 28704 17960 28756
rect 18012 28744 18018 28756
rect 18049 28747 18107 28753
rect 18049 28744 18061 28747
rect 18012 28716 18061 28744
rect 18012 28704 18018 28716
rect 18049 28713 18061 28716
rect 18095 28713 18107 28747
rect 18049 28707 18107 28713
rect 18598 28704 18604 28756
rect 18656 28744 18662 28756
rect 19242 28744 19248 28756
rect 18656 28716 19248 28744
rect 18656 28704 18662 28716
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 21266 28704 21272 28756
rect 21324 28704 21330 28756
rect 21358 28704 21364 28756
rect 21416 28744 21422 28756
rect 21453 28747 21511 28753
rect 21453 28744 21465 28747
rect 21416 28716 21465 28744
rect 21416 28704 21422 28716
rect 21453 28713 21465 28716
rect 21499 28713 21511 28747
rect 21453 28707 21511 28713
rect 21818 28704 21824 28756
rect 21876 28744 21882 28756
rect 22281 28747 22339 28753
rect 22281 28744 22293 28747
rect 21876 28716 22293 28744
rect 21876 28704 21882 28716
rect 22281 28713 22293 28716
rect 22327 28713 22339 28747
rect 22281 28707 22339 28713
rect 22554 28704 22560 28756
rect 22612 28704 22618 28756
rect 22833 28747 22891 28753
rect 22833 28713 22845 28747
rect 22879 28744 22891 28747
rect 23106 28744 23112 28756
rect 22879 28716 23112 28744
rect 22879 28713 22891 28716
rect 22833 28707 22891 28713
rect 23106 28704 23112 28716
rect 23164 28704 23170 28756
rect 23658 28704 23664 28756
rect 23716 28704 23722 28756
rect 25685 28747 25743 28753
rect 25685 28713 25697 28747
rect 25731 28744 25743 28747
rect 25774 28744 25780 28756
rect 25731 28716 25780 28744
rect 25731 28713 25743 28716
rect 25685 28707 25743 28713
rect 25774 28704 25780 28716
rect 25832 28704 25838 28756
rect 26142 28704 26148 28756
rect 26200 28744 26206 28756
rect 29270 28744 29276 28756
rect 26200 28716 29276 28744
rect 26200 28704 26206 28716
rect 29270 28704 29276 28716
rect 29328 28704 29334 28756
rect 29822 28704 29828 28756
rect 29880 28744 29886 28756
rect 30193 28747 30251 28753
rect 30193 28744 30205 28747
rect 29880 28716 30205 28744
rect 29880 28704 29886 28716
rect 30193 28713 30205 28716
rect 30239 28713 30251 28747
rect 30193 28707 30251 28713
rect 30650 28704 30656 28756
rect 30708 28704 30714 28756
rect 30742 28704 30748 28756
rect 30800 28744 30806 28756
rect 31018 28744 31024 28756
rect 30800 28716 31024 28744
rect 30800 28704 30806 28716
rect 31018 28704 31024 28716
rect 31076 28704 31082 28756
rect 34330 28704 34336 28756
rect 34388 28744 34394 28756
rect 34425 28747 34483 28753
rect 34425 28744 34437 28747
rect 34388 28716 34437 28744
rect 34388 28704 34394 28716
rect 34425 28713 34437 28716
rect 34471 28713 34483 28747
rect 34425 28707 34483 28713
rect 34790 28704 34796 28756
rect 34848 28744 34854 28756
rect 35161 28747 35219 28753
rect 35161 28744 35173 28747
rect 34848 28716 35173 28744
rect 34848 28704 34854 28716
rect 35161 28713 35173 28716
rect 35207 28713 35219 28747
rect 35161 28707 35219 28713
rect 36081 28747 36139 28753
rect 36081 28713 36093 28747
rect 36127 28744 36139 28747
rect 36170 28744 36176 28756
rect 36127 28716 36176 28744
rect 36127 28713 36139 28716
rect 36081 28707 36139 28713
rect 36170 28704 36176 28716
rect 36228 28704 36234 28756
rect 41874 28704 41880 28756
rect 41932 28744 41938 28756
rect 42153 28747 42211 28753
rect 42153 28744 42165 28747
rect 41932 28716 42165 28744
rect 41932 28704 41938 28716
rect 42153 28713 42165 28716
rect 42199 28713 42211 28747
rect 42153 28707 42211 28713
rect 3789 28639 3847 28645
rect 4448 28648 4936 28676
rect 1394 28568 1400 28620
rect 1452 28568 1458 28620
rect 1673 28611 1731 28617
rect 1673 28577 1685 28611
rect 1719 28608 1731 28611
rect 2038 28608 2044 28620
rect 1719 28580 2044 28608
rect 1719 28577 1731 28580
rect 1673 28571 1731 28577
rect 2038 28568 2044 28580
rect 2096 28568 2102 28620
rect 3418 28568 3424 28620
rect 3476 28608 3482 28620
rect 4065 28611 4123 28617
rect 4065 28608 4077 28611
rect 3476 28580 4077 28608
rect 3476 28568 3482 28580
rect 4065 28577 4077 28580
rect 4111 28577 4123 28611
rect 4065 28571 4123 28577
rect 2774 28500 2780 28552
rect 2832 28500 2838 28552
rect 3513 28543 3571 28549
rect 3513 28509 3525 28543
rect 3559 28509 3571 28543
rect 3513 28503 3571 28509
rect 3528 28472 3556 28503
rect 4154 28500 4160 28552
rect 4212 28500 4218 28552
rect 4448 28472 4476 28648
rect 5074 28636 5080 28688
rect 5132 28676 5138 28688
rect 5534 28676 5540 28688
rect 5132 28648 5540 28676
rect 5132 28636 5138 28648
rect 5534 28636 5540 28648
rect 5592 28636 5598 28688
rect 10965 28679 11023 28685
rect 10965 28645 10977 28679
rect 11011 28676 11023 28679
rect 11974 28676 11980 28688
rect 11011 28648 11980 28676
rect 11011 28645 11023 28648
rect 10965 28639 11023 28645
rect 11974 28636 11980 28648
rect 12032 28676 12038 28688
rect 12032 28648 12434 28676
rect 12032 28636 12038 28648
rect 4798 28568 4804 28620
rect 4856 28608 4862 28620
rect 9217 28611 9275 28617
rect 4856 28580 6132 28608
rect 4856 28568 4862 28580
rect 4525 28543 4583 28549
rect 4525 28509 4537 28543
rect 4571 28540 4583 28543
rect 4614 28540 4620 28552
rect 4571 28512 4620 28540
rect 4571 28509 4583 28512
rect 4525 28503 4583 28509
rect 4614 28500 4620 28512
rect 4672 28500 4678 28552
rect 4709 28543 4767 28549
rect 4709 28509 4721 28543
rect 4755 28509 4767 28543
rect 4709 28503 4767 28509
rect 5077 28543 5135 28549
rect 5077 28509 5089 28543
rect 5123 28509 5135 28543
rect 5077 28503 5135 28509
rect 4724 28472 4752 28503
rect 4798 28472 4804 28484
rect 3528 28444 4476 28472
rect 4540 28444 4804 28472
rect 3602 28364 3608 28416
rect 3660 28404 3666 28416
rect 4540 28404 4568 28444
rect 4798 28432 4804 28444
rect 4856 28472 4862 28484
rect 5092 28472 5120 28503
rect 5166 28500 5172 28552
rect 5224 28500 5230 28552
rect 5445 28543 5503 28549
rect 5445 28509 5457 28543
rect 5491 28540 5503 28543
rect 5534 28540 5540 28552
rect 5491 28512 5540 28540
rect 5491 28509 5503 28512
rect 5445 28503 5503 28509
rect 5534 28500 5540 28512
rect 5592 28500 5598 28552
rect 6104 28549 6132 28580
rect 9217 28577 9229 28611
rect 9263 28608 9275 28611
rect 9490 28608 9496 28620
rect 9263 28580 9496 28608
rect 9263 28577 9275 28580
rect 9217 28571 9275 28577
rect 9490 28568 9496 28580
rect 9548 28568 9554 28620
rect 12406 28608 12434 28648
rect 12710 28636 12716 28688
rect 12768 28636 12774 28688
rect 14277 28679 14335 28685
rect 14277 28645 14289 28679
rect 14323 28676 14335 28679
rect 14642 28676 14648 28688
rect 14323 28648 14648 28676
rect 14323 28645 14335 28648
rect 14277 28639 14335 28645
rect 14642 28636 14648 28648
rect 14700 28636 14706 28688
rect 14860 28648 15056 28676
rect 14860 28608 14888 28648
rect 12406 28580 13860 28608
rect 6089 28543 6147 28549
rect 6089 28509 6101 28543
rect 6135 28509 6147 28543
rect 6089 28503 6147 28509
rect 6270 28500 6276 28552
rect 6328 28500 6334 28552
rect 7650 28500 7656 28552
rect 7708 28500 7714 28552
rect 11514 28500 11520 28552
rect 11572 28500 11578 28552
rect 12802 28500 12808 28552
rect 12860 28540 12866 28552
rect 13081 28543 13139 28549
rect 13081 28540 13093 28543
rect 12860 28512 13093 28540
rect 12860 28500 12866 28512
rect 13081 28509 13093 28512
rect 13127 28509 13139 28543
rect 13081 28503 13139 28509
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28509 13323 28543
rect 13265 28503 13323 28509
rect 13725 28543 13783 28549
rect 13725 28509 13737 28543
rect 13771 28509 13783 28543
rect 13725 28503 13783 28509
rect 4856 28444 5120 28472
rect 4856 28432 4862 28444
rect 3660 28376 4568 28404
rect 3660 28364 3666 28376
rect 4614 28364 4620 28416
rect 4672 28404 4678 28416
rect 5184 28404 5212 28500
rect 5261 28475 5319 28481
rect 5261 28441 5273 28475
rect 5307 28472 5319 28475
rect 5350 28472 5356 28484
rect 5307 28444 5356 28472
rect 5307 28441 5319 28444
rect 5261 28435 5319 28441
rect 5350 28432 5356 28444
rect 5408 28432 5414 28484
rect 9493 28475 9551 28481
rect 9493 28441 9505 28475
rect 9539 28441 9551 28475
rect 10962 28472 10968 28484
rect 10718 28444 10968 28472
rect 9493 28435 9551 28441
rect 4672 28376 5212 28404
rect 9508 28404 9536 28435
rect 10962 28432 10968 28444
rect 11020 28432 11026 28484
rect 11606 28432 11612 28484
rect 11664 28472 11670 28484
rect 12342 28472 12348 28484
rect 11664 28444 12348 28472
rect 11664 28432 11670 28444
rect 12342 28432 12348 28444
rect 12400 28432 12406 28484
rect 12894 28432 12900 28484
rect 12952 28432 12958 28484
rect 11514 28404 11520 28416
rect 9508 28376 11520 28404
rect 4672 28364 4678 28376
rect 11514 28364 11520 28376
rect 11572 28364 11578 28416
rect 12618 28364 12624 28416
rect 12676 28404 12682 28416
rect 13280 28404 13308 28503
rect 12676 28376 13308 28404
rect 13740 28404 13768 28503
rect 13832 28472 13860 28580
rect 14292 28580 14888 28608
rect 14292 28549 14320 28580
rect 13909 28543 13967 28549
rect 13909 28509 13921 28543
rect 13955 28540 13967 28543
rect 14277 28543 14335 28549
rect 14277 28540 14289 28543
rect 13955 28512 14289 28540
rect 13955 28509 13967 28512
rect 13909 28503 13967 28509
rect 14277 28509 14289 28512
rect 14323 28509 14335 28543
rect 14277 28503 14335 28509
rect 14550 28500 14556 28552
rect 14608 28500 14614 28552
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 14860 28540 14888 28580
rect 14918 28568 14924 28620
rect 14976 28568 14982 28620
rect 15028 28608 15056 28648
rect 18230 28636 18236 28688
rect 18288 28676 18294 28688
rect 18782 28676 18788 28688
rect 18288 28648 18788 28676
rect 18288 28636 18294 28648
rect 18782 28636 18788 28648
rect 18840 28636 18846 28688
rect 18877 28679 18935 28685
rect 18877 28645 18889 28679
rect 18923 28676 18935 28679
rect 20162 28676 20168 28688
rect 18923 28648 20168 28676
rect 18923 28645 18935 28648
rect 18877 28639 18935 28645
rect 15562 28608 15568 28620
rect 15028 28580 15568 28608
rect 15562 28568 15568 28580
rect 15620 28568 15626 28620
rect 16666 28568 16672 28620
rect 16724 28608 16730 28620
rect 16724 28580 17448 28608
rect 16724 28568 16730 28580
rect 17420 28552 17448 28580
rect 18506 28568 18512 28620
rect 18564 28608 18570 28620
rect 18693 28611 18751 28617
rect 18693 28608 18705 28611
rect 18564 28580 18705 28608
rect 18564 28568 18570 28580
rect 18693 28577 18705 28580
rect 18739 28577 18751 28611
rect 18693 28571 18751 28577
rect 17126 28540 17132 28552
rect 14691 28512 14888 28540
rect 16330 28512 17132 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 17126 28500 17132 28512
rect 17184 28500 17190 28552
rect 17402 28500 17408 28552
rect 17460 28540 17466 28552
rect 18138 28540 18144 28552
rect 17460 28512 18144 28540
rect 17460 28500 17466 28512
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 18230 28500 18236 28552
rect 18288 28500 18294 28552
rect 18417 28543 18475 28549
rect 18417 28509 18429 28543
rect 18463 28540 18475 28543
rect 18966 28540 18972 28552
rect 18463 28512 18972 28540
rect 18463 28509 18475 28512
rect 18417 28503 18475 28509
rect 18966 28500 18972 28512
rect 19024 28500 19030 28552
rect 19058 28500 19064 28552
rect 19116 28500 19122 28552
rect 13832 28444 14964 28472
rect 14458 28404 14464 28416
rect 13740 28376 14464 28404
rect 12676 28364 12682 28376
rect 14458 28364 14464 28376
rect 14516 28364 14522 28416
rect 14737 28407 14795 28413
rect 14737 28373 14749 28407
rect 14783 28404 14795 28407
rect 14826 28404 14832 28416
rect 14783 28376 14832 28404
rect 14783 28373 14795 28376
rect 14737 28367 14795 28373
rect 14826 28364 14832 28376
rect 14884 28364 14890 28416
rect 14936 28404 14964 28444
rect 15194 28432 15200 28484
rect 15252 28432 15258 28484
rect 16850 28432 16856 28484
rect 16908 28472 16914 28484
rect 16945 28475 17003 28481
rect 16945 28472 16957 28475
rect 16908 28444 16957 28472
rect 16908 28432 16914 28444
rect 16945 28441 16957 28444
rect 16991 28441 17003 28475
rect 16945 28435 17003 28441
rect 18046 28432 18052 28484
rect 18104 28472 18110 28484
rect 18325 28475 18383 28481
rect 18325 28472 18337 28475
rect 18104 28444 18337 28472
rect 18104 28432 18110 28444
rect 18325 28441 18337 28444
rect 18371 28441 18383 28475
rect 18325 28435 18383 28441
rect 18555 28475 18613 28481
rect 18555 28441 18567 28475
rect 18601 28472 18613 28475
rect 19168 28472 19196 28648
rect 20162 28636 20168 28648
rect 20220 28636 20226 28688
rect 21085 28679 21143 28685
rect 21085 28645 21097 28679
rect 21131 28676 21143 28679
rect 22002 28676 22008 28688
rect 21131 28648 22008 28676
rect 21131 28645 21143 28648
rect 21085 28639 21143 28645
rect 22002 28636 22008 28648
rect 22060 28676 22066 28688
rect 23474 28676 23480 28688
rect 22060 28648 22508 28676
rect 22060 28636 22066 28648
rect 22186 28608 22192 28620
rect 21192 28580 22192 28608
rect 19426 28500 19432 28552
rect 19484 28500 19490 28552
rect 20806 28500 20812 28552
rect 20864 28540 20870 28552
rect 21192 28549 21220 28580
rect 22186 28568 22192 28580
rect 22244 28568 22250 28620
rect 20993 28543 21051 28549
rect 20993 28540 21005 28543
rect 20864 28512 21005 28540
rect 20864 28500 20870 28512
rect 20993 28509 21005 28512
rect 21039 28509 21051 28543
rect 20993 28503 21051 28509
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28509 21235 28543
rect 21821 28543 21879 28549
rect 21177 28503 21235 28509
rect 21284 28512 21588 28540
rect 18601 28444 19196 28472
rect 18601 28441 18613 28444
rect 18555 28435 18613 28441
rect 19610 28432 19616 28484
rect 19668 28432 19674 28484
rect 21008 28472 21036 28503
rect 21284 28472 21312 28512
rect 21560 28484 21588 28512
rect 21821 28509 21833 28543
rect 21867 28540 21879 28543
rect 21928 28540 22048 28542
rect 22370 28540 22376 28552
rect 21867 28514 22376 28540
rect 21867 28512 21956 28514
rect 22020 28512 22376 28514
rect 21867 28509 21879 28512
rect 21821 28503 21879 28509
rect 22370 28500 22376 28512
rect 22428 28500 22434 28552
rect 22480 28549 22508 28648
rect 22756 28648 23480 28676
rect 22756 28549 22784 28648
rect 23474 28636 23480 28648
rect 23532 28676 23538 28688
rect 24302 28676 24308 28688
rect 23532 28648 24308 28676
rect 23532 28636 23538 28648
rect 24302 28636 24308 28648
rect 24360 28636 24366 28688
rect 24394 28636 24400 28688
rect 24452 28676 24458 28688
rect 26050 28676 26056 28688
rect 24452 28648 26056 28676
rect 24452 28636 24458 28648
rect 26050 28636 26056 28648
rect 26108 28636 26114 28688
rect 26418 28636 26424 28688
rect 26476 28676 26482 28688
rect 27157 28679 27215 28685
rect 27157 28676 27169 28679
rect 26476 28648 27169 28676
rect 26476 28636 26482 28648
rect 27157 28645 27169 28648
rect 27203 28645 27215 28679
rect 30558 28676 30564 28688
rect 27157 28639 27215 28645
rect 27264 28648 30564 28676
rect 24118 28568 24124 28620
rect 24176 28568 24182 28620
rect 26329 28611 26387 28617
rect 26329 28577 26341 28611
rect 26375 28608 26387 28611
rect 26878 28608 26884 28620
rect 26375 28580 26884 28608
rect 26375 28577 26387 28580
rect 26329 28571 26387 28577
rect 26878 28568 26884 28580
rect 26936 28608 26942 28620
rect 27264 28608 27292 28648
rect 30558 28636 30564 28648
rect 30616 28636 30622 28688
rect 31202 28636 31208 28688
rect 31260 28676 31266 28688
rect 31389 28679 31447 28685
rect 31389 28676 31401 28679
rect 31260 28648 31401 28676
rect 31260 28636 31266 28648
rect 31389 28645 31401 28648
rect 31435 28645 31447 28679
rect 31389 28639 31447 28645
rect 32030 28636 32036 28688
rect 32088 28676 32094 28688
rect 34698 28676 34704 28688
rect 32088 28648 34704 28676
rect 32088 28636 32094 28648
rect 34698 28636 34704 28648
rect 34756 28676 34762 28688
rect 35526 28676 35532 28688
rect 34756 28648 35532 28676
rect 34756 28636 34762 28648
rect 35526 28636 35532 28648
rect 35584 28676 35590 28688
rect 35621 28679 35679 28685
rect 35621 28676 35633 28679
rect 35584 28648 35633 28676
rect 35584 28636 35590 28648
rect 35621 28645 35633 28648
rect 35667 28645 35679 28679
rect 35621 28639 35679 28645
rect 26936 28580 27292 28608
rect 26936 28568 26942 28580
rect 28718 28568 28724 28620
rect 28776 28608 28782 28620
rect 28776 28580 30052 28608
rect 28776 28568 28782 28580
rect 22465 28543 22523 28549
rect 22465 28509 22477 28543
rect 22511 28509 22523 28543
rect 22465 28503 22523 28509
rect 22741 28543 22799 28549
rect 22741 28509 22753 28543
rect 22787 28509 22799 28543
rect 22741 28503 22799 28509
rect 22925 28543 22983 28549
rect 22925 28509 22937 28543
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 21008 28444 21312 28472
rect 21450 28432 21456 28484
rect 21508 28432 21514 28484
rect 21542 28432 21548 28484
rect 21600 28472 21606 28484
rect 21913 28475 21971 28481
rect 21913 28472 21925 28475
rect 21600 28444 21925 28472
rect 21600 28432 21606 28444
rect 21913 28441 21925 28444
rect 21959 28441 21971 28475
rect 21913 28435 21971 28441
rect 22097 28475 22155 28481
rect 22097 28441 22109 28475
rect 22143 28472 22155 28475
rect 22186 28472 22192 28484
rect 22143 28444 22192 28472
rect 22143 28441 22155 28444
rect 22097 28435 22155 28441
rect 22186 28432 22192 28444
rect 22244 28432 22250 28484
rect 22756 28404 22784 28503
rect 14936 28376 22784 28404
rect 22940 28404 22968 28503
rect 23014 28500 23020 28552
rect 23072 28500 23078 28552
rect 23106 28500 23112 28552
rect 23164 28540 23170 28552
rect 23201 28543 23259 28549
rect 23201 28540 23213 28543
rect 23164 28512 23213 28540
rect 23164 28500 23170 28512
rect 23201 28509 23213 28512
rect 23247 28509 23259 28543
rect 23201 28503 23259 28509
rect 23290 28500 23296 28552
rect 23348 28500 23354 28552
rect 23382 28500 23388 28552
rect 23440 28500 23446 28552
rect 23937 28543 23995 28549
rect 23937 28509 23949 28543
rect 23983 28540 23995 28543
rect 24136 28540 24164 28568
rect 30024 28552 30052 28580
rect 30098 28568 30104 28620
rect 30156 28608 30162 28620
rect 30742 28608 30748 28620
rect 30800 28617 30806 28620
rect 30156 28580 30604 28608
rect 30709 28580 30748 28608
rect 30156 28568 30162 28580
rect 23983 28512 24164 28540
rect 23983 28509 23995 28512
rect 23937 28503 23995 28509
rect 23032 28472 23060 28500
rect 23753 28475 23811 28481
rect 23753 28472 23765 28475
rect 23032 28444 23765 28472
rect 23753 28441 23765 28444
rect 23799 28441 23811 28475
rect 23753 28435 23811 28441
rect 23952 28404 23980 28503
rect 25682 28500 25688 28552
rect 25740 28540 25746 28552
rect 25869 28543 25927 28549
rect 25869 28540 25881 28543
rect 25740 28512 25881 28540
rect 25740 28500 25746 28512
rect 25869 28509 25881 28512
rect 25915 28509 25927 28543
rect 25869 28503 25927 28509
rect 25958 28500 25964 28552
rect 26016 28540 26022 28552
rect 26145 28543 26203 28549
rect 26145 28540 26157 28543
rect 26016 28512 26157 28540
rect 26016 28500 26022 28512
rect 26145 28509 26157 28512
rect 26191 28509 26203 28543
rect 26145 28503 26203 28509
rect 26510 28500 26516 28552
rect 26568 28500 26574 28552
rect 27062 28500 27068 28552
rect 27120 28500 27126 28552
rect 27614 28540 27620 28552
rect 27356 28512 27620 28540
rect 24121 28475 24179 28481
rect 24121 28441 24133 28475
rect 24167 28472 24179 28475
rect 24302 28472 24308 28484
rect 24167 28444 24308 28472
rect 24167 28441 24179 28444
rect 24121 28435 24179 28441
rect 24302 28432 24308 28444
rect 24360 28432 24366 28484
rect 26326 28432 26332 28484
rect 26384 28472 26390 28484
rect 27356 28481 27384 28512
rect 27614 28500 27620 28512
rect 27672 28500 27678 28552
rect 27706 28500 27712 28552
rect 27764 28540 27770 28552
rect 29549 28543 29607 28549
rect 29549 28540 29561 28543
rect 27764 28512 29561 28540
rect 27764 28500 27770 28512
rect 26605 28475 26663 28481
rect 26605 28472 26617 28475
rect 26384 28444 26617 28472
rect 26384 28432 26390 28444
rect 26605 28441 26617 28444
rect 26651 28441 26663 28475
rect 27341 28475 27399 28481
rect 27341 28472 27353 28475
rect 26605 28435 26663 28441
rect 26712 28444 27353 28472
rect 22940 28376 23980 28404
rect 26050 28364 26056 28416
rect 26108 28364 26114 28416
rect 26510 28364 26516 28416
rect 26568 28404 26574 28416
rect 26712 28404 26740 28444
rect 27341 28441 27353 28444
rect 27387 28441 27399 28475
rect 27341 28435 27399 28441
rect 27522 28432 27528 28484
rect 27580 28472 27586 28484
rect 29181 28475 29239 28481
rect 29181 28472 29193 28475
rect 27580 28444 29193 28472
rect 27580 28432 27586 28444
rect 29181 28441 29193 28444
rect 29227 28441 29239 28475
rect 29181 28435 29239 28441
rect 26568 28376 26740 28404
rect 26568 28364 26574 28376
rect 26786 28364 26792 28416
rect 26844 28404 26850 28416
rect 26973 28407 27031 28413
rect 26973 28404 26985 28407
rect 26844 28376 26985 28404
rect 26844 28364 26850 28376
rect 26973 28373 26985 28376
rect 27019 28373 27031 28407
rect 26973 28367 27031 28373
rect 27065 28407 27123 28413
rect 27065 28373 27077 28407
rect 27111 28404 27123 28407
rect 28810 28404 28816 28416
rect 27111 28376 28816 28404
rect 27111 28373 27123 28376
rect 27065 28367 27123 28373
rect 28810 28364 28816 28376
rect 28868 28364 28874 28416
rect 29288 28404 29316 28512
rect 29549 28509 29561 28512
rect 29595 28509 29607 28543
rect 29549 28503 29607 28509
rect 29638 28500 29644 28552
rect 29696 28540 29702 28552
rect 29696 28512 29741 28540
rect 29696 28500 29702 28512
rect 29914 28500 29920 28552
rect 29972 28500 29978 28552
rect 30006 28500 30012 28552
rect 30064 28549 30070 28552
rect 30064 28540 30072 28549
rect 30064 28512 30109 28540
rect 30064 28503 30072 28512
rect 30064 28500 30070 28503
rect 30282 28500 30288 28552
rect 30340 28500 30346 28552
rect 30466 28500 30472 28552
rect 30524 28500 30530 28552
rect 30576 28540 30604 28580
rect 30742 28568 30748 28580
rect 30800 28571 30809 28617
rect 30800 28568 30806 28571
rect 31110 28568 31116 28620
rect 31168 28608 31174 28620
rect 31297 28611 31355 28617
rect 31297 28608 31309 28611
rect 31168 28580 31309 28608
rect 31168 28568 31174 28580
rect 31297 28577 31309 28580
rect 31343 28577 31355 28611
rect 31297 28571 31355 28577
rect 34054 28568 34060 28620
rect 34112 28568 34118 28620
rect 34422 28608 34428 28620
rect 34256 28580 34428 28608
rect 31573 28543 31631 28549
rect 30576 28512 30788 28540
rect 29365 28475 29423 28481
rect 29365 28441 29377 28475
rect 29411 28472 29423 28475
rect 29825 28475 29883 28481
rect 29825 28472 29837 28475
rect 29411 28444 29837 28472
rect 29411 28441 29423 28444
rect 29365 28435 29423 28441
rect 29825 28441 29837 28444
rect 29871 28472 29883 28475
rect 30650 28472 30656 28484
rect 29871 28444 30656 28472
rect 29871 28441 29883 28444
rect 29825 28435 29883 28441
rect 30650 28432 30656 28444
rect 30708 28432 30714 28484
rect 30760 28472 30788 28512
rect 31573 28509 31585 28543
rect 31619 28509 31631 28543
rect 31573 28503 31631 28509
rect 30837 28475 30895 28481
rect 30837 28472 30849 28475
rect 30760 28444 30849 28472
rect 30837 28441 30849 28444
rect 30883 28441 30895 28475
rect 30837 28435 30895 28441
rect 30926 28432 30932 28484
rect 30984 28472 30990 28484
rect 31037 28475 31095 28481
rect 31037 28472 31049 28475
rect 30984 28444 31049 28472
rect 30984 28432 30990 28444
rect 31037 28441 31049 28444
rect 31083 28441 31095 28475
rect 31588 28472 31616 28503
rect 31846 28500 31852 28552
rect 31904 28500 31910 28552
rect 32030 28500 32036 28552
rect 32088 28500 32094 28552
rect 34256 28549 34284 28580
rect 34422 28568 34428 28580
rect 34480 28608 34486 28620
rect 34793 28611 34851 28617
rect 34793 28608 34805 28611
rect 34480 28580 34805 28608
rect 34480 28568 34486 28580
rect 34793 28577 34805 28580
rect 34839 28577 34851 28611
rect 35437 28611 35495 28617
rect 35437 28608 35449 28611
rect 34793 28571 34851 28577
rect 35176 28580 35449 28608
rect 34241 28543 34299 28549
rect 34241 28509 34253 28543
rect 34287 28509 34299 28543
rect 34241 28503 34299 28509
rect 31941 28475 31999 28481
rect 31941 28472 31953 28475
rect 31588 28444 31953 28472
rect 31037 28435 31095 28441
rect 31941 28441 31953 28444
rect 31987 28441 31999 28475
rect 31941 28435 31999 28441
rect 34146 28432 34152 28484
rect 34204 28472 34210 28484
rect 34606 28472 34612 28484
rect 34204 28444 34612 28472
rect 34204 28432 34210 28444
rect 34606 28432 34612 28444
rect 34664 28472 34670 28484
rect 35176 28481 35204 28580
rect 35437 28577 35449 28580
rect 35483 28577 35495 28611
rect 35636 28608 35664 28639
rect 35636 28580 35848 28608
rect 35437 28571 35495 28577
rect 35710 28500 35716 28552
rect 35768 28500 35774 28552
rect 35820 28549 35848 28580
rect 37918 28568 37924 28620
rect 37976 28568 37982 28620
rect 40678 28568 40684 28620
rect 40736 28568 40742 28620
rect 35805 28543 35863 28549
rect 35805 28509 35817 28543
rect 35851 28509 35863 28543
rect 35805 28503 35863 28509
rect 35894 28500 35900 28552
rect 35952 28540 35958 28552
rect 36538 28540 36544 28552
rect 35952 28512 36544 28540
rect 35952 28500 35958 28512
rect 36538 28500 36544 28512
rect 36596 28500 36602 28552
rect 37642 28500 37648 28552
rect 37700 28500 37706 28552
rect 40126 28500 40132 28552
rect 40184 28540 40190 28552
rect 40405 28543 40463 28549
rect 40405 28540 40417 28543
rect 40184 28512 40417 28540
rect 40184 28500 40190 28512
rect 40405 28509 40417 28512
rect 40451 28509 40463 28543
rect 40405 28503 40463 28509
rect 35161 28475 35219 28481
rect 35161 28472 35173 28475
rect 34664 28444 35173 28472
rect 34664 28432 34670 28444
rect 35161 28441 35173 28444
rect 35207 28441 35219 28475
rect 35161 28435 35219 28441
rect 35437 28475 35495 28481
rect 35437 28441 35449 28475
rect 35483 28472 35495 28475
rect 36081 28475 36139 28481
rect 36081 28472 36093 28475
rect 35483 28444 36093 28472
rect 35483 28441 35495 28444
rect 35437 28435 35495 28441
rect 36081 28441 36093 28444
rect 36127 28441 36139 28475
rect 36081 28435 36139 28441
rect 37826 28432 37832 28484
rect 37884 28432 37890 28484
rect 38197 28475 38255 28481
rect 38197 28441 38209 28475
rect 38243 28441 38255 28475
rect 39942 28472 39948 28484
rect 39422 28444 39948 28472
rect 38197 28435 38255 28441
rect 30558 28404 30564 28416
rect 29288 28376 30564 28404
rect 30558 28364 30564 28376
rect 30616 28364 30622 28416
rect 31757 28407 31815 28413
rect 31757 28373 31769 28407
rect 31803 28404 31815 28407
rect 32306 28404 32312 28416
rect 31803 28376 32312 28404
rect 31803 28373 31815 28376
rect 31757 28367 31815 28373
rect 32306 28364 32312 28376
rect 32364 28364 32370 28416
rect 35342 28364 35348 28416
rect 35400 28364 35406 28416
rect 37461 28407 37519 28413
rect 37461 28373 37473 28407
rect 37507 28404 37519 28407
rect 38212 28404 38240 28435
rect 39942 28432 39948 28444
rect 40000 28432 40006 28484
rect 41690 28432 41696 28484
rect 41748 28432 41754 28484
rect 37507 28376 38240 28404
rect 37507 28373 37519 28376
rect 37461 28367 37519 28373
rect 38838 28364 38844 28416
rect 38896 28404 38902 28416
rect 39669 28407 39727 28413
rect 39669 28404 39681 28407
rect 38896 28376 39681 28404
rect 38896 28364 38902 28376
rect 39669 28373 39681 28376
rect 39715 28404 39727 28407
rect 41506 28404 41512 28416
rect 39715 28376 41512 28404
rect 39715 28373 39727 28376
rect 39669 28367 39727 28373
rect 41506 28364 41512 28376
rect 41564 28364 41570 28416
rect 1104 28314 42504 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 42504 28314
rect 1104 28240 42504 28262
rect 3602 28200 3608 28212
rect 1688 28172 3608 28200
rect 1688 28073 1716 28172
rect 3602 28160 3608 28172
rect 3660 28160 3666 28212
rect 3697 28203 3755 28209
rect 3697 28169 3709 28203
rect 3743 28200 3755 28203
rect 4154 28200 4160 28212
rect 3743 28172 4160 28200
rect 3743 28169 3755 28172
rect 3697 28163 3755 28169
rect 4154 28160 4160 28172
rect 4212 28160 4218 28212
rect 4798 28160 4804 28212
rect 4856 28200 4862 28212
rect 5074 28200 5080 28212
rect 4856 28172 5080 28200
rect 4856 28160 4862 28172
rect 5074 28160 5080 28172
rect 5132 28160 5138 28212
rect 5261 28203 5319 28209
rect 5261 28169 5273 28203
rect 5307 28200 5319 28203
rect 5350 28200 5356 28212
rect 5307 28172 5356 28200
rect 5307 28169 5319 28172
rect 5261 28163 5319 28169
rect 5350 28160 5356 28172
rect 5408 28160 5414 28212
rect 5626 28200 5632 28212
rect 5460 28172 5632 28200
rect 2774 28092 2780 28144
rect 2832 28092 2838 28144
rect 3510 28092 3516 28144
rect 3568 28132 3574 28144
rect 5460 28132 5488 28172
rect 5626 28160 5632 28172
rect 5684 28160 5690 28212
rect 9766 28160 9772 28212
rect 9824 28200 9830 28212
rect 10505 28203 10563 28209
rect 10505 28200 10517 28203
rect 9824 28172 10517 28200
rect 9824 28160 9830 28172
rect 10505 28169 10517 28172
rect 10551 28169 10563 28203
rect 10505 28163 10563 28169
rect 10870 28160 10876 28212
rect 10928 28160 10934 28212
rect 10965 28203 11023 28209
rect 10965 28169 10977 28203
rect 11011 28200 11023 28203
rect 11238 28200 11244 28212
rect 11011 28172 11244 28200
rect 11011 28169 11023 28172
rect 10965 28163 11023 28169
rect 11238 28160 11244 28172
rect 11296 28160 11302 28212
rect 11514 28160 11520 28212
rect 11572 28160 11578 28212
rect 11974 28160 11980 28212
rect 12032 28160 12038 28212
rect 13722 28160 13728 28212
rect 13780 28200 13786 28212
rect 14734 28200 14740 28212
rect 13780 28172 14740 28200
rect 13780 28160 13786 28172
rect 5718 28132 5724 28144
rect 3568 28104 5488 28132
rect 5552 28104 5724 28132
rect 3568 28092 3574 28104
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28033 1731 28067
rect 1673 28027 1731 28033
rect 4798 28024 4804 28076
rect 4856 28064 4862 28076
rect 5552 28073 5580 28104
rect 5718 28092 5724 28104
rect 5776 28132 5782 28144
rect 6086 28132 6092 28144
rect 5776 28104 6092 28132
rect 5776 28092 5782 28104
rect 6086 28092 6092 28104
rect 6144 28092 6150 28144
rect 9490 28132 9496 28144
rect 8956 28104 9496 28132
rect 5169 28067 5227 28073
rect 5169 28064 5181 28067
rect 4856 28036 5181 28064
rect 4856 28024 4862 28036
rect 5169 28033 5181 28036
rect 5215 28033 5227 28067
rect 5169 28027 5227 28033
rect 5537 28067 5595 28073
rect 5537 28033 5549 28067
rect 5583 28033 5595 28067
rect 5537 28027 5595 28033
rect 5629 28067 5687 28073
rect 5629 28033 5641 28067
rect 5675 28064 5687 28067
rect 6546 28064 6552 28076
rect 5675 28036 6552 28064
rect 5675 28033 5687 28036
rect 5629 28027 5687 28033
rect 6546 28024 6552 28036
rect 6604 28024 6610 28076
rect 8294 28024 8300 28076
rect 8352 28064 8358 28076
rect 8956 28073 8984 28104
rect 9490 28092 9496 28104
rect 9548 28132 9554 28144
rect 9548 28104 10456 28132
rect 9548 28092 9554 28104
rect 8674 28067 8732 28073
rect 8674 28064 8686 28067
rect 8352 28036 8686 28064
rect 8352 28024 8358 28036
rect 8674 28033 8686 28036
rect 8720 28033 8732 28067
rect 8674 28027 8732 28033
rect 8941 28067 8999 28073
rect 8941 28033 8953 28067
rect 8987 28033 8999 28067
rect 8941 28027 8999 28033
rect 9674 28024 9680 28076
rect 9732 28064 9738 28076
rect 10146 28067 10204 28073
rect 10146 28064 10158 28067
rect 9732 28036 10158 28064
rect 9732 28024 9738 28036
rect 10146 28033 10158 28036
rect 10192 28033 10204 28067
rect 10146 28027 10204 28033
rect 1394 27956 1400 28008
rect 1452 27996 1458 28008
rect 1949 27999 2007 28005
rect 1949 27996 1961 27999
rect 1452 27968 1961 27996
rect 1452 27956 1458 27968
rect 1949 27965 1961 27968
rect 1995 27965 2007 27999
rect 1949 27959 2007 27965
rect 2225 27999 2283 28005
rect 2225 27965 2237 27999
rect 2271 27996 2283 27999
rect 2866 27996 2872 28008
rect 2271 27968 2872 27996
rect 2271 27965 2283 27968
rect 2225 27959 2283 27965
rect 2866 27956 2872 27968
rect 2924 27956 2930 28008
rect 4706 27956 4712 28008
rect 4764 27996 4770 28008
rect 10428 28005 10456 28104
rect 12526 28092 12532 28144
rect 12584 28092 12590 28144
rect 14384 28132 14412 28172
rect 14734 28160 14740 28172
rect 14792 28200 14798 28212
rect 15013 28203 15071 28209
rect 14792 28172 14964 28200
rect 14792 28160 14798 28172
rect 14214 28104 14412 28132
rect 14458 28092 14464 28144
rect 14516 28132 14522 28144
rect 14645 28135 14703 28141
rect 14645 28132 14657 28135
rect 14516 28104 14657 28132
rect 14516 28092 14522 28104
rect 14645 28101 14657 28104
rect 14691 28101 14703 28135
rect 14845 28135 14903 28141
rect 14845 28132 14857 28135
rect 14645 28095 14703 28101
rect 14844 28101 14857 28132
rect 14891 28101 14903 28135
rect 14936 28132 14964 28172
rect 15013 28169 15025 28203
rect 15059 28200 15071 28203
rect 15194 28200 15200 28212
rect 15059 28172 15200 28200
rect 15059 28169 15071 28172
rect 15013 28163 15071 28169
rect 15194 28160 15200 28172
rect 15252 28160 15258 28212
rect 17954 28160 17960 28212
rect 18012 28200 18018 28212
rect 18322 28200 18328 28212
rect 18012 28172 18328 28200
rect 18012 28160 18018 28172
rect 18322 28160 18328 28172
rect 18380 28200 18386 28212
rect 18509 28203 18567 28209
rect 18509 28200 18521 28203
rect 18380 28172 18521 28200
rect 18380 28160 18386 28172
rect 18509 28169 18521 28172
rect 18555 28169 18567 28203
rect 18509 28163 18567 28169
rect 19518 28160 19524 28212
rect 19576 28200 19582 28212
rect 19981 28203 20039 28209
rect 19981 28200 19993 28203
rect 19576 28172 19993 28200
rect 19576 28160 19582 28172
rect 19981 28169 19993 28172
rect 20027 28169 20039 28203
rect 19981 28163 20039 28169
rect 23658 28160 23664 28212
rect 23716 28200 23722 28212
rect 28442 28200 28448 28212
rect 23716 28172 28448 28200
rect 23716 28160 23722 28172
rect 28442 28160 28448 28172
rect 28500 28160 28506 28212
rect 28629 28203 28687 28209
rect 28629 28169 28641 28203
rect 28675 28169 28687 28203
rect 28629 28163 28687 28169
rect 17126 28132 17132 28144
rect 14936 28104 17132 28132
rect 14844 28095 14903 28101
rect 11146 28024 11152 28076
rect 11204 28064 11210 28076
rect 11885 28067 11943 28073
rect 11885 28064 11897 28067
rect 11204 28036 11897 28064
rect 11204 28024 11210 28036
rect 11885 28033 11897 28036
rect 11931 28033 11943 28067
rect 11885 28027 11943 28033
rect 12434 28024 12440 28076
rect 12492 28024 12498 28076
rect 12618 28024 12624 28076
rect 12676 28024 12682 28076
rect 5261 27999 5319 28005
rect 5261 27996 5273 27999
rect 4764 27968 5273 27996
rect 4764 27956 4770 27968
rect 5261 27965 5273 27968
rect 5307 27965 5319 27999
rect 5261 27959 5319 27965
rect 10413 27999 10471 28005
rect 10413 27965 10425 27999
rect 10459 27996 10471 27999
rect 11057 27999 11115 28005
rect 10459 27968 10916 27996
rect 10459 27965 10471 27968
rect 10413 27959 10471 27965
rect 5166 27888 5172 27940
rect 5224 27928 5230 27940
rect 5534 27928 5540 27940
rect 5224 27900 5540 27928
rect 5224 27888 5230 27900
rect 5534 27888 5540 27900
rect 5592 27888 5598 27940
rect 10888 27872 10916 27968
rect 11057 27965 11069 27999
rect 11103 27996 11115 27999
rect 12066 27996 12072 28008
rect 11103 27968 12072 27996
rect 11103 27965 11115 27968
rect 11057 27959 11115 27965
rect 12066 27956 12072 27968
rect 12124 27956 12130 28008
rect 12342 27956 12348 28008
rect 12400 27996 12406 28008
rect 12713 27999 12771 28005
rect 12713 27996 12725 27999
rect 12400 27968 12725 27996
rect 12400 27956 12406 27968
rect 12713 27965 12725 27968
rect 12759 27965 12771 27999
rect 12713 27959 12771 27965
rect 12989 27999 13047 28005
rect 12989 27965 13001 27999
rect 13035 27996 13047 27999
rect 14458 27996 14464 28008
rect 13035 27968 14464 27996
rect 13035 27965 13047 27968
rect 12989 27959 13047 27965
rect 842 27820 848 27872
rect 900 27860 906 27872
rect 1489 27863 1547 27869
rect 1489 27860 1501 27863
rect 900 27832 1501 27860
rect 900 27820 906 27832
rect 1489 27829 1501 27832
rect 1535 27829 1547 27863
rect 1489 27823 1547 27829
rect 4982 27820 4988 27872
rect 5040 27820 5046 27872
rect 5074 27820 5080 27872
rect 5132 27860 5138 27872
rect 5445 27863 5503 27869
rect 5445 27860 5457 27863
rect 5132 27832 5457 27860
rect 5132 27820 5138 27832
rect 5445 27829 5457 27832
rect 5491 27860 5503 27863
rect 5721 27863 5779 27869
rect 5721 27860 5733 27863
rect 5491 27832 5733 27860
rect 5491 27829 5503 27832
rect 5445 27823 5503 27829
rect 5721 27829 5733 27832
rect 5767 27860 5779 27863
rect 5810 27860 5816 27872
rect 5767 27832 5816 27860
rect 5767 27829 5779 27832
rect 5721 27823 5779 27829
rect 5810 27820 5816 27832
rect 5868 27860 5874 27872
rect 6178 27860 6184 27872
rect 5868 27832 6184 27860
rect 5868 27820 5874 27832
rect 6178 27820 6184 27832
rect 6236 27820 6242 27872
rect 7561 27863 7619 27869
rect 7561 27829 7573 27863
rect 7607 27860 7619 27863
rect 7650 27860 7656 27872
rect 7607 27832 7656 27860
rect 7607 27829 7619 27832
rect 7561 27823 7619 27829
rect 7650 27820 7656 27832
rect 7708 27820 7714 27872
rect 9030 27820 9036 27872
rect 9088 27820 9094 27872
rect 10870 27820 10876 27872
rect 10928 27860 10934 27872
rect 11606 27860 11612 27872
rect 10928 27832 11612 27860
rect 10928 27820 10934 27832
rect 11606 27820 11612 27832
rect 11664 27820 11670 27872
rect 12728 27860 12756 27959
rect 14458 27956 14464 27968
rect 14516 27956 14522 28008
rect 14660 27996 14688 28095
rect 14844 28064 14872 28095
rect 17126 28092 17132 28104
rect 17184 28092 17190 28144
rect 18877 28135 18935 28141
rect 18877 28101 18889 28135
rect 18923 28132 18935 28135
rect 25038 28132 25044 28144
rect 18923 28104 20116 28132
rect 18923 28101 18935 28104
rect 18877 28095 18935 28101
rect 20088 28076 20116 28104
rect 24780 28104 25044 28132
rect 15010 28064 15016 28076
rect 14844 28036 15016 28064
rect 15010 28024 15016 28036
rect 15068 28024 15074 28076
rect 15381 28067 15439 28073
rect 15381 28033 15393 28067
rect 15427 28033 15439 28067
rect 15381 28027 15439 28033
rect 15102 27996 15108 28008
rect 14660 27968 15108 27996
rect 15102 27956 15108 27968
rect 15160 27956 15166 28008
rect 15396 27928 15424 28027
rect 18230 28024 18236 28076
rect 18288 28064 18294 28076
rect 18325 28067 18383 28073
rect 18325 28064 18337 28067
rect 18288 28036 18337 28064
rect 18288 28024 18294 28036
rect 18325 28033 18337 28036
rect 18371 28064 18383 28067
rect 18506 28064 18512 28076
rect 18371 28036 18512 28064
rect 18371 28033 18383 28036
rect 18325 28027 18383 28033
rect 18506 28024 18512 28036
rect 18564 28064 18570 28076
rect 18785 28067 18843 28073
rect 18785 28064 18797 28067
rect 18564 28036 18797 28064
rect 18564 28024 18570 28036
rect 18785 28033 18797 28036
rect 18831 28033 18843 28067
rect 18785 28027 18843 28033
rect 18969 28067 19027 28073
rect 18969 28033 18981 28067
rect 19015 28033 19027 28067
rect 18969 28027 19027 28033
rect 16850 27956 16856 28008
rect 16908 27996 16914 28008
rect 18141 27999 18199 28005
rect 18141 27996 18153 27999
rect 16908 27968 18153 27996
rect 16908 27956 16914 27968
rect 18141 27965 18153 27968
rect 18187 27996 18199 27999
rect 18414 27996 18420 28008
rect 18187 27968 18420 27996
rect 18187 27965 18199 27968
rect 18141 27959 18199 27965
rect 18414 27956 18420 27968
rect 18472 27996 18478 28008
rect 18984 27996 19012 28027
rect 19150 28024 19156 28076
rect 19208 28064 19214 28076
rect 19889 28067 19947 28073
rect 19889 28064 19901 28067
rect 19208 28036 19901 28064
rect 19208 28024 19214 28036
rect 19889 28033 19901 28036
rect 19935 28033 19947 28067
rect 19889 28027 19947 28033
rect 20070 28024 20076 28076
rect 20128 28064 20134 28076
rect 21634 28064 21640 28076
rect 20128 28036 21640 28064
rect 20128 28024 20134 28036
rect 21634 28024 21640 28036
rect 21692 28024 21698 28076
rect 23566 28024 23572 28076
rect 23624 28024 23630 28076
rect 23750 28024 23756 28076
rect 23808 28024 23814 28076
rect 24780 28073 24808 28104
rect 25038 28092 25044 28104
rect 25096 28092 25102 28144
rect 25501 28135 25559 28141
rect 25501 28101 25513 28135
rect 25547 28132 25559 28135
rect 26418 28132 26424 28144
rect 25547 28104 26424 28132
rect 25547 28101 25559 28104
rect 25501 28095 25559 28101
rect 26418 28092 26424 28104
rect 26476 28132 26482 28144
rect 27430 28132 27436 28144
rect 26476 28104 27436 28132
rect 26476 28092 26482 28104
rect 27430 28092 27436 28104
rect 27488 28092 27494 28144
rect 28644 28132 28672 28163
rect 28718 28160 28724 28212
rect 28776 28200 28782 28212
rect 28997 28203 29055 28209
rect 28997 28200 29009 28203
rect 28776 28172 29009 28200
rect 28776 28160 28782 28172
rect 28997 28169 29009 28172
rect 29043 28169 29055 28203
rect 28997 28163 29055 28169
rect 29641 28203 29699 28209
rect 29641 28169 29653 28203
rect 29687 28200 29699 28203
rect 30098 28200 30104 28212
rect 29687 28172 30104 28200
rect 29687 28169 29699 28172
rect 29641 28163 29699 28169
rect 30098 28160 30104 28172
rect 30156 28160 30162 28212
rect 30466 28160 30472 28212
rect 30524 28200 30530 28212
rect 30929 28203 30987 28209
rect 30929 28200 30941 28203
rect 30524 28172 30941 28200
rect 30524 28160 30530 28172
rect 30929 28169 30941 28172
rect 30975 28169 30987 28203
rect 33134 28200 33140 28212
rect 30929 28163 30987 28169
rect 31036 28172 33140 28200
rect 27632 28104 28580 28132
rect 28644 28104 29408 28132
rect 24765 28067 24823 28073
rect 24765 28033 24777 28067
rect 24811 28033 24823 28067
rect 24765 28027 24823 28033
rect 24857 28067 24915 28073
rect 24857 28033 24869 28067
rect 24903 28033 24915 28067
rect 24857 28027 24915 28033
rect 25133 28067 25191 28073
rect 25133 28033 25145 28067
rect 25179 28064 25191 28067
rect 25222 28064 25228 28076
rect 25179 28036 25228 28064
rect 25179 28033 25191 28036
rect 25133 28027 25191 28033
rect 18472 27968 19012 27996
rect 18472 27956 18478 27968
rect 19058 27956 19064 28008
rect 19116 27996 19122 28008
rect 23768 27996 23796 28024
rect 19116 27968 23796 27996
rect 24872 27996 24900 28027
rect 25222 28024 25228 28036
rect 25280 28024 25286 28076
rect 25314 28024 25320 28076
rect 25372 28064 25378 28076
rect 25409 28067 25467 28073
rect 25409 28064 25421 28067
rect 25372 28036 25421 28064
rect 25372 28024 25378 28036
rect 25409 28033 25421 28036
rect 25455 28033 25467 28067
rect 25409 28027 25467 28033
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 24872 27968 25268 27996
rect 19116 27956 19122 27968
rect 14476 27900 18644 27928
rect 13998 27860 14004 27872
rect 12728 27832 14004 27860
rect 13998 27820 14004 27832
rect 14056 27820 14062 27872
rect 14476 27869 14504 27900
rect 14461 27863 14519 27869
rect 14461 27829 14473 27863
rect 14507 27829 14519 27863
rect 14461 27823 14519 27829
rect 14826 27820 14832 27872
rect 14884 27820 14890 27872
rect 15102 27820 15108 27872
rect 15160 27860 15166 27872
rect 15197 27863 15255 27869
rect 15197 27860 15209 27863
rect 15160 27832 15209 27860
rect 15160 27820 15166 27832
rect 15197 27829 15209 27832
rect 15243 27829 15255 27863
rect 15197 27823 15255 27829
rect 15378 27820 15384 27872
rect 15436 27860 15442 27872
rect 16482 27860 16488 27872
rect 15436 27832 16488 27860
rect 15436 27820 15442 27832
rect 16482 27820 16488 27832
rect 16540 27820 16546 27872
rect 18616 27860 18644 27900
rect 18690 27888 18696 27940
rect 18748 27928 18754 27940
rect 23658 27928 23664 27940
rect 18748 27900 23664 27928
rect 18748 27888 18754 27900
rect 23658 27888 23664 27900
rect 23716 27888 23722 27940
rect 25240 27937 25268 27968
rect 25498 27956 25504 28008
rect 25556 27996 25562 28008
rect 25608 27996 25636 28027
rect 25774 28024 25780 28076
rect 25832 28024 25838 28076
rect 26602 28024 26608 28076
rect 26660 28064 26666 28076
rect 27632 28064 27660 28104
rect 26660 28036 27660 28064
rect 26660 28024 26666 28036
rect 27706 28024 27712 28076
rect 27764 28024 27770 28076
rect 27798 28024 27804 28076
rect 27856 28064 27862 28076
rect 27985 28067 28043 28073
rect 27856 28036 27901 28064
rect 27856 28024 27862 28036
rect 27985 28033 27997 28067
rect 28031 28033 28043 28067
rect 27985 28027 28043 28033
rect 28077 28067 28135 28073
rect 28077 28033 28089 28067
rect 28123 28033 28135 28067
rect 28077 28027 28135 28033
rect 25556 27968 25636 27996
rect 25556 27956 25562 27968
rect 23753 27931 23811 27937
rect 23753 27897 23765 27931
rect 23799 27928 23811 27931
rect 25225 27931 25283 27937
rect 23799 27900 25176 27928
rect 23799 27897 23811 27900
rect 23753 27891 23811 27897
rect 19518 27860 19524 27872
rect 18616 27832 19524 27860
rect 19518 27820 19524 27832
rect 19576 27820 19582 27872
rect 21726 27820 21732 27872
rect 21784 27860 21790 27872
rect 22002 27860 22008 27872
rect 21784 27832 22008 27860
rect 21784 27820 21790 27832
rect 22002 27820 22008 27832
rect 22060 27820 22066 27872
rect 24486 27820 24492 27872
rect 24544 27860 24550 27872
rect 24581 27863 24639 27869
rect 24581 27860 24593 27863
rect 24544 27832 24593 27860
rect 24544 27820 24550 27832
rect 24581 27829 24593 27832
rect 24627 27829 24639 27863
rect 24581 27823 24639 27829
rect 24946 27820 24952 27872
rect 25004 27860 25010 27872
rect 25041 27863 25099 27869
rect 25041 27860 25053 27863
rect 25004 27832 25053 27860
rect 25004 27820 25010 27832
rect 25041 27829 25053 27832
rect 25087 27829 25099 27863
rect 25148 27860 25176 27900
rect 25225 27897 25237 27931
rect 25271 27897 25283 27931
rect 25608 27928 25636 27968
rect 25682 27956 25688 28008
rect 25740 27996 25746 28008
rect 27724 27996 27752 28024
rect 25740 27968 27752 27996
rect 25740 27956 25746 27968
rect 27246 27928 27252 27940
rect 25608 27900 27252 27928
rect 25225 27891 25283 27897
rect 27246 27888 27252 27900
rect 27304 27928 27310 27940
rect 28000 27928 28028 28027
rect 27304 27900 28028 27928
rect 27304 27888 27310 27900
rect 26510 27860 26516 27872
rect 25148 27832 26516 27860
rect 25041 27823 25099 27829
rect 26510 27820 26516 27832
rect 26568 27820 26574 27872
rect 28092 27860 28120 28027
rect 28166 28024 28172 28076
rect 28224 28073 28230 28076
rect 28224 28064 28232 28073
rect 28224 28036 28396 28064
rect 28224 28027 28232 28036
rect 28224 28024 28230 28027
rect 28368 27996 28396 28036
rect 28442 28024 28448 28076
rect 28500 28024 28506 28076
rect 28552 28064 28580 28104
rect 28813 28067 28871 28073
rect 28813 28064 28825 28067
rect 28552 28036 28825 28064
rect 28813 28033 28825 28036
rect 28859 28033 28871 28067
rect 28813 28027 28871 28033
rect 28534 27996 28540 28008
rect 28368 27968 28540 27996
rect 28534 27956 28540 27968
rect 28592 27956 28598 28008
rect 29380 27996 29408 28104
rect 29546 28092 29552 28144
rect 29604 28132 29610 28144
rect 29604 28104 29868 28132
rect 29604 28092 29610 28104
rect 29454 28024 29460 28076
rect 29512 28064 29518 28076
rect 29733 28067 29791 28073
rect 29733 28064 29745 28067
rect 29512 28036 29745 28064
rect 29512 28024 29518 28036
rect 29733 28033 29745 28036
rect 29779 28033 29791 28067
rect 29840 28064 29868 28104
rect 29914 28092 29920 28144
rect 29972 28132 29978 28144
rect 31036 28132 31064 28172
rect 33134 28160 33140 28172
rect 33192 28160 33198 28212
rect 33870 28160 33876 28212
rect 33928 28200 33934 28212
rect 33928 28172 34468 28200
rect 33928 28160 33934 28172
rect 34440 28144 34468 28172
rect 37734 28160 37740 28212
rect 37792 28160 37798 28212
rect 37826 28160 37832 28212
rect 37884 28200 37890 28212
rect 38289 28203 38347 28209
rect 38289 28200 38301 28203
rect 37884 28172 38301 28200
rect 37884 28160 37890 28172
rect 38289 28169 38301 28172
rect 38335 28169 38347 28203
rect 38289 28163 38347 28169
rect 39022 28160 39028 28212
rect 39080 28200 39086 28212
rect 39669 28203 39727 28209
rect 39669 28200 39681 28203
rect 39080 28172 39681 28200
rect 39080 28160 39086 28172
rect 39669 28169 39681 28172
rect 39715 28169 39727 28203
rect 39669 28163 39727 28169
rect 39758 28160 39764 28212
rect 39816 28160 39822 28212
rect 29972 28104 30512 28132
rect 29972 28092 29978 28104
rect 30193 28067 30251 28073
rect 30193 28064 30205 28067
rect 29840 28036 30205 28064
rect 29733 28027 29791 28033
rect 30193 28033 30205 28036
rect 30239 28033 30251 28067
rect 30193 28027 30251 28033
rect 30374 28024 30380 28076
rect 30432 28024 30438 28076
rect 30484 28073 30512 28104
rect 30576 28104 31064 28132
rect 30576 28073 30604 28104
rect 31110 28092 31116 28144
rect 31168 28132 31174 28144
rect 31168 28104 32720 28132
rect 31168 28092 31174 28104
rect 30469 28067 30527 28073
rect 30469 28033 30481 28067
rect 30515 28033 30527 28067
rect 30469 28027 30527 28033
rect 30561 28067 30619 28073
rect 30561 28033 30573 28067
rect 30607 28033 30619 28067
rect 30561 28027 30619 28033
rect 29549 27999 29607 28005
rect 29549 27996 29561 27999
rect 29380 27968 29561 27996
rect 29549 27965 29561 27968
rect 29595 27996 29607 27999
rect 29638 27996 29644 28008
rect 29595 27968 29644 27996
rect 29595 27965 29607 27968
rect 29549 27959 29607 27965
rect 29638 27956 29644 27968
rect 29696 27956 29702 28008
rect 30006 27956 30012 28008
rect 30064 27996 30070 28008
rect 30576 27996 30604 28027
rect 30834 28024 30840 28076
rect 30892 28024 30898 28076
rect 31021 28067 31079 28073
rect 31021 28033 31033 28067
rect 31067 28064 31079 28067
rect 31202 28064 31208 28076
rect 31067 28036 31208 28064
rect 31067 28033 31079 28036
rect 31021 28027 31079 28033
rect 31202 28024 31208 28036
rect 31260 28024 31266 28076
rect 32306 28024 32312 28076
rect 32364 28024 32370 28076
rect 32692 28073 32720 28104
rect 32766 28092 32772 28144
rect 32824 28132 32830 28144
rect 34241 28135 34299 28141
rect 32824 28104 34099 28132
rect 32824 28092 32830 28104
rect 32401 28067 32459 28073
rect 32401 28033 32413 28067
rect 32447 28033 32459 28067
rect 32401 28027 32459 28033
rect 32677 28067 32735 28073
rect 32677 28033 32689 28067
rect 32723 28064 32735 28067
rect 33594 28064 33600 28076
rect 32723 28036 33600 28064
rect 32723 28033 32735 28036
rect 32677 28027 32735 28033
rect 30064 27968 30604 27996
rect 30852 27996 30880 28024
rect 31846 27996 31852 28008
rect 30852 27968 31852 27996
rect 30064 27956 30070 27968
rect 31846 27956 31852 27968
rect 31904 27956 31910 28008
rect 32416 27996 32444 28027
rect 33594 28024 33600 28036
rect 33652 28024 33658 28076
rect 33689 28067 33747 28073
rect 33689 28033 33701 28067
rect 33735 28064 33747 28067
rect 33870 28064 33876 28076
rect 33735 28036 33876 28064
rect 33735 28033 33747 28036
rect 33689 28027 33747 28033
rect 33870 28024 33876 28036
rect 33928 28024 33934 28076
rect 33965 28067 34023 28073
rect 33965 28033 33977 28067
rect 34011 28033 34023 28067
rect 34071 28064 34099 28104
rect 34241 28101 34253 28135
rect 34287 28132 34299 28135
rect 34330 28132 34336 28144
rect 34287 28104 34336 28132
rect 34287 28101 34299 28104
rect 34241 28095 34299 28101
rect 34330 28092 34336 28104
rect 34388 28092 34394 28144
rect 34422 28092 34428 28144
rect 34480 28092 34486 28144
rect 37366 28092 37372 28144
rect 37424 28132 37430 28144
rect 38565 28135 38623 28141
rect 37424 28104 37872 28132
rect 37424 28092 37430 28104
rect 37844 28073 37872 28104
rect 38565 28101 38577 28135
rect 38611 28132 38623 28135
rect 39390 28132 39396 28144
rect 38611 28104 39396 28132
rect 38611 28101 38623 28104
rect 38565 28095 38623 28101
rect 39390 28092 39396 28104
rect 39448 28092 39454 28144
rect 37829 28067 37887 28073
rect 34071 28036 37688 28064
rect 33965 28027 34023 28033
rect 33502 27996 33508 28008
rect 32416 27968 33508 27996
rect 33502 27956 33508 27968
rect 33560 27956 33566 28008
rect 33980 27996 34008 28027
rect 34698 27996 34704 28008
rect 33980 27968 34704 27996
rect 34698 27956 34704 27968
rect 34756 27956 34762 28008
rect 37550 27956 37556 28008
rect 37608 27956 37614 28008
rect 37660 27996 37688 28036
rect 37829 28033 37841 28067
rect 37875 28064 37887 28067
rect 38010 28064 38016 28076
rect 37875 28036 38016 28064
rect 37875 28033 37887 28036
rect 37829 28027 37887 28033
rect 38010 28024 38016 28036
rect 38068 28024 38074 28076
rect 38470 28024 38476 28076
rect 38528 28024 38534 28076
rect 38654 28024 38660 28076
rect 38712 28024 38718 28076
rect 38838 28024 38844 28076
rect 38896 28024 38902 28076
rect 39022 28024 39028 28076
rect 39080 28024 39086 28076
rect 40034 28024 40040 28076
rect 40092 28064 40098 28076
rect 40221 28067 40279 28073
rect 40221 28064 40233 28067
rect 40092 28036 40233 28064
rect 40092 28024 40098 28036
rect 40221 28033 40233 28036
rect 40267 28033 40279 28067
rect 40221 28027 40279 28033
rect 40405 28067 40463 28073
rect 40405 28033 40417 28067
rect 40451 28033 40463 28067
rect 40405 28027 40463 28033
rect 39485 27999 39543 28005
rect 39485 27996 39497 27999
rect 37660 27968 39497 27996
rect 39485 27965 39497 27968
rect 39531 27965 39543 27999
rect 39485 27959 39543 27965
rect 28353 27931 28411 27937
rect 28353 27897 28365 27931
rect 28399 27928 28411 27931
rect 28626 27928 28632 27940
rect 28399 27900 28632 27928
rect 28399 27897 28411 27900
rect 28353 27891 28411 27897
rect 28626 27888 28632 27900
rect 28684 27888 28690 27940
rect 29086 27928 29092 27940
rect 28920 27900 29092 27928
rect 28920 27860 28948 27900
rect 29086 27888 29092 27900
rect 29144 27928 29150 27940
rect 30190 27928 30196 27940
rect 29144 27900 30196 27928
rect 29144 27888 29150 27900
rect 30190 27888 30196 27900
rect 30248 27888 30254 27940
rect 30745 27931 30803 27937
rect 30745 27897 30757 27931
rect 30791 27928 30803 27931
rect 40420 27928 40448 28027
rect 41506 28024 41512 28076
rect 41564 28024 41570 28076
rect 41874 28024 41880 28076
rect 41932 28024 41938 28076
rect 30791 27900 40448 27928
rect 30791 27897 30803 27900
rect 30745 27891 30803 27897
rect 41690 27888 41696 27940
rect 41748 27888 41754 27940
rect 28092 27832 28948 27860
rect 30098 27820 30104 27872
rect 30156 27820 30162 27872
rect 32122 27820 32128 27872
rect 32180 27820 32186 27872
rect 32582 27820 32588 27872
rect 32640 27860 32646 27872
rect 33778 27860 33784 27872
rect 32640 27832 33784 27860
rect 32640 27820 32646 27832
rect 33778 27820 33784 27832
rect 33836 27820 33842 27872
rect 34149 27863 34207 27869
rect 34149 27829 34161 27863
rect 34195 27860 34207 27863
rect 34514 27860 34520 27872
rect 34195 27832 34520 27860
rect 34195 27829 34207 27832
rect 34149 27823 34207 27829
rect 34514 27820 34520 27832
rect 34572 27820 34578 27872
rect 34606 27820 34612 27872
rect 34664 27820 34670 27872
rect 35158 27820 35164 27872
rect 35216 27860 35222 27872
rect 35526 27860 35532 27872
rect 35216 27832 35532 27860
rect 35216 27820 35222 27832
rect 35526 27820 35532 27832
rect 35584 27820 35590 27872
rect 38194 27820 38200 27872
rect 38252 27820 38258 27872
rect 39117 27863 39175 27869
rect 39117 27829 39129 27863
rect 39163 27860 39175 27863
rect 39390 27860 39396 27872
rect 39163 27832 39396 27860
rect 39163 27829 39175 27832
rect 39117 27823 39175 27829
rect 39390 27820 39396 27832
rect 39448 27820 39454 27872
rect 40129 27863 40187 27869
rect 40129 27829 40141 27863
rect 40175 27860 40187 27863
rect 40402 27860 40408 27872
rect 40175 27832 40408 27860
rect 40175 27829 40187 27832
rect 40129 27823 40187 27829
rect 40402 27820 40408 27832
rect 40460 27820 40466 27872
rect 40586 27820 40592 27872
rect 40644 27820 40650 27872
rect 42058 27820 42064 27872
rect 42116 27820 42122 27872
rect 1104 27770 42504 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 42504 27770
rect 1104 27696 42504 27718
rect 4154 27616 4160 27668
rect 4212 27656 4218 27668
rect 4982 27656 4988 27668
rect 4212 27628 4988 27656
rect 4212 27616 4218 27628
rect 4982 27616 4988 27628
rect 5040 27616 5046 27668
rect 5718 27656 5724 27668
rect 5092 27628 5724 27656
rect 4614 27548 4620 27600
rect 4672 27548 4678 27600
rect 5092 27588 5120 27628
rect 5718 27616 5724 27628
rect 5776 27616 5782 27668
rect 10962 27616 10968 27668
rect 11020 27616 11026 27668
rect 14921 27659 14979 27665
rect 14921 27625 14933 27659
rect 14967 27625 14979 27659
rect 14921 27619 14979 27625
rect 17129 27659 17187 27665
rect 17129 27625 17141 27659
rect 17175 27656 17187 27659
rect 18230 27656 18236 27668
rect 17175 27628 18236 27656
rect 17175 27625 17187 27628
rect 17129 27619 17187 27625
rect 4908 27560 5120 27588
rect 7653 27591 7711 27597
rect 3602 27412 3608 27464
rect 3660 27452 3666 27464
rect 4908 27461 4936 27560
rect 7653 27557 7665 27591
rect 7699 27588 7711 27591
rect 8294 27588 8300 27600
rect 7699 27560 8300 27588
rect 7699 27557 7711 27560
rect 7653 27551 7711 27557
rect 8294 27548 8300 27560
rect 8352 27548 8358 27600
rect 8389 27591 8447 27597
rect 8389 27557 8401 27591
rect 8435 27588 8447 27591
rect 9674 27588 9680 27600
rect 8435 27560 9680 27588
rect 8435 27557 8447 27560
rect 8389 27551 8447 27557
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 4985 27523 5043 27529
rect 4985 27489 4997 27523
rect 5031 27520 5043 27523
rect 6638 27520 6644 27532
rect 5031 27492 6644 27520
rect 5031 27489 5043 27492
rect 4985 27483 5043 27489
rect 6638 27480 6644 27492
rect 6696 27480 6702 27532
rect 7745 27523 7803 27529
rect 7745 27520 7757 27523
rect 7392 27492 7757 27520
rect 4617 27455 4675 27461
rect 4617 27452 4629 27455
rect 3660 27424 4629 27452
rect 3660 27412 3666 27424
rect 4617 27421 4629 27424
rect 4663 27421 4675 27455
rect 4617 27415 4675 27421
rect 4893 27455 4951 27461
rect 4893 27421 4905 27455
rect 4939 27421 4951 27455
rect 4893 27415 4951 27421
rect 2774 27344 2780 27396
rect 2832 27384 2838 27396
rect 4522 27384 4528 27396
rect 2832 27356 4528 27384
rect 2832 27344 2838 27356
rect 4522 27344 4528 27356
rect 4580 27344 4586 27396
rect 4632 27384 4660 27415
rect 7098 27412 7104 27464
rect 7156 27412 7162 27464
rect 7392 27461 7420 27492
rect 7745 27489 7757 27492
rect 7791 27520 7803 27523
rect 8018 27520 8024 27532
rect 7791 27492 8024 27520
rect 7791 27489 7803 27492
rect 7745 27483 7803 27489
rect 8018 27480 8024 27492
rect 8076 27480 8082 27532
rect 8128 27492 8432 27520
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27421 7435 27455
rect 7377 27415 7435 27421
rect 7466 27412 7472 27464
rect 7524 27412 7530 27464
rect 7903 27455 7961 27461
rect 7903 27421 7915 27455
rect 7949 27452 7961 27455
rect 8128 27452 8156 27492
rect 7949 27424 8156 27452
rect 8205 27455 8263 27461
rect 7949 27421 7961 27424
rect 7903 27415 7961 27421
rect 8205 27421 8217 27455
rect 8251 27421 8263 27455
rect 8404 27452 8432 27492
rect 9030 27480 9036 27532
rect 9088 27480 9094 27532
rect 10870 27480 10876 27532
rect 10928 27480 10934 27532
rect 10980 27520 11008 27616
rect 12897 27591 12955 27597
rect 12897 27588 12909 27591
rect 12406 27560 12909 27588
rect 12406 27520 12434 27560
rect 12897 27557 12909 27560
rect 12943 27557 12955 27591
rect 12897 27551 12955 27557
rect 14458 27548 14464 27600
rect 14516 27548 14522 27600
rect 14936 27588 14964 27619
rect 18230 27616 18236 27628
rect 18288 27616 18294 27668
rect 18874 27656 18880 27668
rect 18340 27628 18880 27656
rect 15194 27588 15200 27600
rect 14936 27560 15200 27588
rect 15194 27548 15200 27560
rect 15252 27548 15258 27600
rect 15286 27548 15292 27600
rect 15344 27548 15350 27600
rect 16850 27548 16856 27600
rect 16908 27588 16914 27600
rect 17773 27591 17831 27597
rect 16908 27560 16988 27588
rect 16908 27548 16914 27560
rect 10980 27492 12434 27520
rect 8404 27424 9352 27452
rect 8205 27415 8263 27421
rect 5166 27384 5172 27396
rect 4632 27356 5172 27384
rect 5166 27344 5172 27356
rect 5224 27344 5230 27396
rect 5261 27387 5319 27393
rect 5261 27353 5273 27387
rect 5307 27384 5319 27387
rect 5350 27384 5356 27396
rect 5307 27356 5356 27384
rect 5307 27353 5319 27356
rect 5261 27347 5319 27353
rect 5350 27344 5356 27356
rect 5408 27344 5414 27396
rect 5718 27344 5724 27396
rect 5776 27344 5782 27396
rect 7285 27387 7343 27393
rect 7285 27353 7297 27387
rect 7331 27384 7343 27387
rect 8021 27387 8079 27393
rect 8021 27384 8033 27387
rect 7331 27356 8033 27384
rect 7331 27353 7343 27356
rect 7285 27347 7343 27353
rect 7944 27328 7972 27356
rect 8021 27353 8033 27356
rect 8067 27353 8079 27387
rect 8021 27347 8079 27353
rect 8110 27344 8116 27396
rect 8168 27344 8174 27396
rect 4798 27276 4804 27328
rect 4856 27316 4862 27328
rect 6733 27319 6791 27325
rect 6733 27316 6745 27319
rect 4856 27288 6745 27316
rect 4856 27276 4862 27288
rect 6733 27285 6745 27288
rect 6779 27316 6791 27319
rect 6914 27316 6920 27328
rect 6779 27288 6920 27316
rect 6779 27285 6791 27288
rect 6733 27279 6791 27285
rect 6914 27276 6920 27288
rect 6972 27276 6978 27328
rect 7926 27276 7932 27328
rect 7984 27276 7990 27328
rect 8220 27316 8248 27415
rect 9324 27384 9352 27424
rect 9398 27412 9404 27464
rect 9456 27452 9462 27464
rect 9769 27455 9827 27461
rect 9769 27452 9781 27455
rect 9456 27424 9781 27452
rect 9456 27412 9462 27424
rect 9769 27421 9781 27424
rect 9815 27421 9827 27455
rect 12406 27452 12434 27492
rect 13906 27480 13912 27532
rect 13964 27520 13970 27532
rect 14918 27520 14924 27532
rect 13964 27492 14924 27520
rect 13964 27480 13970 27492
rect 14918 27480 14924 27492
rect 14976 27520 14982 27532
rect 15381 27523 15439 27529
rect 15381 27520 15393 27523
rect 14976 27492 15393 27520
rect 14976 27480 14982 27492
rect 15381 27489 15393 27492
rect 15427 27489 15439 27523
rect 15381 27483 15439 27489
rect 12282 27424 12434 27452
rect 9769 27415 9827 27421
rect 12710 27412 12716 27464
rect 12768 27412 12774 27464
rect 14642 27412 14648 27464
rect 14700 27412 14706 27464
rect 14737 27455 14795 27461
rect 14737 27421 14749 27455
rect 14783 27421 14795 27455
rect 14737 27415 14795 27421
rect 9677 27387 9735 27393
rect 9677 27384 9689 27387
rect 9324 27356 9689 27384
rect 9677 27353 9689 27356
rect 9723 27384 9735 27387
rect 11054 27384 11060 27396
rect 9723 27356 11060 27384
rect 9723 27353 9735 27356
rect 9677 27347 9735 27353
rect 11054 27344 11060 27356
rect 11112 27344 11118 27396
rect 11146 27344 11152 27396
rect 11204 27344 11210 27396
rect 13354 27344 13360 27396
rect 13412 27384 13418 27396
rect 14752 27384 14780 27415
rect 15010 27412 15016 27464
rect 15068 27412 15074 27464
rect 16960 27452 16988 27560
rect 17773 27557 17785 27591
rect 17819 27588 17831 27591
rect 17862 27588 17868 27600
rect 17819 27560 17868 27588
rect 17819 27557 17831 27560
rect 17773 27551 17831 27557
rect 17862 27548 17868 27560
rect 17920 27548 17926 27600
rect 18340 27588 18368 27628
rect 18874 27616 18880 27628
rect 18932 27616 18938 27668
rect 19426 27616 19432 27668
rect 19484 27656 19490 27668
rect 19521 27659 19579 27665
rect 19521 27656 19533 27659
rect 19484 27628 19533 27656
rect 19484 27616 19490 27628
rect 19521 27625 19533 27628
rect 19567 27625 19579 27659
rect 19521 27619 19579 27625
rect 21729 27659 21787 27665
rect 21729 27625 21741 27659
rect 21775 27656 21787 27659
rect 22370 27656 22376 27668
rect 21775 27628 22376 27656
rect 21775 27625 21787 27628
rect 21729 27619 21787 27625
rect 22370 27616 22376 27628
rect 22428 27656 22434 27668
rect 23106 27656 23112 27668
rect 22428 27628 23112 27656
rect 22428 27616 22434 27628
rect 23106 27616 23112 27628
rect 23164 27616 23170 27668
rect 24486 27616 24492 27668
rect 24544 27656 24550 27668
rect 24654 27659 24712 27665
rect 24654 27656 24666 27659
rect 24544 27628 24666 27656
rect 24544 27616 24550 27628
rect 24654 27625 24666 27628
rect 24700 27625 24712 27659
rect 24654 27619 24712 27625
rect 25222 27616 25228 27668
rect 25280 27656 25286 27668
rect 26145 27659 26203 27665
rect 26145 27656 26157 27659
rect 25280 27628 26157 27656
rect 25280 27616 25286 27628
rect 26145 27625 26157 27628
rect 26191 27625 26203 27659
rect 27246 27656 27252 27668
rect 26145 27619 26203 27625
rect 26344 27628 27252 27656
rect 18008 27560 18368 27588
rect 18008 27520 18036 27560
rect 18414 27548 18420 27600
rect 18472 27588 18478 27600
rect 19889 27591 19947 27597
rect 19889 27588 19901 27591
rect 18472 27560 19901 27588
rect 18472 27548 18478 27560
rect 19889 27557 19901 27560
rect 19935 27557 19947 27591
rect 19889 27551 19947 27557
rect 19981 27591 20039 27597
rect 19981 27557 19993 27591
rect 20027 27588 20039 27591
rect 20070 27588 20076 27600
rect 20027 27560 20076 27588
rect 20027 27557 20039 27560
rect 19981 27551 20039 27557
rect 18008 27492 18092 27520
rect 17497 27455 17555 27461
rect 17497 27452 17509 27455
rect 16960 27424 17509 27452
rect 17497 27421 17509 27424
rect 17543 27421 17555 27455
rect 17954 27452 17960 27464
rect 17497 27415 17555 27421
rect 17604 27424 17960 27452
rect 14826 27384 14832 27396
rect 13412 27356 14832 27384
rect 13412 27344 13418 27356
rect 14826 27344 14832 27356
rect 14884 27344 14890 27396
rect 14918 27344 14924 27396
rect 14976 27344 14982 27396
rect 15289 27387 15347 27393
rect 15289 27353 15301 27387
rect 15335 27384 15347 27387
rect 15562 27384 15568 27396
rect 15335 27356 15568 27384
rect 15335 27353 15347 27356
rect 15289 27347 15347 27353
rect 15562 27344 15568 27356
rect 15620 27344 15626 27396
rect 15654 27344 15660 27396
rect 15712 27344 15718 27396
rect 16882 27356 16988 27384
rect 9306 27316 9312 27328
rect 8220 27288 9312 27316
rect 9306 27276 9312 27288
rect 9364 27276 9370 27328
rect 10134 27276 10140 27328
rect 10192 27316 10198 27328
rect 10413 27319 10471 27325
rect 10413 27316 10425 27319
rect 10192 27288 10425 27316
rect 10192 27276 10198 27288
rect 10413 27285 10425 27288
rect 10459 27285 10471 27319
rect 10413 27279 10471 27285
rect 11974 27276 11980 27328
rect 12032 27316 12038 27328
rect 12621 27319 12679 27325
rect 12621 27316 12633 27319
rect 12032 27288 12633 27316
rect 12032 27276 12038 27288
rect 12621 27285 12633 27288
rect 12667 27316 12679 27319
rect 14366 27316 14372 27328
rect 12667 27288 14372 27316
rect 12667 27285 12679 27288
rect 12621 27279 12679 27285
rect 14366 27276 14372 27288
rect 14424 27276 14430 27328
rect 14458 27276 14464 27328
rect 14516 27316 14522 27328
rect 15102 27316 15108 27328
rect 14516 27288 15108 27316
rect 14516 27276 14522 27288
rect 15102 27276 15108 27288
rect 15160 27276 15166 27328
rect 16960 27316 16988 27356
rect 17034 27344 17040 27396
rect 17092 27384 17098 27396
rect 17313 27387 17371 27393
rect 17313 27384 17325 27387
rect 17092 27356 17325 27384
rect 17092 27344 17098 27356
rect 17313 27353 17325 27356
rect 17359 27353 17371 27387
rect 17313 27347 17371 27353
rect 17126 27316 17132 27328
rect 16960 27288 17132 27316
rect 17126 27276 17132 27288
rect 17184 27276 17190 27328
rect 17402 27276 17408 27328
rect 17460 27316 17466 27328
rect 17604 27316 17632 27424
rect 17954 27412 17960 27424
rect 18012 27412 18018 27464
rect 18064 27461 18092 27492
rect 18230 27480 18236 27532
rect 18288 27520 18294 27532
rect 18288 27492 18644 27520
rect 18288 27480 18294 27492
rect 18616 27461 18644 27492
rect 19150 27480 19156 27532
rect 19208 27520 19214 27532
rect 19797 27523 19855 27529
rect 19797 27520 19809 27523
rect 19208 27492 19809 27520
rect 19208 27480 19214 27492
rect 19797 27489 19809 27492
rect 19843 27489 19855 27523
rect 19904 27520 19932 27551
rect 20070 27548 20076 27560
rect 20128 27548 20134 27600
rect 22002 27548 22008 27600
rect 22060 27548 22066 27600
rect 26344 27597 26372 27628
rect 27246 27616 27252 27628
rect 27304 27616 27310 27668
rect 27614 27616 27620 27668
rect 27672 27656 27678 27668
rect 30834 27656 30840 27668
rect 27672 27628 30840 27656
rect 27672 27616 27678 27628
rect 30834 27616 30840 27628
rect 30892 27616 30898 27668
rect 31928 27659 31986 27665
rect 31928 27625 31940 27659
rect 31974 27656 31986 27659
rect 32122 27656 32128 27668
rect 31974 27628 32128 27656
rect 31974 27625 31986 27628
rect 31928 27619 31986 27625
rect 32122 27616 32128 27628
rect 32180 27616 32186 27668
rect 33594 27656 33600 27668
rect 33428 27628 33600 27656
rect 26329 27591 26387 27597
rect 26329 27557 26341 27591
rect 26375 27557 26387 27591
rect 26329 27551 26387 27557
rect 26789 27591 26847 27597
rect 26789 27557 26801 27591
rect 26835 27588 26847 27591
rect 27154 27588 27160 27600
rect 26835 27560 27160 27588
rect 26835 27557 26847 27560
rect 26789 27551 26847 27557
rect 27154 27548 27160 27560
rect 27212 27548 27218 27600
rect 29178 27588 29184 27600
rect 28552 27560 29184 27588
rect 19904 27492 20668 27520
rect 19797 27483 19855 27489
rect 18049 27455 18107 27461
rect 18049 27421 18061 27455
rect 18095 27421 18107 27455
rect 18049 27415 18107 27421
rect 18141 27455 18199 27461
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 18325 27455 18383 27461
rect 18187 27424 18276 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 17681 27387 17739 27393
rect 17681 27353 17693 27387
rect 17727 27353 17739 27387
rect 17681 27347 17739 27353
rect 17460 27288 17632 27316
rect 17696 27316 17724 27347
rect 17770 27344 17776 27396
rect 17828 27344 17834 27396
rect 17954 27316 17960 27328
rect 17696 27288 17960 27316
rect 17460 27276 17466 27288
rect 17954 27276 17960 27288
rect 18012 27276 18018 27328
rect 18138 27276 18144 27328
rect 18196 27276 18202 27328
rect 18248 27316 18276 27424
rect 18325 27421 18337 27455
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18417 27455 18475 27461
rect 18417 27421 18429 27455
rect 18463 27452 18475 27455
rect 18601 27455 18659 27461
rect 18463 27424 18552 27452
rect 18463 27421 18475 27424
rect 18417 27415 18475 27421
rect 18340 27384 18368 27415
rect 18524 27384 18552 27424
rect 18601 27421 18613 27455
rect 18647 27452 18659 27455
rect 20349 27455 20407 27461
rect 20349 27452 20361 27455
rect 18647 27424 20361 27452
rect 18647 27421 18659 27424
rect 18601 27415 18659 27421
rect 20349 27421 20361 27424
rect 20395 27421 20407 27455
rect 20349 27415 20407 27421
rect 20530 27412 20536 27464
rect 20588 27412 20594 27464
rect 20640 27461 20668 27492
rect 21634 27480 21640 27532
rect 21692 27520 21698 27532
rect 23014 27520 23020 27532
rect 21692 27492 21772 27520
rect 21692 27480 21698 27492
rect 21744 27461 21772 27492
rect 22480 27492 23020 27520
rect 20625 27455 20683 27461
rect 20625 27421 20637 27455
rect 20671 27421 20683 27455
rect 20625 27415 20683 27421
rect 21545 27455 21603 27461
rect 21545 27421 21557 27455
rect 21591 27421 21603 27455
rect 21545 27415 21603 27421
rect 21729 27455 21787 27461
rect 21729 27421 21741 27455
rect 21775 27421 21787 27455
rect 21729 27415 21787 27421
rect 20070 27384 20076 27396
rect 18340 27356 18460 27384
rect 18524 27356 20076 27384
rect 18322 27316 18328 27328
rect 18248 27288 18328 27316
rect 18322 27276 18328 27288
rect 18380 27276 18386 27328
rect 18432 27316 18460 27356
rect 18616 27328 18644 27356
rect 20070 27344 20076 27356
rect 20128 27344 20134 27396
rect 20438 27344 20444 27396
rect 20496 27384 20502 27396
rect 21560 27384 21588 27415
rect 21818 27412 21824 27464
rect 21876 27412 21882 27464
rect 22005 27455 22063 27461
rect 22005 27421 22017 27455
rect 22051 27452 22063 27455
rect 22094 27452 22100 27464
rect 22051 27424 22100 27452
rect 22051 27421 22063 27424
rect 22005 27415 22063 27421
rect 22094 27412 22100 27424
rect 22152 27452 22158 27464
rect 22480 27461 22508 27492
rect 23014 27480 23020 27492
rect 23072 27480 23078 27532
rect 23842 27480 23848 27532
rect 23900 27520 23906 27532
rect 24394 27520 24400 27532
rect 23900 27492 24400 27520
rect 23900 27480 23906 27492
rect 24044 27461 24072 27492
rect 24394 27480 24400 27492
rect 24452 27520 24458 27532
rect 24670 27520 24676 27532
rect 24452 27492 24676 27520
rect 24452 27480 24458 27492
rect 24670 27480 24676 27492
rect 24728 27480 24734 27532
rect 27522 27520 27528 27532
rect 26620 27492 27528 27520
rect 22465 27455 22523 27461
rect 22152 27424 22197 27452
rect 22152 27412 22158 27424
rect 22465 27421 22477 27455
rect 22511 27421 22523 27455
rect 22465 27415 22523 27421
rect 24029 27455 24087 27461
rect 24029 27421 24041 27455
rect 24075 27421 24087 27455
rect 24029 27415 24087 27421
rect 26510 27412 26516 27464
rect 26568 27446 26574 27464
rect 26620 27446 26648 27492
rect 27522 27480 27528 27492
rect 27580 27480 27586 27532
rect 28552 27529 28580 27560
rect 29178 27548 29184 27560
rect 29236 27588 29242 27600
rect 29236 27560 29960 27588
rect 29236 27548 29242 27560
rect 29932 27532 29960 27560
rect 30650 27548 30656 27600
rect 30708 27588 30714 27600
rect 33428 27597 33456 27628
rect 33594 27616 33600 27628
rect 33652 27656 33658 27668
rect 33652 27628 33732 27656
rect 33652 27616 33658 27628
rect 33413 27591 33471 27597
rect 30708 27560 31800 27588
rect 30708 27548 30714 27560
rect 28537 27523 28595 27529
rect 28537 27489 28549 27523
rect 28583 27489 28595 27523
rect 28537 27483 28595 27489
rect 28626 27480 28632 27532
rect 28684 27520 28690 27532
rect 29089 27523 29147 27529
rect 28684 27492 28948 27520
rect 28684 27480 28690 27492
rect 26568 27418 26648 27446
rect 26568 27412 26574 27418
rect 28810 27412 28816 27464
rect 28868 27412 28874 27464
rect 28920 27461 28948 27492
rect 29089 27489 29101 27523
rect 29135 27520 29147 27523
rect 29270 27520 29276 27532
rect 29135 27492 29276 27520
rect 29135 27489 29147 27492
rect 29089 27483 29147 27489
rect 29270 27480 29276 27492
rect 29328 27480 29334 27532
rect 29914 27480 29920 27532
rect 29972 27520 29978 27532
rect 31662 27520 31668 27532
rect 29972 27492 31668 27520
rect 29972 27480 29978 27492
rect 31662 27480 31668 27492
rect 31720 27480 31726 27532
rect 31772 27520 31800 27560
rect 33413 27557 33425 27591
rect 33459 27557 33471 27591
rect 33413 27551 33471 27557
rect 33502 27548 33508 27600
rect 33560 27548 33566 27600
rect 33704 27588 33732 27628
rect 33778 27616 33784 27668
rect 33836 27656 33842 27668
rect 35526 27656 35532 27668
rect 33836 27628 35532 27656
rect 33836 27616 33842 27628
rect 35526 27616 35532 27628
rect 35584 27616 35590 27668
rect 35986 27616 35992 27668
rect 36044 27656 36050 27668
rect 37734 27656 37740 27668
rect 36044 27628 37740 27656
rect 36044 27616 36050 27628
rect 37734 27616 37740 27628
rect 37792 27616 37798 27668
rect 40392 27659 40450 27665
rect 40392 27625 40404 27659
rect 40438 27656 40450 27659
rect 40586 27656 40592 27668
rect 40438 27628 40592 27656
rect 40438 27625 40450 27628
rect 40392 27619 40450 27625
rect 40586 27616 40592 27628
rect 40644 27616 40650 27668
rect 41874 27616 41880 27668
rect 41932 27616 41938 27668
rect 33870 27588 33876 27600
rect 33704 27560 33876 27588
rect 33870 27548 33876 27560
rect 33928 27548 33934 27600
rect 33962 27548 33968 27600
rect 34020 27548 34026 27600
rect 34146 27548 34152 27600
rect 34204 27588 34210 27600
rect 34204 27560 35112 27588
rect 34204 27548 34210 27560
rect 33980 27520 34008 27548
rect 34330 27520 34336 27532
rect 31772 27492 33916 27520
rect 33980 27492 34192 27520
rect 28905 27455 28963 27461
rect 28905 27421 28917 27455
rect 28951 27421 28963 27455
rect 28905 27415 28963 27421
rect 29178 27412 29184 27464
rect 29236 27412 29242 27464
rect 30650 27412 30656 27464
rect 30708 27412 30714 27464
rect 30745 27455 30803 27461
rect 30745 27421 30757 27455
rect 30791 27452 30803 27455
rect 30834 27452 30840 27464
rect 30791 27424 30840 27452
rect 30791 27421 30803 27424
rect 30745 27415 30803 27421
rect 30834 27412 30840 27424
rect 30892 27412 30898 27464
rect 30926 27412 30932 27464
rect 30984 27412 30990 27464
rect 31031 27433 31089 27439
rect 31031 27399 31043 27433
rect 31077 27399 31089 27433
rect 33042 27412 33048 27464
rect 33100 27412 33106 27464
rect 33226 27412 33232 27464
rect 33284 27452 33290 27464
rect 33643 27455 33701 27461
rect 33643 27452 33655 27455
rect 33284 27424 33655 27452
rect 33284 27412 33290 27424
rect 33643 27421 33655 27424
rect 33689 27421 33701 27455
rect 33643 27415 33701 27421
rect 33778 27412 33784 27464
rect 33836 27412 33842 27464
rect 33888 27461 33916 27492
rect 34164 27461 34192 27492
rect 34256 27492 34336 27520
rect 34256 27461 34284 27492
rect 34330 27480 34336 27492
rect 34388 27480 34394 27532
rect 34606 27480 34612 27532
rect 34664 27520 34670 27532
rect 35084 27529 35112 27560
rect 35342 27548 35348 27600
rect 35400 27588 35406 27600
rect 35400 27560 35756 27588
rect 35400 27548 35406 27560
rect 34885 27523 34943 27529
rect 34885 27520 34897 27523
rect 34664 27492 34897 27520
rect 34664 27480 34670 27492
rect 34885 27489 34897 27492
rect 34931 27489 34943 27523
rect 34885 27483 34943 27489
rect 35069 27523 35127 27529
rect 35069 27489 35081 27523
rect 35115 27489 35127 27523
rect 35069 27483 35127 27489
rect 35437 27523 35495 27529
rect 35437 27489 35449 27523
rect 35483 27520 35495 27523
rect 35526 27520 35532 27532
rect 35483 27492 35532 27520
rect 35483 27489 35495 27492
rect 35437 27483 35495 27489
rect 35526 27480 35532 27492
rect 35584 27480 35590 27532
rect 33873 27455 33931 27461
rect 33873 27421 33885 27455
rect 33919 27421 33931 27455
rect 34001 27455 34059 27461
rect 34001 27452 34013 27455
rect 33873 27415 33931 27421
rect 33980 27421 34013 27452
rect 34047 27421 34059 27455
rect 33980 27415 34059 27421
rect 34149 27455 34207 27461
rect 34149 27421 34161 27455
rect 34195 27421 34207 27455
rect 34149 27415 34207 27421
rect 34241 27455 34299 27461
rect 34241 27421 34253 27455
rect 34287 27421 34299 27455
rect 34241 27415 34299 27421
rect 31031 27396 31089 27399
rect 20496 27356 21588 27384
rect 20496 27344 20502 27356
rect 22554 27344 22560 27396
rect 22612 27384 22618 27396
rect 22649 27387 22707 27393
rect 22649 27384 22661 27387
rect 22612 27356 22661 27384
rect 22612 27344 22618 27356
rect 22649 27353 22661 27356
rect 22695 27353 22707 27387
rect 22649 27347 22707 27353
rect 22830 27344 22836 27396
rect 22888 27344 22894 27396
rect 26234 27384 26240 27396
rect 25898 27356 26240 27384
rect 26234 27344 26240 27356
rect 26292 27384 26298 27396
rect 28261 27387 28319 27393
rect 26292 27356 27094 27384
rect 26292 27344 26298 27356
rect 28261 27353 28273 27387
rect 28307 27384 28319 27387
rect 28629 27387 28687 27393
rect 28629 27384 28641 27387
rect 28307 27356 28641 27384
rect 28307 27353 28319 27356
rect 28261 27347 28319 27353
rect 28629 27353 28641 27356
rect 28675 27353 28687 27387
rect 31018 27384 31024 27396
rect 28629 27347 28687 27353
rect 28966 27356 31024 27384
rect 18506 27316 18512 27328
rect 18432 27288 18512 27316
rect 18506 27276 18512 27288
rect 18564 27276 18570 27328
rect 18598 27276 18604 27328
rect 18656 27276 18662 27328
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 22848 27316 22876 27344
rect 19116 27288 22876 27316
rect 19116 27276 19122 27288
rect 23014 27276 23020 27328
rect 23072 27316 23078 27328
rect 28966 27316 28994 27356
rect 31018 27344 31024 27356
rect 31076 27393 31089 27396
rect 31076 27344 31082 27393
rect 31478 27344 31484 27396
rect 31536 27344 31542 27396
rect 33888 27328 33916 27415
rect 23072 27288 28994 27316
rect 23072 27276 23078 27288
rect 30374 27276 30380 27328
rect 30432 27316 30438 27328
rect 30469 27319 30527 27325
rect 30469 27316 30481 27319
rect 30432 27288 30481 27316
rect 30432 27276 30438 27288
rect 30469 27285 30481 27288
rect 30515 27285 30527 27319
rect 30469 27279 30527 27285
rect 31202 27276 31208 27328
rect 31260 27276 31266 27328
rect 33870 27276 33876 27328
rect 33928 27276 33934 27328
rect 33980 27316 34008 27415
rect 34422 27412 34428 27464
rect 34480 27412 34486 27464
rect 34977 27455 35035 27461
rect 34977 27421 34989 27455
rect 35023 27421 35035 27455
rect 34977 27415 35035 27421
rect 35161 27455 35219 27461
rect 35161 27421 35173 27455
rect 35207 27452 35219 27455
rect 35250 27452 35256 27464
rect 35207 27424 35256 27452
rect 35207 27421 35219 27424
rect 35161 27415 35219 27421
rect 34333 27387 34391 27393
rect 34333 27353 34345 27387
rect 34379 27384 34391 27387
rect 34992 27384 35020 27415
rect 35250 27412 35256 27424
rect 35308 27412 35314 27464
rect 35728 27461 35756 27560
rect 37274 27548 37280 27600
rect 37332 27588 37338 27600
rect 38378 27588 38384 27600
rect 37332 27560 38384 27588
rect 37332 27548 37338 27560
rect 38378 27548 38384 27560
rect 38436 27548 38442 27600
rect 39117 27591 39175 27597
rect 39117 27557 39129 27591
rect 39163 27588 39175 27591
rect 40034 27588 40040 27600
rect 39163 27560 40040 27588
rect 39163 27557 39175 27560
rect 39117 27551 39175 27557
rect 40034 27548 40040 27560
rect 40092 27548 40098 27600
rect 38654 27480 38660 27532
rect 38712 27520 38718 27532
rect 41892 27520 41920 27616
rect 38712 27492 39528 27520
rect 38712 27480 38718 27492
rect 35345 27455 35403 27461
rect 35345 27421 35357 27455
rect 35391 27421 35403 27455
rect 35345 27415 35403 27421
rect 35621 27455 35679 27461
rect 35621 27421 35633 27455
rect 35667 27421 35679 27455
rect 35621 27415 35679 27421
rect 35713 27455 35771 27461
rect 35713 27421 35725 27455
rect 35759 27421 35771 27455
rect 35713 27415 35771 27421
rect 34379 27356 35020 27384
rect 35360 27384 35388 27415
rect 35526 27384 35532 27396
rect 35360 27356 35532 27384
rect 34379 27353 34391 27356
rect 34333 27347 34391 27353
rect 35526 27344 35532 27356
rect 35584 27344 35590 27396
rect 34054 27316 34060 27328
rect 33980 27288 34060 27316
rect 34054 27276 34060 27288
rect 34112 27276 34118 27328
rect 34698 27276 34704 27328
rect 34756 27276 34762 27328
rect 35636 27316 35664 27415
rect 35986 27412 35992 27464
rect 36044 27412 36050 27464
rect 39298 27412 39304 27464
rect 39356 27412 39362 27464
rect 39500 27396 39528 27492
rect 39684 27492 41920 27520
rect 39684 27461 39712 27492
rect 39669 27455 39727 27461
rect 39669 27421 39681 27455
rect 39715 27421 39727 27455
rect 39669 27415 39727 27421
rect 40126 27412 40132 27464
rect 40184 27412 40190 27464
rect 35897 27387 35955 27393
rect 35897 27353 35909 27387
rect 35943 27384 35955 27387
rect 36265 27387 36323 27393
rect 36265 27384 36277 27387
rect 35943 27356 36277 27384
rect 35943 27353 35955 27356
rect 35897 27347 35955 27353
rect 36265 27353 36277 27356
rect 36311 27353 36323 27387
rect 39022 27384 39028 27396
rect 37490 27356 39028 27384
rect 36265 27347 36323 27353
rect 39022 27344 39028 27356
rect 39080 27344 39086 27396
rect 39390 27344 39396 27396
rect 39448 27344 39454 27396
rect 39482 27344 39488 27396
rect 39540 27384 39546 27396
rect 39850 27384 39856 27396
rect 39540 27356 39856 27384
rect 39540 27344 39546 27356
rect 39850 27344 39856 27356
rect 39908 27344 39914 27396
rect 39942 27344 39948 27396
rect 40000 27384 40006 27396
rect 40000 27356 40894 27384
rect 40000 27344 40006 27356
rect 36630 27316 36636 27328
rect 35636 27288 36636 27316
rect 36630 27276 36636 27288
rect 36688 27276 36694 27328
rect 1104 27226 42504 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 42504 27226
rect 1104 27152 42504 27174
rect 4614 27072 4620 27124
rect 4672 27072 4678 27124
rect 4890 27072 4896 27124
rect 4948 27112 4954 27124
rect 4948 27084 5304 27112
rect 4948 27072 4954 27084
rect 4632 27044 4660 27072
rect 5276 27053 5304 27084
rect 5442 27072 5448 27124
rect 5500 27072 5506 27124
rect 5718 27072 5724 27124
rect 5776 27112 5782 27124
rect 6457 27115 6515 27121
rect 6457 27112 6469 27115
rect 5776 27084 6469 27112
rect 5776 27072 5782 27084
rect 6457 27081 6469 27084
rect 6503 27081 6515 27115
rect 6457 27075 6515 27081
rect 6748 27084 9260 27112
rect 6748 27053 6776 27084
rect 5077 27047 5135 27053
rect 5077 27044 5089 27047
rect 4356 27016 5089 27044
rect 4154 26936 4160 26988
rect 4212 26936 4218 26988
rect 4356 26985 4384 27016
rect 5077 27013 5089 27016
rect 5123 27013 5135 27047
rect 5077 27007 5135 27013
rect 5261 27047 5319 27053
rect 5261 27013 5273 27047
rect 5307 27013 5319 27047
rect 5261 27007 5319 27013
rect 6733 27047 6791 27053
rect 6733 27013 6745 27047
rect 6779 27013 6791 27047
rect 6733 27007 6791 27013
rect 9030 27004 9036 27056
rect 9088 27044 9094 27056
rect 9125 27047 9183 27053
rect 9125 27044 9137 27047
rect 9088 27016 9137 27044
rect 9088 27004 9094 27016
rect 9125 27013 9137 27016
rect 9171 27013 9183 27047
rect 9232 27044 9260 27084
rect 9306 27072 9312 27124
rect 9364 27072 9370 27124
rect 11146 27072 11152 27124
rect 11204 27112 11210 27124
rect 11517 27115 11575 27121
rect 11517 27112 11529 27115
rect 11204 27084 11529 27112
rect 11204 27072 11210 27084
rect 11517 27081 11529 27084
rect 11563 27081 11575 27115
rect 11517 27075 11575 27081
rect 11974 27072 11980 27124
rect 12032 27072 12038 27124
rect 15010 27072 15016 27124
rect 15068 27072 15074 27124
rect 15473 27115 15531 27121
rect 15473 27081 15485 27115
rect 15519 27112 15531 27115
rect 15654 27112 15660 27124
rect 15519 27084 15660 27112
rect 15519 27081 15531 27084
rect 15473 27075 15531 27081
rect 15654 27072 15660 27084
rect 15712 27072 15718 27124
rect 16298 27072 16304 27124
rect 16356 27072 16362 27124
rect 16758 27072 16764 27124
rect 16816 27112 16822 27124
rect 16853 27115 16911 27121
rect 16853 27112 16865 27115
rect 16816 27084 16865 27112
rect 16816 27072 16822 27084
rect 16853 27081 16865 27084
rect 16899 27081 16911 27115
rect 16853 27075 16911 27081
rect 16942 27072 16948 27124
rect 17000 27112 17006 27124
rect 17313 27115 17371 27121
rect 17313 27112 17325 27115
rect 17000 27084 17325 27112
rect 17000 27072 17006 27084
rect 17313 27081 17325 27084
rect 17359 27081 17371 27115
rect 17313 27075 17371 27081
rect 18322 27072 18328 27124
rect 18380 27112 18386 27124
rect 19426 27112 19432 27124
rect 18380 27084 19432 27112
rect 18380 27072 18386 27084
rect 19426 27072 19432 27084
rect 19484 27072 19490 27124
rect 19518 27072 19524 27124
rect 19576 27112 19582 27124
rect 19797 27115 19855 27121
rect 19797 27112 19809 27115
rect 19576 27084 19809 27112
rect 19576 27072 19582 27084
rect 19797 27081 19809 27084
rect 19843 27081 19855 27115
rect 20622 27112 20628 27124
rect 19797 27075 19855 27081
rect 19996 27084 20628 27112
rect 12710 27044 12716 27056
rect 9232 27016 12716 27044
rect 9125 27007 9183 27013
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 14550 27004 14556 27056
rect 14608 27044 14614 27056
rect 14645 27047 14703 27053
rect 14645 27044 14657 27047
rect 14608 27016 14657 27044
rect 14608 27004 14614 27016
rect 14645 27013 14657 27016
rect 14691 27013 14703 27047
rect 14645 27007 14703 27013
rect 14829 27047 14887 27053
rect 14829 27013 14841 27047
rect 14875 27044 14887 27047
rect 15930 27044 15936 27056
rect 14875 27016 15936 27044
rect 14875 27013 14887 27016
rect 14829 27007 14887 27013
rect 15930 27004 15936 27016
rect 15988 27004 15994 27056
rect 16393 27047 16451 27053
rect 16393 27013 16405 27047
rect 16439 27044 16451 27047
rect 17862 27044 17868 27056
rect 16439 27016 17868 27044
rect 16439 27013 16451 27016
rect 16393 27007 16451 27013
rect 17862 27004 17868 27016
rect 17920 27004 17926 27056
rect 18049 27047 18107 27053
rect 18049 27013 18061 27047
rect 18095 27044 18107 27047
rect 18874 27044 18880 27056
rect 18095 27016 18880 27044
rect 18095 27013 18107 27016
rect 18049 27007 18107 27013
rect 18874 27004 18880 27016
rect 18932 27004 18938 27056
rect 19996 27053 20024 27084
rect 20622 27072 20628 27084
rect 20680 27112 20686 27124
rect 20809 27115 20867 27121
rect 20809 27112 20821 27115
rect 20680 27084 20821 27112
rect 20680 27072 20686 27084
rect 20809 27081 20821 27084
rect 20855 27081 20867 27115
rect 20809 27075 20867 27081
rect 21818 27072 21824 27124
rect 21876 27112 21882 27124
rect 22849 27115 22907 27121
rect 22849 27112 22861 27115
rect 21876 27084 22861 27112
rect 21876 27072 21882 27084
rect 22849 27081 22861 27084
rect 22895 27081 22907 27115
rect 22849 27075 22907 27081
rect 23014 27072 23020 27124
rect 23072 27072 23078 27124
rect 25222 27072 25228 27124
rect 25280 27112 25286 27124
rect 25501 27115 25559 27121
rect 25501 27112 25513 27115
rect 25280 27084 25513 27112
rect 25280 27072 25286 27084
rect 25501 27081 25513 27084
rect 25547 27081 25559 27115
rect 25501 27075 25559 27081
rect 27154 27072 27160 27124
rect 27212 27112 27218 27124
rect 28169 27115 28227 27121
rect 28169 27112 28181 27115
rect 27212 27084 28181 27112
rect 27212 27072 27218 27084
rect 28169 27081 28181 27084
rect 28215 27112 28227 27115
rect 29178 27112 29184 27124
rect 28215 27084 29184 27112
rect 28215 27081 28227 27084
rect 28169 27075 28227 27081
rect 29178 27072 29184 27084
rect 29236 27072 29242 27124
rect 29638 27072 29644 27124
rect 29696 27112 29702 27124
rect 32122 27112 32128 27124
rect 29696 27084 32128 27112
rect 29696 27072 29702 27084
rect 32122 27072 32128 27084
rect 32180 27072 32186 27124
rect 33137 27115 33195 27121
rect 33137 27081 33149 27115
rect 33183 27112 33195 27115
rect 34422 27112 34428 27124
rect 33183 27084 34428 27112
rect 33183 27081 33195 27084
rect 33137 27075 33195 27081
rect 34422 27072 34428 27084
rect 34480 27072 34486 27124
rect 35802 27112 35808 27124
rect 34900 27084 35808 27112
rect 19981 27047 20039 27053
rect 19981 27013 19993 27047
rect 20027 27013 20039 27047
rect 20530 27044 20536 27056
rect 19981 27007 20039 27013
rect 20088 27016 20536 27044
rect 4341 26979 4399 26985
rect 4341 26945 4353 26979
rect 4387 26945 4399 26979
rect 4341 26939 4399 26945
rect 4617 26979 4675 26985
rect 4617 26945 4629 26979
rect 4663 26945 4675 26979
rect 4617 26939 4675 26945
rect 4709 26979 4767 26985
rect 4709 26945 4721 26979
rect 4755 26976 4767 26979
rect 4893 26979 4951 26985
rect 4755 26948 4844 26976
rect 4755 26945 4767 26948
rect 4709 26939 4767 26945
rect 2409 26911 2467 26917
rect 2409 26877 2421 26911
rect 2455 26908 2467 26911
rect 2774 26908 2780 26920
rect 2455 26880 2780 26908
rect 2455 26877 2467 26880
rect 2409 26871 2467 26877
rect 2774 26868 2780 26880
rect 2832 26868 2838 26920
rect 4249 26911 4307 26917
rect 4249 26877 4261 26911
rect 4295 26908 4307 26911
rect 4632 26908 4660 26939
rect 4295 26880 4660 26908
rect 4295 26877 4307 26880
rect 4249 26871 4307 26877
rect 3418 26800 3424 26852
rect 3476 26840 3482 26852
rect 4433 26843 4491 26849
rect 4433 26840 4445 26843
rect 3476 26812 4445 26840
rect 3476 26800 3482 26812
rect 4433 26809 4445 26812
rect 4479 26809 4491 26843
rect 4632 26840 4660 26880
rect 4706 26840 4712 26852
rect 4632 26812 4712 26840
rect 4433 26803 4491 26809
rect 4706 26800 4712 26812
rect 4764 26800 4770 26852
rect 4816 26840 4844 26948
rect 4893 26945 4905 26979
rect 4939 26945 4951 26979
rect 4893 26939 4951 26945
rect 4908 26908 4936 26939
rect 4982 26936 4988 26988
rect 5040 26936 5046 26988
rect 6546 26936 6552 26988
rect 6604 26976 6610 26988
rect 8941 26979 8999 26985
rect 8941 26976 8953 26979
rect 6604 26948 8953 26976
rect 6604 26936 6610 26948
rect 8941 26945 8953 26948
rect 8987 26945 8999 26979
rect 8941 26939 8999 26945
rect 9490 26936 9496 26988
rect 9548 26976 9554 26988
rect 10514 26979 10572 26985
rect 10514 26976 10526 26979
rect 9548 26948 10526 26976
rect 9548 26936 9554 26948
rect 10514 26945 10526 26948
rect 10560 26945 10572 26979
rect 10514 26939 10572 26945
rect 10686 26936 10692 26988
rect 10744 26976 10750 26988
rect 10781 26979 10839 26985
rect 10781 26976 10793 26979
rect 10744 26948 10793 26976
rect 10744 26936 10750 26948
rect 10781 26945 10793 26948
rect 10827 26976 10839 26979
rect 10870 26976 10876 26988
rect 10827 26948 10876 26976
rect 10827 26945 10839 26948
rect 10781 26939 10839 26945
rect 10870 26936 10876 26948
rect 10928 26936 10934 26988
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26945 11943 26979
rect 11885 26939 11943 26945
rect 15105 26979 15163 26985
rect 15105 26945 15117 26979
rect 15151 26976 15163 26979
rect 16298 26976 16304 26988
rect 15151 26948 16304 26976
rect 15151 26945 15163 26948
rect 15105 26939 15163 26945
rect 5626 26908 5632 26920
rect 4908 26880 5632 26908
rect 5626 26868 5632 26880
rect 5684 26868 5690 26920
rect 5534 26840 5540 26852
rect 4816 26812 5540 26840
rect 5534 26800 5540 26812
rect 5592 26840 5598 26852
rect 5718 26840 5724 26852
rect 5592 26812 5724 26840
rect 5592 26800 5598 26812
rect 5718 26800 5724 26812
rect 5776 26800 5782 26852
rect 2866 26732 2872 26784
rect 2924 26772 2930 26784
rect 2961 26775 3019 26781
rect 2961 26772 2973 26775
rect 2924 26744 2973 26772
rect 2924 26732 2930 26744
rect 2961 26741 2973 26744
rect 3007 26741 3019 26775
rect 2961 26735 3019 26741
rect 4522 26732 4528 26784
rect 4580 26772 4586 26784
rect 4982 26772 4988 26784
rect 4580 26744 4988 26772
rect 4580 26732 4586 26744
rect 4982 26732 4988 26744
rect 5040 26772 5046 26784
rect 5442 26772 5448 26784
rect 5040 26744 5448 26772
rect 5040 26732 5046 26744
rect 5442 26732 5448 26744
rect 5500 26732 5506 26784
rect 8662 26732 8668 26784
rect 8720 26772 8726 26784
rect 9398 26772 9404 26784
rect 8720 26744 9404 26772
rect 8720 26732 8726 26744
rect 9398 26732 9404 26744
rect 9456 26732 9462 26784
rect 10134 26732 10140 26784
rect 10192 26772 10198 26784
rect 11900 26772 11928 26939
rect 16298 26936 16304 26948
rect 16356 26936 16362 26988
rect 16850 26936 16856 26988
rect 16908 26976 16914 26988
rect 17770 26976 17776 26988
rect 16908 26948 17776 26976
rect 16908 26936 16914 26948
rect 17770 26936 17776 26948
rect 17828 26936 17834 26988
rect 17954 26936 17960 26988
rect 18012 26936 18018 26988
rect 18138 26936 18144 26988
rect 18196 26976 18202 26988
rect 18233 26979 18291 26985
rect 18233 26976 18245 26979
rect 18196 26948 18245 26976
rect 18196 26936 18202 26948
rect 18233 26945 18245 26948
rect 18279 26945 18291 26979
rect 18233 26939 18291 26945
rect 18414 26936 18420 26988
rect 18472 26976 18478 26988
rect 18966 26976 18972 26988
rect 18472 26948 18972 26976
rect 18472 26936 18478 26948
rect 18966 26936 18972 26948
rect 19024 26936 19030 26988
rect 19150 26936 19156 26988
rect 19208 26976 19214 26988
rect 19337 26979 19395 26985
rect 19337 26976 19349 26979
rect 19208 26948 19349 26976
rect 19208 26936 19214 26948
rect 19337 26945 19349 26948
rect 19383 26945 19395 26979
rect 19337 26939 19395 26945
rect 19886 26936 19892 26988
rect 19944 26976 19950 26988
rect 20088 26976 20116 27016
rect 20530 27004 20536 27016
rect 20588 27044 20594 27056
rect 20717 27047 20775 27053
rect 20717 27044 20729 27047
rect 20588 27016 20729 27044
rect 20588 27004 20594 27016
rect 20717 27013 20729 27016
rect 20763 27013 20775 27047
rect 22649 27047 22707 27053
rect 22649 27044 22661 27047
rect 20717 27007 20775 27013
rect 22066 27016 22661 27044
rect 20441 26979 20499 26985
rect 20441 26976 20453 26979
rect 19944 26948 20116 26976
rect 20272 26948 20453 26976
rect 19944 26936 19950 26948
rect 12066 26868 12072 26920
rect 12124 26868 12130 26920
rect 15197 26911 15255 26917
rect 15197 26877 15209 26911
rect 15243 26908 15255 26911
rect 15378 26908 15384 26920
rect 15243 26880 15384 26908
rect 15243 26877 15255 26880
rect 15197 26871 15255 26877
rect 15378 26868 15384 26880
rect 15436 26868 15442 26920
rect 16666 26868 16672 26920
rect 16724 26868 16730 26920
rect 16761 26911 16819 26917
rect 16761 26877 16773 26911
rect 16807 26908 16819 26911
rect 16942 26908 16948 26920
rect 16807 26880 16948 26908
rect 16807 26877 16819 26880
rect 16761 26871 16819 26877
rect 12618 26800 12624 26852
rect 12676 26840 12682 26852
rect 15746 26840 15752 26852
rect 12676 26812 15752 26840
rect 12676 26800 12682 26812
rect 15746 26800 15752 26812
rect 15804 26840 15810 26852
rect 16776 26840 16804 26871
rect 16942 26868 16948 26880
rect 17000 26868 17006 26920
rect 17037 26911 17095 26917
rect 17037 26877 17049 26911
rect 17083 26877 17095 26911
rect 17037 26871 17095 26877
rect 17129 26911 17187 26917
rect 17129 26877 17141 26911
rect 17175 26908 17187 26911
rect 17310 26908 17316 26920
rect 17175 26880 17316 26908
rect 17175 26877 17187 26880
rect 17129 26871 17187 26877
rect 15804 26812 16804 26840
rect 15804 26800 15810 26812
rect 10192 26744 11928 26772
rect 10192 26732 10198 26744
rect 14826 26732 14832 26784
rect 14884 26772 14890 26784
rect 15105 26775 15163 26781
rect 15105 26772 15117 26775
rect 14884 26744 15117 26772
rect 14884 26732 14890 26744
rect 15105 26741 15117 26744
rect 15151 26741 15163 26775
rect 15105 26735 15163 26741
rect 15286 26732 15292 26784
rect 15344 26772 15350 26784
rect 15838 26772 15844 26784
rect 15344 26744 15844 26772
rect 15344 26732 15350 26744
rect 15838 26732 15844 26744
rect 15896 26732 15902 26784
rect 16942 26732 16948 26784
rect 17000 26772 17006 26784
rect 17052 26772 17080 26871
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 18322 26868 18328 26920
rect 18380 26908 18386 26920
rect 19429 26911 19487 26917
rect 19429 26908 19441 26911
rect 18380 26880 19441 26908
rect 18380 26868 18386 26880
rect 19429 26877 19441 26880
rect 19475 26908 19487 26911
rect 19613 26911 19671 26917
rect 19613 26908 19625 26911
rect 19475 26880 19625 26908
rect 19475 26877 19487 26880
rect 19429 26871 19487 26877
rect 19613 26877 19625 26880
rect 19659 26908 19671 26911
rect 20272 26908 20300 26948
rect 20441 26945 20453 26948
rect 20487 26945 20499 26979
rect 20441 26939 20499 26945
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26976 20683 26979
rect 22066 26976 22094 27016
rect 22649 27013 22661 27016
rect 22695 27013 22707 27047
rect 22649 27007 22707 27013
rect 24121 27047 24179 27053
rect 24121 27013 24133 27047
rect 24167 27044 24179 27047
rect 26694 27044 26700 27056
rect 24167 27016 26700 27044
rect 24167 27013 24179 27016
rect 24121 27007 24179 27013
rect 26694 27004 26700 27016
rect 26752 27004 26758 27056
rect 29656 27044 29684 27072
rect 28092 27016 29684 27044
rect 20671 26948 22094 26976
rect 23385 26979 23443 26985
rect 20671 26945 20683 26948
rect 20625 26939 20683 26945
rect 23385 26945 23397 26979
rect 23431 26976 23443 26979
rect 23474 26976 23480 26988
rect 23431 26948 23480 26976
rect 23431 26945 23443 26948
rect 23385 26939 23443 26945
rect 19659 26880 20300 26908
rect 20349 26911 20407 26917
rect 19659 26877 19671 26880
rect 19613 26871 19671 26877
rect 20349 26877 20361 26911
rect 20395 26877 20407 26911
rect 20640 26908 20668 26939
rect 23474 26936 23480 26948
rect 23532 26976 23538 26988
rect 24394 26976 24400 26988
rect 23532 26948 24400 26976
rect 23532 26936 23538 26948
rect 24394 26936 24400 26948
rect 24452 26936 24458 26988
rect 25498 26936 25504 26988
rect 25556 26976 25562 26988
rect 25593 26979 25651 26985
rect 25593 26976 25605 26979
rect 25556 26948 25605 26976
rect 25556 26936 25562 26948
rect 25593 26945 25605 26948
rect 25639 26945 25651 26979
rect 25593 26939 25651 26945
rect 26145 26979 26203 26985
rect 26145 26945 26157 26979
rect 26191 26945 26203 26979
rect 26145 26939 26203 26945
rect 26329 26979 26387 26985
rect 26329 26945 26341 26979
rect 26375 26945 26387 26979
rect 26329 26939 26387 26945
rect 20349 26871 20407 26877
rect 20456 26880 20668 26908
rect 17494 26800 17500 26852
rect 17552 26840 17558 26852
rect 18233 26843 18291 26849
rect 18233 26840 18245 26843
rect 17552 26812 18245 26840
rect 17552 26800 17558 26812
rect 18233 26809 18245 26812
rect 18279 26809 18291 26843
rect 18233 26803 18291 26809
rect 18598 26800 18604 26852
rect 18656 26840 18662 26852
rect 18656 26812 19012 26840
rect 18656 26800 18662 26812
rect 17000 26744 17080 26772
rect 17589 26775 17647 26781
rect 17000 26732 17006 26744
rect 17589 26741 17601 26775
rect 17635 26772 17647 26775
rect 17678 26772 17684 26784
rect 17635 26744 17684 26772
rect 17635 26741 17647 26744
rect 17589 26735 17647 26741
rect 17678 26732 17684 26744
rect 17736 26732 17742 26784
rect 17770 26732 17776 26784
rect 17828 26772 17834 26784
rect 18616 26772 18644 26800
rect 17828 26744 18644 26772
rect 17828 26732 17834 26744
rect 18690 26732 18696 26784
rect 18748 26772 18754 26784
rect 18984 26781 19012 26812
rect 20254 26800 20260 26852
rect 20312 26840 20318 26852
rect 20364 26840 20392 26871
rect 20456 26852 20484 26880
rect 20714 26868 20720 26920
rect 20772 26908 20778 26920
rect 20993 26911 21051 26917
rect 20993 26908 21005 26911
rect 20772 26880 21005 26908
rect 20772 26868 20778 26880
rect 20993 26877 21005 26880
rect 21039 26877 21051 26911
rect 20993 26871 21051 26877
rect 21174 26868 21180 26920
rect 21232 26908 21238 26920
rect 22554 26908 22560 26920
rect 21232 26880 22560 26908
rect 21232 26868 21238 26880
rect 22554 26868 22560 26880
rect 22612 26868 22618 26920
rect 23106 26868 23112 26920
rect 23164 26908 23170 26920
rect 23164 26880 24801 26908
rect 23164 26868 23170 26880
rect 20312 26812 20392 26840
rect 20312 26800 20318 26812
rect 20438 26800 20444 26852
rect 20496 26800 20502 26852
rect 20806 26800 20812 26852
rect 20864 26840 20870 26852
rect 22094 26840 22100 26852
rect 20864 26812 22100 26840
rect 20864 26800 20870 26812
rect 22066 26800 22100 26812
rect 22152 26800 22158 26852
rect 24773 26840 24801 26880
rect 25314 26868 25320 26920
rect 25372 26868 25378 26920
rect 25406 26868 25412 26920
rect 25464 26908 25470 26920
rect 25774 26908 25780 26920
rect 25464 26880 25780 26908
rect 25464 26868 25470 26880
rect 25774 26868 25780 26880
rect 25832 26908 25838 26920
rect 26160 26908 26188 26939
rect 25832 26880 26188 26908
rect 26344 26908 26372 26939
rect 26418 26936 26424 26988
rect 26476 26936 26482 26988
rect 26510 26936 26516 26988
rect 26568 26936 26574 26988
rect 27890 26908 27896 26920
rect 26344 26880 27896 26908
rect 25832 26868 25838 26880
rect 27890 26868 27896 26880
rect 27948 26868 27954 26920
rect 28092 26917 28120 27016
rect 29730 27004 29736 27056
rect 29788 27044 29794 27056
rect 30650 27044 30656 27056
rect 29788 27016 30656 27044
rect 29788 27004 29794 27016
rect 30650 27004 30656 27016
rect 30708 27004 30714 27056
rect 33870 27004 33876 27056
rect 33928 27004 33934 27056
rect 34514 27004 34520 27056
rect 34572 27044 34578 27056
rect 34609 27047 34667 27053
rect 34609 27044 34621 27047
rect 34572 27016 34621 27044
rect 34572 27004 34578 27016
rect 34609 27013 34621 27016
rect 34655 27013 34667 27047
rect 34609 27007 34667 27013
rect 28261 26979 28319 26985
rect 28261 26945 28273 26979
rect 28307 26976 28319 26979
rect 28350 26976 28356 26988
rect 28307 26948 28356 26976
rect 28307 26945 28319 26948
rect 28261 26939 28319 26945
rect 28350 26936 28356 26948
rect 28408 26936 28414 26988
rect 28721 26979 28779 26985
rect 28721 26976 28733 26979
rect 28460 26948 28733 26976
rect 28077 26911 28135 26917
rect 28077 26877 28089 26911
rect 28123 26877 28135 26911
rect 28077 26871 28135 26877
rect 24773 26812 26832 26840
rect 18785 26775 18843 26781
rect 18785 26772 18797 26775
rect 18748 26744 18797 26772
rect 18748 26732 18754 26744
rect 18785 26741 18797 26744
rect 18831 26741 18843 26775
rect 18785 26735 18843 26741
rect 18969 26775 19027 26781
rect 18969 26741 18981 26775
rect 19015 26741 19027 26775
rect 22066 26772 22094 26800
rect 22462 26772 22468 26784
rect 22066 26744 22468 26772
rect 18969 26735 19027 26741
rect 22462 26732 22468 26744
rect 22520 26732 22526 26784
rect 22833 26775 22891 26781
rect 22833 26741 22845 26775
rect 22879 26772 22891 26775
rect 22922 26772 22928 26784
rect 22879 26744 22928 26772
rect 22879 26741 22891 26744
rect 22833 26735 22891 26741
rect 22922 26732 22928 26744
rect 22980 26732 22986 26784
rect 23106 26732 23112 26784
rect 23164 26772 23170 26784
rect 24210 26772 24216 26784
rect 23164 26744 24216 26772
rect 23164 26732 23170 26744
rect 24210 26732 24216 26744
rect 24268 26732 24274 26784
rect 25590 26732 25596 26784
rect 25648 26772 25654 26784
rect 25961 26775 26019 26781
rect 25961 26772 25973 26775
rect 25648 26744 25973 26772
rect 25648 26732 25654 26744
rect 25961 26741 25973 26744
rect 26007 26741 26019 26775
rect 25961 26735 26019 26741
rect 26694 26732 26700 26784
rect 26752 26732 26758 26784
rect 26804 26772 26832 26812
rect 27798 26800 27804 26852
rect 27856 26840 27862 26852
rect 28460 26840 28488 26948
rect 28721 26945 28733 26948
rect 28767 26945 28779 26979
rect 28721 26939 28779 26945
rect 28902 26936 28908 26988
rect 28960 26936 28966 26988
rect 28994 26936 29000 26988
rect 29052 26936 29058 26988
rect 29089 26979 29147 26985
rect 29089 26945 29101 26979
rect 29135 26945 29147 26979
rect 29089 26939 29147 26945
rect 28810 26868 28816 26920
rect 28868 26908 28874 26920
rect 29104 26908 29132 26939
rect 29914 26936 29920 26988
rect 29972 26936 29978 26988
rect 34900 26985 34928 27084
rect 35802 27072 35808 27084
rect 35860 27072 35866 27124
rect 36262 27112 36268 27124
rect 35912 27084 36268 27112
rect 35526 27004 35532 27056
rect 35584 27004 35590 27056
rect 34885 26979 34943 26985
rect 34885 26945 34897 26979
rect 34931 26945 34943 26979
rect 35391 26979 35449 26985
rect 35391 26976 35403 26979
rect 34885 26939 34943 26945
rect 35268 26948 35403 26976
rect 32125 26911 32183 26917
rect 32125 26908 32137 26911
rect 28868 26880 29132 26908
rect 29196 26880 32137 26908
rect 28868 26868 28874 26880
rect 29196 26840 29224 26880
rect 32125 26877 32137 26880
rect 32171 26877 32183 26911
rect 32125 26871 32183 26877
rect 32401 26911 32459 26917
rect 32401 26877 32413 26911
rect 32447 26908 32459 26911
rect 32766 26908 32772 26920
rect 32447 26880 32772 26908
rect 32447 26877 32459 26880
rect 32401 26871 32459 26877
rect 32766 26868 32772 26880
rect 32824 26868 32830 26920
rect 33594 26868 33600 26920
rect 33652 26908 33658 26920
rect 34054 26908 34060 26920
rect 33652 26880 34060 26908
rect 33652 26868 33658 26880
rect 34054 26868 34060 26880
rect 34112 26868 34118 26920
rect 34514 26868 34520 26920
rect 34572 26908 34578 26920
rect 34900 26908 34928 26939
rect 34572 26880 34928 26908
rect 35268 26908 35296 26948
rect 35391 26945 35403 26948
rect 35437 26945 35449 26979
rect 35391 26939 35449 26945
rect 35618 26936 35624 26988
rect 35676 26936 35682 26988
rect 35912 26985 35940 27084
rect 36262 27072 36268 27084
rect 36320 27072 36326 27124
rect 36630 27072 36636 27124
rect 36688 27072 36694 27124
rect 37734 27072 37740 27124
rect 37792 27112 37798 27124
rect 40034 27112 40040 27124
rect 37792 27084 40040 27112
rect 37792 27072 37798 27084
rect 40034 27072 40040 27084
rect 40092 27072 40098 27124
rect 40129 27115 40187 27121
rect 40129 27081 40141 27115
rect 40175 27112 40187 27115
rect 40862 27112 40868 27124
rect 40175 27084 40868 27112
rect 40175 27081 40187 27084
rect 40129 27075 40187 27081
rect 40862 27072 40868 27084
rect 40920 27112 40926 27124
rect 41598 27112 41604 27124
rect 40920 27084 41604 27112
rect 40920 27072 40926 27084
rect 41598 27072 41604 27084
rect 41656 27072 41662 27124
rect 36538 27044 36544 27056
rect 36280 27016 36544 27044
rect 36170 26985 36176 26988
rect 35804 26979 35862 26985
rect 35804 26945 35816 26979
rect 35850 26945 35862 26979
rect 35804 26939 35862 26945
rect 35897 26979 35955 26985
rect 35897 26945 35909 26979
rect 35943 26976 35955 26979
rect 35989 26979 36047 26985
rect 35989 26976 36001 26979
rect 35943 26948 36001 26976
rect 35943 26945 35955 26948
rect 35897 26939 35955 26945
rect 35989 26945 36001 26948
rect 36035 26945 36047 26979
rect 35989 26939 36047 26945
rect 36137 26979 36176 26985
rect 36137 26945 36149 26979
rect 36137 26939 36176 26945
rect 35820 26908 35848 26939
rect 36170 26936 36176 26939
rect 36228 26936 36234 26988
rect 36280 26985 36308 27016
rect 36538 27004 36544 27016
rect 36596 27004 36602 27056
rect 38378 27004 38384 27056
rect 38436 27004 38442 27056
rect 38473 27047 38531 27053
rect 38473 27013 38485 27047
rect 38519 27044 38531 27047
rect 38562 27044 38568 27056
rect 38519 27016 38568 27044
rect 38519 27013 38531 27016
rect 38473 27007 38531 27013
rect 38562 27004 38568 27016
rect 38620 27004 38626 27056
rect 36265 26979 36323 26985
rect 36265 26945 36277 26979
rect 36311 26945 36323 26979
rect 36265 26939 36323 26945
rect 36354 26936 36360 26988
rect 36412 26936 36418 26988
rect 36446 26936 36452 26988
rect 36504 26985 36510 26988
rect 36504 26976 36512 26985
rect 36504 26948 36549 26976
rect 36504 26939 36512 26948
rect 36504 26936 36510 26939
rect 40586 26936 40592 26988
rect 40644 26936 40650 26988
rect 40770 26936 40776 26988
rect 40828 26936 40834 26988
rect 41046 26936 41052 26988
rect 41104 26976 41110 26988
rect 41877 26979 41935 26985
rect 41877 26976 41889 26979
rect 41104 26948 41889 26976
rect 41104 26936 41110 26948
rect 41877 26945 41889 26948
rect 41923 26945 41935 26979
rect 41877 26939 41935 26945
rect 36722 26908 36728 26920
rect 35268 26880 35480 26908
rect 35820 26880 36728 26908
rect 34572 26868 34578 26880
rect 27856 26812 28488 26840
rect 28552 26812 29224 26840
rect 27856 26800 27862 26812
rect 28552 26772 28580 26812
rect 35250 26800 35256 26852
rect 35308 26800 35314 26852
rect 26804 26744 28580 26772
rect 28629 26775 28687 26781
rect 28629 26741 28641 26775
rect 28675 26772 28687 26775
rect 28718 26772 28724 26784
rect 28675 26744 28724 26772
rect 28675 26741 28687 26744
rect 28629 26735 28687 26741
rect 28718 26732 28724 26744
rect 28776 26732 28782 26784
rect 29273 26775 29331 26781
rect 29273 26741 29285 26775
rect 29319 26772 29331 26775
rect 30006 26772 30012 26784
rect 29319 26744 30012 26772
rect 29319 26741 29331 26744
rect 29273 26735 29331 26741
rect 30006 26732 30012 26744
rect 30064 26732 30070 26784
rect 30190 26781 30196 26784
rect 30180 26775 30196 26781
rect 30180 26741 30192 26775
rect 30180 26735 30196 26741
rect 30190 26732 30196 26735
rect 30248 26732 30254 26784
rect 30650 26732 30656 26784
rect 30708 26772 30714 26784
rect 31202 26772 31208 26784
rect 30708 26744 31208 26772
rect 30708 26732 30714 26744
rect 31202 26732 31208 26744
rect 31260 26732 31266 26784
rect 31662 26772 31668 26784
rect 31623 26744 31668 26772
rect 31662 26732 31668 26744
rect 31720 26772 31726 26784
rect 34606 26772 34612 26784
rect 31720 26744 34612 26772
rect 31720 26732 31726 26744
rect 34606 26732 34612 26744
rect 34664 26732 34670 26784
rect 35452 26772 35480 26880
rect 36722 26868 36728 26880
rect 36780 26868 36786 26920
rect 38197 26911 38255 26917
rect 38197 26877 38209 26911
rect 38243 26877 38255 26911
rect 38197 26871 38255 26877
rect 39853 26911 39911 26917
rect 39853 26877 39865 26911
rect 39899 26877 39911 26911
rect 39853 26871 39911 26877
rect 35710 26800 35716 26852
rect 35768 26840 35774 26852
rect 37550 26840 37556 26852
rect 35768 26812 37556 26840
rect 35768 26800 35774 26812
rect 37550 26800 37556 26812
rect 37608 26840 37614 26852
rect 38212 26840 38240 26871
rect 39868 26840 39896 26871
rect 37608 26812 39896 26840
rect 40497 26843 40555 26849
rect 37608 26800 37614 26812
rect 40497 26809 40509 26843
rect 40543 26840 40555 26843
rect 41230 26840 41236 26852
rect 40543 26812 41236 26840
rect 40543 26809 40555 26812
rect 40497 26803 40555 26809
rect 41230 26800 41236 26812
rect 41288 26800 41294 26852
rect 36078 26772 36084 26784
rect 35452 26744 36084 26772
rect 36078 26732 36084 26744
rect 36136 26732 36142 26784
rect 38841 26775 38899 26781
rect 38841 26741 38853 26775
rect 38887 26772 38899 26775
rect 39206 26772 39212 26784
rect 38887 26744 39212 26772
rect 38887 26741 38899 26744
rect 38841 26735 38899 26741
rect 39206 26732 39212 26744
rect 39264 26732 39270 26784
rect 40678 26732 40684 26784
rect 40736 26772 40742 26784
rect 40957 26775 41015 26781
rect 40957 26772 40969 26775
rect 40736 26744 40969 26772
rect 40736 26732 40742 26744
rect 40957 26741 40969 26744
rect 41003 26741 41015 26775
rect 40957 26735 41015 26741
rect 42058 26732 42064 26784
rect 42116 26732 42122 26784
rect 1104 26682 42504 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 42504 26682
rect 1104 26608 42504 26630
rect 3255 26571 3313 26577
rect 3255 26537 3267 26571
rect 3301 26568 3313 26571
rect 3418 26568 3424 26580
rect 3301 26540 3424 26568
rect 3301 26537 3313 26540
rect 3255 26531 3313 26537
rect 3418 26528 3424 26540
rect 3476 26528 3482 26580
rect 4430 26528 4436 26580
rect 4488 26528 4494 26580
rect 4617 26571 4675 26577
rect 4617 26537 4629 26571
rect 4663 26568 4675 26571
rect 4706 26568 4712 26580
rect 4663 26540 4712 26568
rect 4663 26537 4675 26540
rect 4617 26531 4675 26537
rect 4706 26528 4712 26540
rect 4764 26528 4770 26580
rect 4893 26571 4951 26577
rect 4893 26537 4905 26571
rect 4939 26568 4951 26571
rect 5350 26568 5356 26580
rect 4939 26540 5356 26568
rect 4939 26537 4951 26540
rect 4893 26531 4951 26537
rect 5350 26528 5356 26540
rect 5408 26528 5414 26580
rect 8478 26528 8484 26580
rect 8536 26568 8542 26580
rect 9214 26568 9220 26580
rect 8536 26540 9220 26568
rect 8536 26528 8542 26540
rect 9214 26528 9220 26540
rect 9272 26528 9278 26580
rect 9490 26528 9496 26580
rect 9548 26528 9554 26580
rect 9582 26528 9588 26580
rect 9640 26568 9646 26580
rect 11330 26568 11336 26580
rect 9640 26540 11336 26568
rect 9640 26528 9646 26540
rect 11330 26528 11336 26540
rect 11388 26528 11394 26580
rect 12069 26571 12127 26577
rect 12069 26537 12081 26571
rect 12115 26568 12127 26571
rect 12158 26568 12164 26580
rect 12115 26540 12164 26568
rect 12115 26537 12127 26540
rect 12069 26531 12127 26537
rect 12158 26528 12164 26540
rect 12216 26568 12222 26580
rect 12986 26568 12992 26580
rect 12216 26540 12992 26568
rect 12216 26528 12222 26540
rect 12986 26528 12992 26540
rect 13044 26528 13050 26580
rect 14918 26528 14924 26580
rect 14976 26568 14982 26580
rect 15013 26571 15071 26577
rect 15013 26568 15025 26571
rect 14976 26540 15025 26568
rect 14976 26528 14982 26540
rect 15013 26537 15025 26540
rect 15059 26537 15071 26571
rect 15013 26531 15071 26537
rect 15856 26540 16068 26568
rect 7926 26460 7932 26512
rect 7984 26460 7990 26512
rect 8757 26503 8815 26509
rect 8757 26469 8769 26503
rect 8803 26500 8815 26503
rect 10226 26500 10232 26512
rect 8803 26472 10232 26500
rect 8803 26469 8815 26472
rect 8757 26463 8815 26469
rect 10226 26460 10232 26472
rect 10284 26460 10290 26512
rect 15856 26500 15884 26540
rect 13832 26472 15884 26500
rect 16040 26500 16068 26540
rect 16298 26528 16304 26580
rect 16356 26568 16362 26580
rect 16485 26571 16543 26577
rect 16485 26568 16497 26571
rect 16356 26540 16497 26568
rect 16356 26528 16362 26540
rect 16485 26537 16497 26540
rect 16531 26537 16543 26571
rect 16485 26531 16543 26537
rect 17954 26528 17960 26580
rect 18012 26568 18018 26580
rect 18417 26571 18475 26577
rect 18417 26568 18429 26571
rect 18012 26540 18429 26568
rect 18012 26528 18018 26540
rect 18417 26537 18429 26540
rect 18463 26537 18475 26571
rect 18417 26531 18475 26537
rect 20438 26528 20444 26580
rect 20496 26568 20502 26580
rect 20809 26571 20867 26577
rect 20809 26568 20821 26571
rect 20496 26540 20821 26568
rect 20496 26528 20502 26540
rect 20809 26537 20821 26540
rect 20855 26537 20867 26571
rect 20809 26531 20867 26537
rect 21192 26540 22508 26568
rect 16945 26503 17003 26509
rect 16945 26500 16957 26503
rect 16040 26472 16957 26500
rect 1489 26435 1547 26441
rect 1489 26401 1501 26435
rect 1535 26432 1547 26435
rect 2774 26432 2780 26444
rect 1535 26404 2780 26432
rect 1535 26401 1547 26404
rect 1489 26395 1547 26401
rect 2774 26392 2780 26404
rect 2832 26392 2838 26444
rect 7006 26432 7012 26444
rect 5276 26404 7012 26432
rect 3510 26324 3516 26376
rect 3568 26324 3574 26376
rect 3970 26324 3976 26376
rect 4028 26364 4034 26376
rect 4065 26367 4123 26373
rect 4065 26364 4077 26367
rect 4028 26336 4077 26364
rect 4028 26324 4034 26336
rect 4065 26333 4077 26336
rect 4111 26333 4123 26367
rect 4890 26364 4896 26376
rect 4065 26327 4123 26333
rect 4540 26336 4896 26364
rect 2958 26296 2964 26308
rect 2806 26268 2964 26296
rect 2958 26256 2964 26268
rect 3016 26256 3022 26308
rect 4540 26240 4568 26336
rect 4890 26324 4896 26336
rect 4948 26324 4954 26376
rect 5074 26373 5080 26376
rect 5072 26364 5080 26373
rect 5035 26336 5080 26364
rect 5072 26327 5080 26336
rect 5074 26324 5080 26327
rect 5132 26324 5138 26376
rect 5276 26373 5304 26404
rect 7006 26392 7012 26404
rect 7064 26392 7070 26444
rect 7944 26432 7972 26460
rect 10134 26432 10140 26444
rect 7944 26404 9168 26432
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5444 26367 5502 26373
rect 5444 26333 5456 26367
rect 5490 26333 5502 26367
rect 5444 26327 5502 26333
rect 4798 26256 4804 26308
rect 4856 26296 4862 26308
rect 5169 26299 5227 26305
rect 5169 26296 5181 26299
rect 4856 26268 5181 26296
rect 4856 26256 4862 26268
rect 5169 26265 5181 26268
rect 5215 26265 5227 26299
rect 5169 26259 5227 26265
rect 5459 26240 5487 26327
rect 5534 26324 5540 26376
rect 5592 26324 5598 26376
rect 5718 26324 5724 26376
rect 5776 26324 5782 26376
rect 5813 26367 5871 26373
rect 5813 26333 5825 26367
rect 5859 26364 5871 26367
rect 5994 26364 6000 26376
rect 5859 26336 6000 26364
rect 5859 26333 5871 26336
rect 5813 26327 5871 26333
rect 5994 26324 6000 26336
rect 6052 26324 6058 26376
rect 6178 26324 6184 26376
rect 6236 26324 6242 26376
rect 6638 26324 6644 26376
rect 6696 26324 6702 26376
rect 6914 26324 6920 26376
rect 6972 26324 6978 26376
rect 7190 26324 7196 26376
rect 7248 26364 7254 26376
rect 7285 26367 7343 26373
rect 7285 26364 7297 26367
rect 7248 26336 7297 26364
rect 7248 26324 7254 26336
rect 7285 26333 7297 26336
rect 7331 26333 7343 26367
rect 7285 26327 7343 26333
rect 8021 26367 8079 26373
rect 8021 26333 8033 26367
rect 8067 26333 8079 26367
rect 8021 26327 8079 26333
rect 8205 26367 8263 26373
rect 8205 26333 8217 26367
rect 8251 26364 8263 26367
rect 8294 26364 8300 26376
rect 8251 26336 8300 26364
rect 8251 26333 8263 26336
rect 8205 26327 8263 26333
rect 7208 26296 7236 26324
rect 6012 26268 7236 26296
rect 8036 26296 8064 26327
rect 8294 26324 8300 26336
rect 8352 26324 8358 26376
rect 8404 26373 8432 26404
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26333 8447 26367
rect 8389 26327 8447 26333
rect 8478 26324 8484 26376
rect 8536 26324 8542 26376
rect 8573 26367 8631 26373
rect 8573 26333 8585 26367
rect 8619 26333 8631 26367
rect 8573 26327 8631 26333
rect 8496 26296 8524 26324
rect 8036 26268 8524 26296
rect 8588 26296 8616 26327
rect 8938 26324 8944 26376
rect 8996 26324 9002 26376
rect 9140 26373 9168 26404
rect 9324 26404 10140 26432
rect 9125 26367 9183 26373
rect 9125 26333 9137 26367
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 9214 26324 9220 26376
rect 9272 26324 9278 26376
rect 9324 26373 9352 26404
rect 10134 26392 10140 26404
rect 10192 26392 10198 26444
rect 10321 26435 10379 26441
rect 10321 26401 10333 26435
rect 10367 26432 10379 26435
rect 10686 26432 10692 26444
rect 10367 26404 10692 26432
rect 10367 26401 10379 26404
rect 10321 26395 10379 26401
rect 10686 26392 10692 26404
rect 10744 26392 10750 26444
rect 13170 26432 13176 26444
rect 11716 26404 13176 26432
rect 9309 26367 9367 26373
rect 9309 26333 9321 26367
rect 9355 26333 9367 26367
rect 9309 26327 9367 26333
rect 9582 26324 9588 26376
rect 9640 26324 9646 26376
rect 11716 26350 11744 26404
rect 13170 26392 13176 26404
rect 13228 26392 13234 26444
rect 13633 26435 13691 26441
rect 13633 26401 13645 26435
rect 13679 26432 13691 26435
rect 13832 26432 13860 26472
rect 16945 26469 16957 26472
rect 16991 26469 17003 26503
rect 16945 26463 17003 26469
rect 17402 26460 17408 26512
rect 17460 26500 17466 26512
rect 18322 26500 18328 26512
rect 17460 26472 18328 26500
rect 17460 26460 17466 26472
rect 18322 26460 18328 26472
rect 18380 26460 18386 26512
rect 18966 26460 18972 26512
rect 19024 26500 19030 26512
rect 19024 26472 20944 26500
rect 19024 26460 19030 26472
rect 13679 26404 13860 26432
rect 13679 26401 13691 26404
rect 13633 26395 13691 26401
rect 13906 26392 13912 26444
rect 13964 26392 13970 26444
rect 14918 26392 14924 26444
rect 14976 26432 14982 26444
rect 15381 26435 15439 26441
rect 15381 26432 15393 26435
rect 14976 26404 15393 26432
rect 14976 26392 14982 26404
rect 15381 26401 15393 26404
rect 15427 26401 15439 26435
rect 15381 26395 15439 26401
rect 15470 26392 15476 26444
rect 15528 26392 15534 26444
rect 16390 26392 16396 26444
rect 16448 26432 16454 26444
rect 16669 26435 16727 26441
rect 16669 26432 16681 26435
rect 16448 26404 16681 26432
rect 16448 26392 16454 26404
rect 16669 26401 16681 26404
rect 16715 26432 16727 26435
rect 16850 26432 16856 26444
rect 16715 26404 16856 26432
rect 16715 26401 16727 26404
rect 16669 26395 16727 26401
rect 16850 26392 16856 26404
rect 16908 26392 16914 26444
rect 17129 26435 17187 26441
rect 17129 26401 17141 26435
rect 17175 26432 17187 26435
rect 18138 26432 18144 26444
rect 17175 26404 18144 26432
rect 17175 26401 17187 26404
rect 17129 26395 17187 26401
rect 18138 26392 18144 26404
rect 18196 26392 18202 26444
rect 18230 26392 18236 26444
rect 18288 26432 18294 26444
rect 19720 26441 19748 26472
rect 19245 26435 19303 26441
rect 19245 26432 19257 26435
rect 18288 26404 19257 26432
rect 18288 26392 18294 26404
rect 19245 26401 19257 26404
rect 19291 26401 19303 26435
rect 19245 26395 19303 26401
rect 19705 26435 19763 26441
rect 19705 26401 19717 26435
rect 19751 26401 19763 26435
rect 19705 26395 19763 26401
rect 19797 26435 19855 26441
rect 19797 26401 19809 26435
rect 19843 26432 19855 26435
rect 20254 26432 20260 26444
rect 19843 26404 20260 26432
rect 19843 26401 19855 26404
rect 19797 26395 19855 26401
rect 15289 26367 15347 26373
rect 15289 26333 15301 26367
rect 15335 26364 15347 26367
rect 15654 26364 15660 26376
rect 15335 26336 15660 26364
rect 15335 26333 15347 26336
rect 15289 26327 15347 26333
rect 15654 26324 15660 26336
rect 15712 26324 15718 26376
rect 15746 26324 15752 26376
rect 15804 26324 15810 26376
rect 15838 26324 15844 26376
rect 15896 26324 15902 26376
rect 15934 26367 15992 26373
rect 15934 26333 15946 26367
rect 15980 26333 15992 26367
rect 15934 26327 15992 26333
rect 10229 26299 10287 26305
rect 10229 26296 10241 26299
rect 8588 26268 9076 26296
rect 4154 26188 4160 26240
rect 4212 26228 4218 26240
rect 4433 26231 4491 26237
rect 4433 26228 4445 26231
rect 4212 26200 4445 26228
rect 4212 26188 4218 26200
rect 4433 26197 4445 26200
rect 4479 26228 4491 26231
rect 4522 26228 4528 26240
rect 4479 26200 4528 26228
rect 4479 26197 4491 26200
rect 4433 26191 4491 26197
rect 4522 26188 4528 26200
rect 4580 26188 4586 26240
rect 5442 26188 5448 26240
rect 5500 26188 5506 26240
rect 6012 26237 6040 26268
rect 5997 26231 6055 26237
rect 5997 26197 6009 26231
rect 6043 26197 6055 26231
rect 9048 26228 9076 26268
rect 9324 26268 10241 26296
rect 9324 26228 9352 26268
rect 10229 26265 10241 26268
rect 10275 26265 10287 26299
rect 10229 26259 10287 26265
rect 10597 26299 10655 26305
rect 10597 26265 10609 26299
rect 10643 26296 10655 26299
rect 10643 26268 11008 26296
rect 10643 26265 10655 26268
rect 10597 26259 10655 26265
rect 9048 26200 9352 26228
rect 10244 26228 10272 26259
rect 10686 26228 10692 26240
rect 10244 26200 10692 26228
rect 5997 26191 6055 26197
rect 10686 26188 10692 26200
rect 10744 26188 10750 26240
rect 10980 26228 11008 26268
rect 13170 26256 13176 26308
rect 13228 26296 13234 26308
rect 13722 26296 13728 26308
rect 13228 26268 13728 26296
rect 13228 26256 13234 26268
rect 13722 26256 13728 26268
rect 13780 26256 13786 26308
rect 15949 26296 15977 26327
rect 16022 26324 16028 26376
rect 16080 26364 16086 26376
rect 16209 26367 16267 26373
rect 16209 26364 16221 26367
rect 16080 26336 16221 26364
rect 16080 26324 16086 26336
rect 16209 26333 16221 26336
rect 16255 26333 16267 26367
rect 16209 26327 16267 26333
rect 15764 26268 15977 26296
rect 15764 26240 15792 26268
rect 16114 26256 16120 26308
rect 16172 26256 16178 26308
rect 16224 26296 16252 26327
rect 16298 26324 16304 26376
rect 16356 26373 16362 26376
rect 16356 26327 16364 26373
rect 16577 26367 16635 26373
rect 16577 26333 16589 26367
rect 16623 26333 16635 26367
rect 16577 26327 16635 26333
rect 16761 26367 16819 26373
rect 16761 26333 16773 26367
rect 16807 26364 16819 26367
rect 17034 26364 17040 26376
rect 16807 26336 17040 26364
rect 16807 26333 16819 26336
rect 16761 26327 16819 26333
rect 16356 26324 16362 26327
rect 16592 26296 16620 26327
rect 17034 26324 17040 26336
rect 17092 26324 17098 26376
rect 17218 26324 17224 26376
rect 17276 26324 17282 26376
rect 17313 26367 17371 26373
rect 17313 26333 17325 26367
rect 17359 26333 17371 26367
rect 17313 26327 17371 26333
rect 16224 26268 16620 26296
rect 17328 26296 17356 26327
rect 17402 26324 17408 26376
rect 17460 26324 17466 26376
rect 17865 26367 17923 26373
rect 17865 26364 17877 26367
rect 17604 26336 17877 26364
rect 17604 26296 17632 26336
rect 17865 26333 17877 26336
rect 17911 26333 17923 26367
rect 17865 26327 17923 26333
rect 17770 26305 17776 26308
rect 17328 26268 17632 26296
rect 17748 26299 17776 26305
rect 17748 26265 17760 26299
rect 17748 26259 17776 26265
rect 17770 26256 17776 26259
rect 17828 26256 17834 26308
rect 17880 26296 17908 26327
rect 17954 26324 17960 26376
rect 18012 26324 18018 26376
rect 18325 26367 18383 26373
rect 18325 26333 18337 26367
rect 18371 26364 18383 26367
rect 18414 26364 18420 26376
rect 18371 26336 18420 26364
rect 18371 26333 18383 26336
rect 18325 26327 18383 26333
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 18506 26324 18512 26376
rect 18564 26324 18570 26376
rect 19260 26364 19288 26395
rect 20254 26392 20260 26404
rect 20312 26432 20318 26444
rect 20622 26432 20628 26444
rect 20312 26404 20628 26432
rect 20312 26392 20318 26404
rect 20622 26392 20628 26404
rect 20680 26432 20686 26444
rect 20916 26441 20944 26472
rect 20901 26435 20959 26441
rect 20680 26404 20852 26432
rect 20680 26392 20686 26404
rect 20824 26373 20852 26404
rect 20901 26401 20913 26435
rect 20947 26401 20959 26435
rect 20901 26395 20959 26401
rect 20073 26367 20131 26373
rect 20073 26364 20085 26367
rect 19260 26336 20085 26364
rect 20073 26333 20085 26336
rect 20119 26364 20131 26367
rect 20809 26367 20867 26373
rect 20119 26336 20760 26364
rect 20119 26333 20131 26336
rect 20073 26327 20131 26333
rect 19886 26296 19892 26308
rect 17880 26268 19892 26296
rect 19886 26256 19892 26268
rect 19944 26296 19950 26308
rect 20441 26299 20499 26305
rect 20441 26296 20453 26299
rect 19944 26268 20453 26296
rect 19944 26256 19950 26268
rect 20441 26265 20453 26268
rect 20487 26265 20499 26299
rect 20441 26259 20499 26265
rect 20530 26256 20536 26308
rect 20588 26305 20594 26308
rect 20588 26299 20616 26305
rect 20604 26265 20616 26299
rect 20732 26296 20760 26336
rect 20809 26333 20821 26367
rect 20855 26333 20867 26367
rect 20809 26327 20867 26333
rect 21085 26367 21143 26373
rect 21085 26333 21097 26367
rect 21131 26333 21143 26367
rect 21085 26327 21143 26333
rect 21100 26296 21128 26327
rect 20732 26268 21128 26296
rect 20588 26259 20616 26265
rect 20588 26256 20594 26259
rect 11514 26228 11520 26240
rect 10980 26200 11520 26228
rect 11514 26188 11520 26200
rect 11572 26188 11578 26240
rect 11974 26188 11980 26240
rect 12032 26228 12038 26240
rect 12161 26231 12219 26237
rect 12161 26228 12173 26231
rect 12032 26200 12173 26228
rect 12032 26188 12038 26200
rect 12161 26197 12173 26200
rect 12207 26197 12219 26231
rect 12161 26191 12219 26197
rect 14550 26188 14556 26240
rect 14608 26228 14614 26240
rect 15657 26231 15715 26237
rect 15657 26228 15669 26231
rect 14608 26200 15669 26228
rect 14608 26188 14614 26200
rect 15657 26197 15669 26200
rect 15703 26197 15715 26231
rect 15657 26191 15715 26197
rect 15746 26188 15752 26240
rect 15804 26188 15810 26240
rect 17586 26188 17592 26240
rect 17644 26188 17650 26240
rect 17862 26188 17868 26240
rect 17920 26228 17926 26240
rect 19429 26231 19487 26237
rect 19429 26228 19441 26231
rect 17920 26200 19441 26228
rect 17920 26188 17926 26200
rect 19429 26197 19441 26200
rect 19475 26197 19487 26231
rect 19429 26191 19487 26197
rect 19518 26188 19524 26240
rect 19576 26228 19582 26240
rect 20349 26231 20407 26237
rect 20349 26228 20361 26231
rect 19576 26200 20361 26228
rect 19576 26188 19582 26200
rect 20349 26197 20361 26200
rect 20395 26197 20407 26231
rect 20349 26191 20407 26197
rect 20717 26231 20775 26237
rect 20717 26197 20729 26231
rect 20763 26228 20775 26231
rect 21192 26228 21220 26540
rect 21468 26404 21956 26432
rect 21468 26373 21496 26404
rect 21453 26367 21511 26373
rect 21453 26333 21465 26367
rect 21499 26333 21511 26367
rect 21453 26327 21511 26333
rect 21542 26324 21548 26376
rect 21600 26364 21606 26376
rect 21928 26373 21956 26404
rect 21637 26367 21695 26373
rect 21637 26364 21649 26367
rect 21600 26336 21649 26364
rect 21600 26324 21606 26336
rect 21637 26333 21649 26336
rect 21683 26364 21695 26367
rect 21729 26367 21787 26373
rect 21729 26364 21741 26367
rect 21683 26336 21741 26364
rect 21683 26333 21695 26336
rect 21637 26327 21695 26333
rect 21729 26333 21741 26336
rect 21775 26333 21787 26367
rect 21729 26327 21787 26333
rect 21913 26367 21971 26373
rect 21913 26333 21925 26367
rect 21959 26364 21971 26367
rect 22278 26364 22284 26376
rect 21959 26336 22284 26364
rect 21959 26333 21971 26336
rect 21913 26327 21971 26333
rect 22278 26324 22284 26336
rect 22336 26324 22342 26376
rect 22480 26373 22508 26540
rect 22554 26528 22560 26580
rect 22612 26568 22618 26580
rect 30101 26571 30159 26577
rect 22612 26540 30052 26568
rect 22612 26528 22618 26540
rect 23382 26460 23388 26512
rect 23440 26500 23446 26512
rect 23753 26503 23811 26509
rect 23440 26472 23704 26500
rect 23440 26460 23446 26472
rect 23106 26392 23112 26444
rect 23164 26392 23170 26444
rect 23566 26392 23572 26444
rect 23624 26392 23630 26444
rect 23676 26432 23704 26472
rect 23753 26469 23765 26503
rect 23799 26500 23811 26503
rect 23842 26500 23848 26512
rect 23799 26472 23848 26500
rect 23799 26469 23811 26472
rect 23753 26463 23811 26469
rect 23842 26460 23848 26472
rect 23900 26500 23906 26512
rect 23937 26503 23995 26509
rect 23937 26500 23949 26503
rect 23900 26472 23949 26500
rect 23900 26460 23906 26472
rect 23937 26469 23949 26472
rect 23983 26469 23995 26503
rect 23937 26463 23995 26469
rect 24044 26472 24624 26500
rect 23676 26404 23980 26432
rect 22465 26367 22523 26373
rect 22465 26333 22477 26367
rect 22511 26333 22523 26367
rect 22465 26327 22523 26333
rect 23293 26367 23351 26373
rect 23293 26333 23305 26367
rect 23339 26364 23351 26367
rect 23382 26364 23388 26376
rect 23339 26336 23388 26364
rect 23339 26333 23351 26336
rect 23293 26327 23351 26333
rect 22480 26296 22508 26327
rect 23382 26324 23388 26336
rect 23440 26324 23446 26376
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26364 23535 26367
rect 23750 26364 23756 26376
rect 23523 26336 23756 26364
rect 23523 26333 23535 26336
rect 23477 26327 23535 26333
rect 23750 26324 23756 26336
rect 23808 26364 23814 26376
rect 23952 26373 23980 26404
rect 23845 26367 23903 26373
rect 23845 26364 23857 26367
rect 23808 26336 23857 26364
rect 23808 26324 23814 26336
rect 23845 26333 23857 26336
rect 23891 26333 23903 26367
rect 23845 26327 23903 26333
rect 23937 26367 23995 26373
rect 23937 26333 23949 26367
rect 23983 26333 23995 26367
rect 23937 26327 23995 26333
rect 24044 26296 24072 26472
rect 24394 26392 24400 26444
rect 24452 26432 24458 26444
rect 24489 26435 24547 26441
rect 24489 26432 24501 26435
rect 24452 26404 24501 26432
rect 24452 26392 24458 26404
rect 24489 26401 24501 26404
rect 24535 26401 24547 26435
rect 24596 26432 24624 26472
rect 27890 26460 27896 26512
rect 27948 26500 27954 26512
rect 28902 26500 28908 26512
rect 27948 26472 28908 26500
rect 27948 26460 27954 26472
rect 28902 26460 28908 26472
rect 28960 26460 28966 26512
rect 30024 26500 30052 26540
rect 30101 26537 30113 26571
rect 30147 26568 30159 26571
rect 30190 26568 30196 26580
rect 30147 26540 30196 26568
rect 30147 26537 30159 26540
rect 30101 26531 30159 26537
rect 30190 26528 30196 26540
rect 30248 26528 30254 26580
rect 31294 26528 31300 26580
rect 31352 26568 31358 26580
rect 31478 26568 31484 26580
rect 31352 26540 31484 26568
rect 31352 26528 31358 26540
rect 31478 26528 31484 26540
rect 31536 26528 31542 26580
rect 32950 26568 32956 26580
rect 31726 26540 32956 26568
rect 31726 26512 31754 26540
rect 32950 26528 32956 26540
rect 33008 26528 33014 26580
rect 33134 26528 33140 26580
rect 33192 26568 33198 26580
rect 33686 26568 33692 26580
rect 33192 26540 33692 26568
rect 33192 26528 33198 26540
rect 33686 26528 33692 26540
rect 33744 26568 33750 26580
rect 33870 26568 33876 26580
rect 33744 26540 33876 26568
rect 33744 26528 33750 26540
rect 33870 26528 33876 26540
rect 33928 26528 33934 26580
rect 34146 26528 34152 26580
rect 34204 26528 34210 26580
rect 34238 26528 34244 26580
rect 34296 26568 34302 26580
rect 35805 26571 35863 26577
rect 35805 26568 35817 26571
rect 34296 26540 35817 26568
rect 34296 26528 34302 26540
rect 35805 26537 35817 26540
rect 35851 26537 35863 26571
rect 40034 26568 40040 26580
rect 35805 26531 35863 26537
rect 35912 26540 40040 26568
rect 31726 26500 31760 26512
rect 30024 26472 31760 26500
rect 31754 26460 31760 26472
rect 31812 26460 31818 26512
rect 31938 26460 31944 26512
rect 31996 26460 32002 26512
rect 32122 26460 32128 26512
rect 32180 26500 32186 26512
rect 35437 26503 35495 26509
rect 32180 26472 34836 26500
rect 32180 26460 32186 26472
rect 29086 26432 29092 26444
rect 24596 26404 29092 26432
rect 24489 26395 24547 26401
rect 29086 26392 29092 26404
rect 29144 26392 29150 26444
rect 29270 26392 29276 26444
rect 29328 26432 29334 26444
rect 30561 26435 30619 26441
rect 30561 26432 30573 26435
rect 29328 26404 30573 26432
rect 29328 26392 29334 26404
rect 30561 26401 30573 26404
rect 30607 26401 30619 26435
rect 30561 26395 30619 26401
rect 30834 26392 30840 26444
rect 30892 26432 30898 26444
rect 32674 26432 32680 26444
rect 30892 26404 31488 26432
rect 30892 26392 30898 26404
rect 31460 26376 31488 26404
rect 31680 26404 32680 26432
rect 24121 26367 24179 26373
rect 24121 26333 24133 26367
rect 24167 26364 24179 26367
rect 24210 26364 24216 26376
rect 24167 26336 24216 26364
rect 24167 26333 24179 26336
rect 24121 26327 24179 26333
rect 24210 26324 24216 26336
rect 24268 26324 24274 26376
rect 26234 26364 26240 26376
rect 25898 26336 26240 26364
rect 26234 26324 26240 26336
rect 26292 26364 26298 26376
rect 29730 26364 29736 26376
rect 26292 26336 29736 26364
rect 26292 26324 26298 26336
rect 29730 26324 29736 26336
rect 29788 26324 29794 26376
rect 30282 26324 30288 26376
rect 30340 26324 30346 26376
rect 30374 26324 30380 26376
rect 30432 26324 30438 26376
rect 30653 26367 30711 26373
rect 30653 26333 30665 26367
rect 30699 26364 30711 26367
rect 30742 26364 30748 26376
rect 30699 26336 30748 26364
rect 30699 26333 30711 26336
rect 30653 26327 30711 26333
rect 30742 26324 30748 26336
rect 30800 26364 30806 26376
rect 30800 26336 30972 26364
rect 30800 26324 30806 26336
rect 22112 26268 22416 26296
rect 22480 26268 24072 26296
rect 24765 26299 24823 26305
rect 22112 26240 22140 26268
rect 20763 26200 21220 26228
rect 20763 26197 20775 26200
rect 20717 26191 20775 26197
rect 21266 26188 21272 26240
rect 21324 26188 21330 26240
rect 21450 26188 21456 26240
rect 21508 26188 21514 26240
rect 22094 26188 22100 26240
rect 22152 26188 22158 26240
rect 22186 26188 22192 26240
rect 22244 26228 22250 26240
rect 22281 26231 22339 26237
rect 22281 26228 22293 26231
rect 22244 26200 22293 26228
rect 22244 26188 22250 26200
rect 22281 26197 22293 26200
rect 22327 26197 22339 26231
rect 22388 26228 22416 26268
rect 24765 26265 24777 26299
rect 24811 26296 24823 26299
rect 24854 26296 24860 26308
rect 24811 26268 24860 26296
rect 24811 26265 24823 26268
rect 24765 26259 24823 26265
rect 24854 26256 24860 26268
rect 24912 26256 24918 26308
rect 22554 26228 22560 26240
rect 22388 26200 22560 26228
rect 22281 26191 22339 26197
rect 22554 26188 22560 26200
rect 22612 26188 22618 26240
rect 23566 26188 23572 26240
rect 23624 26188 23630 26240
rect 25498 26188 25504 26240
rect 25556 26228 25562 26240
rect 26237 26231 26295 26237
rect 26237 26228 26249 26231
rect 25556 26200 26249 26228
rect 25556 26188 25562 26200
rect 26237 26197 26249 26200
rect 26283 26197 26295 26231
rect 30944 26228 30972 26336
rect 31018 26324 31024 26376
rect 31076 26364 31082 26376
rect 31460 26373 31484 26376
rect 31297 26367 31355 26373
rect 31297 26364 31309 26367
rect 31076 26336 31309 26364
rect 31076 26324 31082 26336
rect 31297 26333 31309 26336
rect 31343 26333 31355 26367
rect 31297 26327 31355 26333
rect 31445 26367 31484 26373
rect 31445 26333 31457 26367
rect 31445 26327 31484 26333
rect 31478 26324 31484 26327
rect 31536 26324 31542 26376
rect 31680 26373 31708 26404
rect 32674 26392 32680 26404
rect 32732 26392 32738 26444
rect 33778 26392 33784 26444
rect 33836 26432 33842 26444
rect 34808 26441 34836 26472
rect 35437 26469 35449 26503
rect 35483 26500 35495 26503
rect 35912 26500 35940 26540
rect 40034 26528 40040 26540
rect 40092 26528 40098 26580
rect 35483 26472 35940 26500
rect 35989 26503 36047 26509
rect 35483 26469 35495 26472
rect 35437 26463 35495 26469
rect 35989 26469 36001 26503
rect 36035 26469 36047 26503
rect 35989 26463 36047 26469
rect 36633 26503 36691 26509
rect 36633 26469 36645 26503
rect 36679 26500 36691 26503
rect 37090 26500 37096 26512
rect 36679 26472 37096 26500
rect 36679 26469 36691 26472
rect 36633 26463 36691 26469
rect 34793 26435 34851 26441
rect 33836 26404 33916 26432
rect 33836 26392 33842 26404
rect 31665 26367 31723 26373
rect 31665 26333 31677 26367
rect 31711 26333 31723 26367
rect 31665 26327 31723 26333
rect 31754 26324 31760 26376
rect 31812 26373 31818 26376
rect 31812 26364 31820 26373
rect 31812 26336 31857 26364
rect 31812 26327 31820 26336
rect 31812 26324 31818 26327
rect 33594 26324 33600 26376
rect 33652 26324 33658 26376
rect 33888 26373 33916 26404
rect 34793 26401 34805 26435
rect 34839 26432 34851 26435
rect 35710 26432 35716 26444
rect 34839 26404 35716 26432
rect 34839 26401 34851 26404
rect 34793 26395 34851 26401
rect 35710 26392 35716 26404
rect 35768 26392 35774 26444
rect 36004 26432 36032 26463
rect 37090 26460 37096 26472
rect 37148 26460 37154 26512
rect 37277 26503 37335 26509
rect 37277 26469 37289 26503
rect 37323 26500 37335 26503
rect 39298 26500 39304 26512
rect 37323 26472 39304 26500
rect 37323 26469 37335 26472
rect 37277 26463 37335 26469
rect 39298 26460 39304 26472
rect 39356 26460 39362 26512
rect 38381 26435 38439 26441
rect 38381 26432 38393 26435
rect 36004 26404 37412 26432
rect 33873 26367 33931 26373
rect 33873 26333 33885 26367
rect 33919 26333 33931 26367
rect 33873 26327 33931 26333
rect 33965 26367 34023 26373
rect 33965 26333 33977 26367
rect 34011 26333 34023 26367
rect 33965 26327 34023 26333
rect 31573 26299 31631 26305
rect 31573 26265 31585 26299
rect 31619 26296 31631 26299
rect 32766 26296 32772 26308
rect 31619 26268 32772 26296
rect 31619 26265 31631 26268
rect 31573 26259 31631 26265
rect 32766 26256 32772 26268
rect 32824 26256 32830 26308
rect 33778 26256 33784 26308
rect 33836 26256 33842 26308
rect 31662 26228 31668 26240
rect 30944 26200 31668 26228
rect 26237 26191 26295 26197
rect 31662 26188 31668 26200
rect 31720 26188 31726 26240
rect 33226 26188 33232 26240
rect 33284 26228 33290 26240
rect 33980 26228 34008 26327
rect 34422 26324 34428 26376
rect 34480 26364 34486 26376
rect 34977 26367 35035 26373
rect 34977 26364 34989 26367
rect 34480 26336 34989 26364
rect 34480 26324 34486 26336
rect 34977 26333 34989 26336
rect 35023 26333 35035 26367
rect 34977 26327 35035 26333
rect 34606 26256 34612 26308
rect 34664 26296 34670 26308
rect 34664 26268 34744 26296
rect 34664 26256 34670 26268
rect 33284 26200 34008 26228
rect 34716 26228 34744 26268
rect 34790 26256 34796 26308
rect 34848 26296 34854 26308
rect 35069 26299 35127 26305
rect 35069 26296 35081 26299
rect 34848 26268 35081 26296
rect 34848 26256 34854 26268
rect 35069 26265 35081 26268
rect 35115 26265 35127 26299
rect 35621 26299 35679 26305
rect 35621 26296 35633 26299
rect 35069 26259 35127 26265
rect 35176 26268 35633 26296
rect 35176 26228 35204 26268
rect 35621 26265 35633 26268
rect 35667 26265 35679 26299
rect 35728 26296 35756 26392
rect 36078 26324 36084 26376
rect 36136 26324 36142 26376
rect 36354 26324 36360 26376
rect 36412 26324 36418 26376
rect 36446 26324 36452 26376
rect 36504 26324 36510 26376
rect 36722 26324 36728 26376
rect 36780 26324 36786 26376
rect 36814 26324 36820 26376
rect 36872 26364 36878 26376
rect 36909 26367 36967 26373
rect 36909 26364 36921 26367
rect 36872 26336 36921 26364
rect 36872 26324 36878 26336
rect 36909 26333 36921 26336
rect 36955 26333 36967 26367
rect 36909 26327 36967 26333
rect 36998 26324 37004 26376
rect 37056 26324 37062 26376
rect 37384 26373 37412 26404
rect 37660 26404 38393 26432
rect 37660 26373 37688 26404
rect 38381 26401 38393 26404
rect 38427 26401 38439 26435
rect 38381 26395 38439 26401
rect 40126 26392 40132 26444
rect 40184 26432 40190 26444
rect 40405 26435 40463 26441
rect 40405 26432 40417 26435
rect 40184 26404 40417 26432
rect 40184 26392 40190 26404
rect 40405 26401 40417 26404
rect 40451 26401 40463 26435
rect 40405 26395 40463 26401
rect 40678 26392 40684 26444
rect 40736 26392 40742 26444
rect 41046 26392 41052 26444
rect 41104 26432 41110 26444
rect 42153 26435 42211 26441
rect 42153 26432 42165 26435
rect 41104 26404 42165 26432
rect 41104 26392 41110 26404
rect 42153 26401 42165 26404
rect 42199 26401 42211 26435
rect 42153 26395 42211 26401
rect 37093 26367 37151 26373
rect 37093 26333 37105 26367
rect 37139 26333 37151 26367
rect 37093 26327 37151 26333
rect 37369 26367 37427 26373
rect 37369 26333 37381 26367
rect 37415 26333 37427 26367
rect 37369 26327 37427 26333
rect 37461 26367 37519 26373
rect 37461 26333 37473 26367
rect 37507 26333 37519 26367
rect 37461 26327 37519 26333
rect 37645 26367 37703 26373
rect 37645 26333 37657 26367
rect 37691 26333 37703 26367
rect 37645 26327 37703 26333
rect 37737 26367 37795 26373
rect 37737 26333 37749 26367
rect 37783 26333 37795 26367
rect 37737 26327 37795 26333
rect 35821 26299 35879 26305
rect 35821 26296 35833 26299
rect 35728 26268 35833 26296
rect 35621 26259 35679 26265
rect 35821 26265 35833 26268
rect 35867 26265 35879 26299
rect 35821 26259 35879 26265
rect 36262 26256 36268 26308
rect 36320 26296 36326 26308
rect 36832 26296 36860 26324
rect 36320 26268 36860 26296
rect 36320 26256 36326 26268
rect 34716 26200 35204 26228
rect 33284 26188 33290 26200
rect 36446 26188 36452 26240
rect 36504 26228 36510 26240
rect 37108 26228 37136 26327
rect 37182 26256 37188 26308
rect 37240 26296 37246 26308
rect 37476 26296 37504 26327
rect 37240 26268 37504 26296
rect 37752 26296 37780 26327
rect 38286 26324 38292 26376
rect 38344 26324 38350 26376
rect 39022 26324 39028 26376
rect 39080 26324 39086 26376
rect 37752 26268 38654 26296
rect 37240 26256 37246 26268
rect 36504 26200 37136 26228
rect 36504 26188 36510 26200
rect 37550 26188 37556 26240
rect 37608 26228 37614 26240
rect 38120 26237 38148 26268
rect 37921 26231 37979 26237
rect 37921 26228 37933 26231
rect 37608 26200 37933 26228
rect 37608 26188 37614 26200
rect 37921 26197 37933 26200
rect 37967 26197 37979 26231
rect 37921 26191 37979 26197
rect 38105 26231 38163 26237
rect 38105 26197 38117 26231
rect 38151 26197 38163 26231
rect 38626 26228 38654 26268
rect 39114 26256 39120 26308
rect 39172 26296 39178 26308
rect 39574 26296 39580 26308
rect 39172 26268 39580 26296
rect 39172 26256 39178 26268
rect 39574 26256 39580 26268
rect 39632 26296 39638 26308
rect 39942 26296 39948 26308
rect 39632 26268 39948 26296
rect 39632 26256 39638 26268
rect 39942 26256 39948 26268
rect 40000 26296 40006 26308
rect 40000 26268 41170 26296
rect 40000 26256 40006 26268
rect 39482 26228 39488 26240
rect 38626 26200 39488 26228
rect 38105 26191 38163 26197
rect 39482 26188 39488 26200
rect 39540 26228 39546 26240
rect 40218 26228 40224 26240
rect 39540 26200 40224 26228
rect 39540 26188 39546 26200
rect 40218 26188 40224 26200
rect 40276 26188 40282 26240
rect 1104 26138 42504 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 42504 26138
rect 1104 26064 42504 26086
rect 842 25984 848 26036
rect 900 26024 906 26036
rect 1489 26027 1547 26033
rect 1489 26024 1501 26027
rect 900 25996 1501 26024
rect 900 25984 906 25996
rect 1489 25993 1501 25996
rect 1535 25993 1547 26027
rect 4433 26027 4491 26033
rect 1489 25987 1547 25993
rect 1688 25996 2774 26024
rect 1688 25897 1716 25996
rect 2746 25956 2774 25996
rect 4433 25993 4445 26027
rect 4479 26024 4491 26027
rect 4617 26027 4675 26033
rect 4617 26024 4629 26027
rect 4479 25996 4629 26024
rect 4479 25993 4491 25996
rect 4433 25987 4491 25993
rect 4617 25993 4629 25996
rect 4663 26024 4675 26027
rect 4706 26024 4712 26036
rect 4663 25996 4712 26024
rect 4663 25993 4675 25996
rect 4617 25987 4675 25993
rect 4706 25984 4712 25996
rect 4764 25984 4770 26036
rect 5718 25984 5724 26036
rect 5776 26024 5782 26036
rect 6086 26024 6092 26036
rect 5776 25996 6092 26024
rect 5776 25984 5782 25996
rect 6086 25984 6092 25996
rect 6144 25984 6150 26036
rect 7098 25984 7104 26036
rect 7156 25984 7162 26036
rect 8294 25984 8300 26036
rect 8352 25984 8358 26036
rect 8588 25996 8800 26024
rect 8021 25959 8079 25965
rect 2746 25928 7052 25956
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25857 1731 25891
rect 1673 25851 1731 25857
rect 2682 25848 2688 25900
rect 2740 25848 2746 25900
rect 2774 25848 2780 25900
rect 2832 25888 2838 25900
rect 3145 25891 3203 25897
rect 3145 25888 3157 25891
rect 2832 25860 3157 25888
rect 2832 25848 2838 25860
rect 3145 25857 3157 25860
rect 3191 25857 3203 25891
rect 3145 25851 3203 25857
rect 3697 25891 3755 25897
rect 3697 25857 3709 25891
rect 3743 25888 3755 25891
rect 3786 25888 3792 25900
rect 3743 25860 3792 25888
rect 3743 25857 3755 25860
rect 3697 25851 3755 25857
rect 3160 25752 3188 25851
rect 3786 25848 3792 25860
rect 3844 25848 3850 25900
rect 3881 25891 3939 25897
rect 3881 25857 3893 25891
rect 3927 25857 3939 25891
rect 3881 25851 3939 25857
rect 3513 25823 3571 25829
rect 3513 25789 3525 25823
rect 3559 25820 3571 25823
rect 3602 25820 3608 25832
rect 3559 25792 3608 25820
rect 3559 25789 3571 25792
rect 3513 25783 3571 25789
rect 3602 25780 3608 25792
rect 3660 25780 3666 25832
rect 3896 25752 3924 25851
rect 3970 25848 3976 25900
rect 4028 25888 4034 25900
rect 4341 25891 4399 25897
rect 4341 25888 4353 25891
rect 4028 25860 4353 25888
rect 4028 25848 4034 25860
rect 4341 25857 4353 25860
rect 4387 25857 4399 25891
rect 4341 25851 4399 25857
rect 4430 25848 4436 25900
rect 4488 25888 4494 25900
rect 4525 25891 4583 25897
rect 4525 25888 4537 25891
rect 4488 25860 4537 25888
rect 4488 25848 4494 25860
rect 4525 25857 4537 25860
rect 4571 25888 4583 25891
rect 4706 25888 4712 25900
rect 4571 25860 4712 25888
rect 4571 25857 4583 25860
rect 4525 25851 4583 25857
rect 4706 25848 4712 25860
rect 4764 25848 4770 25900
rect 5077 25891 5135 25897
rect 5077 25857 5089 25891
rect 5123 25888 5135 25891
rect 5350 25888 5356 25900
rect 5123 25860 5356 25888
rect 5123 25857 5135 25860
rect 5077 25851 5135 25857
rect 5350 25848 5356 25860
rect 5408 25848 5414 25900
rect 5810 25848 5816 25900
rect 5868 25848 5874 25900
rect 5905 25891 5963 25897
rect 5905 25857 5917 25891
rect 5951 25888 5963 25891
rect 5994 25888 6000 25900
rect 5951 25860 6000 25888
rect 5951 25857 5963 25860
rect 5905 25851 5963 25857
rect 5994 25848 6000 25860
rect 6052 25848 6058 25900
rect 6086 25848 6092 25900
rect 6144 25848 6150 25900
rect 4249 25823 4307 25829
rect 4249 25789 4261 25823
rect 4295 25820 4307 25823
rect 4614 25820 4620 25832
rect 4295 25792 4620 25820
rect 4295 25789 4307 25792
rect 4249 25783 4307 25789
rect 4614 25780 4620 25792
rect 4672 25780 4678 25832
rect 4798 25780 4804 25832
rect 4856 25820 4862 25832
rect 4985 25823 5043 25829
rect 4985 25820 4997 25823
rect 4856 25792 4997 25820
rect 4856 25780 4862 25792
rect 4985 25789 4997 25792
rect 5031 25789 5043 25823
rect 4985 25783 5043 25789
rect 5261 25823 5319 25829
rect 5261 25789 5273 25823
rect 5307 25820 5319 25823
rect 5445 25823 5503 25829
rect 5445 25820 5457 25823
rect 5307 25792 5457 25820
rect 5307 25789 5319 25792
rect 5261 25783 5319 25789
rect 5445 25789 5457 25792
rect 5491 25789 5503 25823
rect 5445 25783 5503 25789
rect 5537 25823 5595 25829
rect 5537 25789 5549 25823
rect 5583 25820 5595 25823
rect 5583 25792 5948 25820
rect 5583 25789 5595 25792
rect 5537 25783 5595 25789
rect 3160 25724 3924 25752
rect 3896 25684 3924 25724
rect 4522 25712 4528 25764
rect 4580 25752 4586 25764
rect 4816 25752 4844 25780
rect 5920 25764 5948 25792
rect 4580 25724 4844 25752
rect 4580 25712 4586 25724
rect 5626 25712 5632 25764
rect 5684 25712 5690 25764
rect 5902 25712 5908 25764
rect 5960 25712 5966 25764
rect 4706 25684 4712 25696
rect 3896 25656 4712 25684
rect 4706 25644 4712 25656
rect 4764 25644 4770 25696
rect 5718 25644 5724 25696
rect 5776 25644 5782 25696
rect 5997 25687 6055 25693
rect 5997 25653 6009 25687
rect 6043 25684 6055 25687
rect 6362 25684 6368 25696
rect 6043 25656 6368 25684
rect 6043 25653 6055 25656
rect 5997 25647 6055 25653
rect 6362 25644 6368 25656
rect 6420 25644 6426 25696
rect 7024 25684 7052 25928
rect 8021 25925 8033 25959
rect 8067 25956 8079 25959
rect 8588 25956 8616 25996
rect 8067 25928 8616 25956
rect 8067 25925 8079 25928
rect 8021 25919 8079 25925
rect 8662 25916 8668 25968
rect 8720 25916 8726 25968
rect 8772 25956 8800 25996
rect 8938 25984 8944 26036
rect 8996 25984 9002 26036
rect 9401 26027 9459 26033
rect 9401 25993 9413 26027
rect 9447 26024 9459 26027
rect 9582 26024 9588 26036
rect 9447 25996 9588 26024
rect 9447 25993 9459 25996
rect 9401 25987 9459 25993
rect 9416 25956 9444 25987
rect 9582 25984 9588 25996
rect 9640 25984 9646 26036
rect 11514 25984 11520 26036
rect 11572 25984 11578 26036
rect 11977 26027 12035 26033
rect 11977 25993 11989 26027
rect 12023 26024 12035 26027
rect 12158 26024 12164 26036
rect 12023 25996 12164 26024
rect 12023 25993 12035 25996
rect 11977 25987 12035 25993
rect 12158 25984 12164 25996
rect 12216 25984 12222 26036
rect 14734 25984 14740 26036
rect 14792 25984 14798 26036
rect 14918 25984 14924 26036
rect 14976 25984 14982 26036
rect 16025 26027 16083 26033
rect 16025 25993 16037 26027
rect 16071 26024 16083 26027
rect 16298 26024 16304 26036
rect 16071 25996 16304 26024
rect 16071 25993 16083 25996
rect 16025 25987 16083 25993
rect 16298 25984 16304 25996
rect 16356 25984 16362 26036
rect 16482 25984 16488 26036
rect 16540 26024 16546 26036
rect 18230 26024 18236 26036
rect 16540 25996 18236 26024
rect 16540 25984 16546 25996
rect 18230 25984 18236 25996
rect 18288 26024 18294 26036
rect 21818 26024 21824 26036
rect 18288 25996 21128 26024
rect 18288 25984 18294 25996
rect 8772 25928 9444 25956
rect 10226 25916 10232 25968
rect 10284 25956 10290 25968
rect 10514 25959 10572 25965
rect 10514 25956 10526 25959
rect 10284 25928 10526 25956
rect 10284 25916 10290 25928
rect 10514 25925 10526 25928
rect 10560 25925 10572 25959
rect 10514 25919 10572 25925
rect 10686 25916 10692 25968
rect 10744 25956 10750 25968
rect 11885 25959 11943 25965
rect 11885 25956 11897 25959
rect 10744 25928 11897 25956
rect 10744 25916 10750 25928
rect 11885 25925 11897 25928
rect 11931 25925 11943 25959
rect 11885 25919 11943 25925
rect 15562 25916 15568 25968
rect 15620 25956 15626 25968
rect 16390 25956 16396 25968
rect 15620 25928 16396 25956
rect 15620 25916 15626 25928
rect 16390 25916 16396 25928
rect 16448 25916 16454 25968
rect 20438 25956 20444 25968
rect 19996 25928 20444 25956
rect 7282 25848 7288 25900
rect 7340 25848 7346 25900
rect 7374 25848 7380 25900
rect 7432 25848 7438 25900
rect 7650 25848 7656 25900
rect 7708 25848 7714 25900
rect 7745 25891 7803 25897
rect 7745 25857 7757 25891
rect 7791 25857 7803 25891
rect 7745 25851 7803 25857
rect 7760 25820 7788 25851
rect 7926 25848 7932 25900
rect 7984 25848 7990 25900
rect 8113 25891 8171 25897
rect 8113 25857 8125 25891
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 8018 25820 8024 25832
rect 7760 25792 8024 25820
rect 8018 25780 8024 25792
rect 8076 25780 8082 25832
rect 8128 25820 8156 25851
rect 8386 25848 8392 25900
rect 8444 25848 8450 25900
rect 8570 25848 8576 25900
rect 8628 25848 8634 25900
rect 8757 25891 8815 25897
rect 8757 25857 8769 25891
rect 8803 25888 8815 25891
rect 8846 25888 8852 25900
rect 8803 25860 8852 25888
rect 8803 25857 8815 25860
rect 8757 25851 8815 25857
rect 8772 25820 8800 25851
rect 8846 25848 8852 25860
rect 8904 25848 8910 25900
rect 10778 25848 10784 25900
rect 10836 25848 10842 25900
rect 12434 25848 12440 25900
rect 12492 25888 12498 25900
rect 12529 25891 12587 25897
rect 12529 25888 12541 25891
rect 12492 25860 12541 25888
rect 12492 25848 12498 25860
rect 12529 25857 12541 25860
rect 12575 25857 12587 25891
rect 12529 25851 12587 25857
rect 12713 25891 12771 25897
rect 12713 25857 12725 25891
rect 12759 25888 12771 25891
rect 12802 25888 12808 25900
rect 12759 25860 12808 25888
rect 12759 25857 12771 25860
rect 12713 25851 12771 25857
rect 12802 25848 12808 25860
rect 12860 25848 12866 25900
rect 14366 25848 14372 25900
rect 14424 25848 14430 25900
rect 14550 25897 14556 25900
rect 14523 25891 14556 25897
rect 14523 25857 14535 25891
rect 14523 25851 14556 25857
rect 14550 25848 14556 25851
rect 14608 25848 14614 25900
rect 14826 25848 14832 25900
rect 14884 25848 14890 25900
rect 15010 25848 15016 25900
rect 15068 25848 15074 25900
rect 15105 25891 15163 25897
rect 15105 25857 15117 25891
rect 15151 25857 15163 25891
rect 15105 25851 15163 25857
rect 15197 25891 15255 25897
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 15286 25888 15292 25900
rect 15243 25860 15292 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 8128 25792 8800 25820
rect 12158 25780 12164 25832
rect 12216 25780 12222 25832
rect 14918 25780 14924 25832
rect 14976 25820 14982 25832
rect 15120 25820 15148 25851
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 15381 25891 15439 25897
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 14976 25792 15148 25820
rect 15396 25820 15424 25851
rect 15470 25848 15476 25900
rect 15528 25848 15534 25900
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25857 16175 25891
rect 16117 25851 16175 25857
rect 16945 25891 17003 25897
rect 16945 25857 16957 25891
rect 16991 25888 17003 25891
rect 17954 25888 17960 25900
rect 16991 25860 17960 25888
rect 16991 25857 17003 25860
rect 16945 25851 17003 25857
rect 16022 25820 16028 25832
rect 15396 25792 16028 25820
rect 14976 25780 14982 25792
rect 16022 25780 16028 25792
rect 16080 25780 16086 25832
rect 16132 25820 16160 25851
rect 17954 25848 17960 25860
rect 18012 25888 18018 25900
rect 19426 25888 19432 25900
rect 18012 25860 19432 25888
rect 18012 25848 18018 25860
rect 19426 25848 19432 25860
rect 19484 25888 19490 25900
rect 19996 25897 20024 25928
rect 20438 25916 20444 25928
rect 20496 25916 20502 25968
rect 21100 25956 21128 25996
rect 21284 25996 21824 26024
rect 21174 25956 21180 25968
rect 21100 25928 21180 25956
rect 19981 25891 20039 25897
rect 19981 25888 19993 25891
rect 19484 25860 19993 25888
rect 19484 25848 19490 25860
rect 19981 25857 19993 25860
rect 20027 25857 20039 25891
rect 19981 25851 20039 25857
rect 20073 25891 20131 25897
rect 20073 25857 20085 25891
rect 20119 25857 20131 25891
rect 20073 25851 20131 25857
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 16132 25792 16681 25820
rect 16669 25789 16681 25792
rect 16715 25820 16727 25823
rect 17034 25820 17040 25832
rect 16715 25792 17040 25820
rect 16715 25789 16727 25792
rect 16669 25783 16727 25789
rect 17034 25780 17040 25792
rect 17092 25780 17098 25832
rect 19518 25780 19524 25832
rect 19576 25820 19582 25832
rect 20088 25820 20116 25851
rect 20162 25848 20168 25900
rect 20220 25888 20226 25900
rect 20349 25891 20407 25897
rect 20349 25888 20361 25891
rect 20220 25860 20361 25888
rect 20220 25848 20226 25860
rect 20349 25857 20361 25860
rect 20395 25888 20407 25891
rect 20530 25888 20536 25900
rect 20395 25860 20536 25888
rect 20395 25857 20407 25860
rect 20349 25851 20407 25857
rect 20530 25848 20536 25860
rect 20588 25848 20594 25900
rect 21100 25897 21128 25928
rect 21174 25916 21180 25928
rect 21232 25916 21238 25968
rect 21284 25897 21312 25996
rect 21818 25984 21824 25996
rect 21876 25984 21882 26036
rect 22281 26027 22339 26033
rect 22281 25993 22293 26027
rect 22327 26024 22339 26027
rect 23569 26027 23627 26033
rect 22327 25996 23336 26024
rect 22327 25993 22339 25996
rect 22281 25987 22339 25993
rect 21450 25916 21456 25968
rect 21508 25916 21514 25968
rect 21637 25959 21695 25965
rect 21637 25925 21649 25959
rect 21683 25956 21695 25959
rect 22094 25956 22100 25968
rect 21683 25928 22100 25956
rect 21683 25925 21695 25928
rect 21637 25919 21695 25925
rect 22094 25916 22100 25928
rect 22152 25916 22158 25968
rect 22373 25959 22431 25965
rect 22373 25956 22385 25959
rect 22296 25928 22385 25956
rect 21085 25891 21143 25897
rect 21085 25857 21097 25891
rect 21131 25857 21143 25891
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 21085 25851 21143 25857
rect 21192 25860 21281 25888
rect 19576 25792 20116 25820
rect 19576 25780 19582 25792
rect 20254 25780 20260 25832
rect 20312 25780 20318 25832
rect 7098 25712 7104 25764
rect 7156 25752 7162 25764
rect 7561 25755 7619 25761
rect 7561 25752 7573 25755
rect 7156 25724 7573 25752
rect 7156 25712 7162 25724
rect 7561 25721 7573 25724
rect 7607 25721 7619 25755
rect 8036 25752 8064 25780
rect 8570 25752 8576 25764
rect 8036 25724 8576 25752
rect 7561 25715 7619 25721
rect 8570 25712 8576 25724
rect 8628 25712 8634 25764
rect 15102 25712 15108 25764
rect 15160 25752 15166 25764
rect 16761 25755 16819 25761
rect 16761 25752 16773 25755
rect 15160 25724 16773 25752
rect 15160 25712 15166 25724
rect 16761 25721 16773 25724
rect 16807 25721 16819 25755
rect 16761 25715 16819 25721
rect 16853 25755 16911 25761
rect 16853 25721 16865 25755
rect 16899 25752 16911 25755
rect 17862 25752 17868 25764
rect 16899 25724 17868 25752
rect 16899 25721 16911 25724
rect 16853 25715 16911 25721
rect 11974 25684 11980 25696
rect 7024 25656 11980 25684
rect 11974 25644 11980 25656
rect 12032 25644 12038 25696
rect 12529 25687 12587 25693
rect 12529 25653 12541 25687
rect 12575 25684 12587 25687
rect 12710 25684 12716 25696
rect 12575 25656 12716 25684
rect 12575 25653 12587 25656
rect 12529 25647 12587 25653
rect 12710 25644 12716 25656
rect 12768 25644 12774 25696
rect 14826 25644 14832 25696
rect 14884 25684 14890 25696
rect 15470 25684 15476 25696
rect 14884 25656 15476 25684
rect 14884 25644 14890 25656
rect 15470 25644 15476 25656
rect 15528 25644 15534 25696
rect 15657 25687 15715 25693
rect 15657 25653 15669 25687
rect 15703 25684 15715 25687
rect 15838 25684 15844 25696
rect 15703 25656 15844 25684
rect 15703 25653 15715 25656
rect 15657 25647 15715 25653
rect 15838 25644 15844 25656
rect 15896 25644 15902 25696
rect 16390 25644 16396 25696
rect 16448 25684 16454 25696
rect 16868 25684 16896 25715
rect 17862 25712 17868 25724
rect 17920 25712 17926 25764
rect 18322 25712 18328 25764
rect 18380 25752 18386 25764
rect 21192 25752 21220 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 21358 25848 21364 25900
rect 21416 25848 21422 25900
rect 21468 25888 21496 25916
rect 22002 25888 22008 25900
rect 21468 25860 22008 25888
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 21376 25820 21404 25848
rect 22296 25820 22324 25928
rect 22373 25925 22385 25928
rect 22419 25925 22431 25959
rect 22373 25919 22431 25925
rect 22649 25959 22707 25965
rect 22649 25925 22661 25959
rect 22695 25956 22707 25959
rect 22695 25928 22968 25956
rect 22695 25925 22707 25928
rect 22649 25919 22707 25925
rect 22554 25897 22560 25900
rect 22458 25891 22516 25897
rect 22458 25857 22470 25891
rect 22504 25888 22516 25891
rect 22547 25891 22560 25897
rect 22547 25888 22559 25891
rect 22504 25860 22559 25888
rect 22504 25857 22516 25860
rect 22458 25851 22516 25857
rect 22547 25857 22559 25860
rect 22547 25851 22560 25857
rect 22554 25848 22560 25851
rect 22612 25848 22618 25900
rect 22833 25891 22891 25897
rect 22833 25888 22845 25891
rect 22664 25860 22845 25888
rect 22664 25820 22692 25860
rect 22833 25857 22845 25860
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 21376 25792 22692 25820
rect 18380 25724 21220 25752
rect 21269 25755 21327 25761
rect 18380 25712 18386 25724
rect 21269 25721 21281 25755
rect 21315 25752 21327 25755
rect 22278 25752 22284 25764
rect 21315 25724 22284 25752
rect 21315 25721 21327 25724
rect 21269 25715 21327 25721
rect 22278 25712 22284 25724
rect 22336 25712 22342 25764
rect 16448 25656 16896 25684
rect 21545 25687 21603 25693
rect 16448 25644 16454 25656
rect 21545 25653 21557 25687
rect 21591 25684 21603 25687
rect 21634 25684 21640 25696
rect 21591 25656 21640 25684
rect 21591 25653 21603 25656
rect 21545 25647 21603 25653
rect 21634 25644 21640 25656
rect 21692 25644 21698 25696
rect 22002 25644 22008 25696
rect 22060 25684 22066 25696
rect 22940 25684 22968 25928
rect 23308 25897 23336 25996
rect 23569 25993 23581 26027
rect 23615 25993 23627 26027
rect 23569 25987 23627 25993
rect 23584 25956 23612 25987
rect 24854 25984 24860 26036
rect 24912 26024 24918 26036
rect 24949 26027 25007 26033
rect 24949 26024 24961 26027
rect 24912 25996 24961 26024
rect 24912 25984 24918 25996
rect 24949 25993 24961 25996
rect 24995 25993 25007 26027
rect 24949 25987 25007 25993
rect 29365 26027 29423 26033
rect 29365 25993 29377 26027
rect 29411 26024 29423 26027
rect 29454 26024 29460 26036
rect 29411 25996 29460 26024
rect 29411 25993 29423 25996
rect 29365 25987 29423 25993
rect 29454 25984 29460 25996
rect 29512 26024 29518 26036
rect 29638 26024 29644 26036
rect 29512 25996 29644 26024
rect 29512 25984 29518 25996
rect 29638 25984 29644 25996
rect 29696 25984 29702 26036
rect 31662 25984 31668 26036
rect 31720 26024 31726 26036
rect 32401 26027 32459 26033
rect 32401 26024 32413 26027
rect 31720 25996 32413 26024
rect 31720 25984 31726 25996
rect 32401 25993 32413 25996
rect 32447 25993 32459 26027
rect 32401 25987 32459 25993
rect 32493 26027 32551 26033
rect 32493 25993 32505 26027
rect 32539 26024 32551 26027
rect 32674 26024 32680 26036
rect 32539 25996 32680 26024
rect 32539 25993 32551 25996
rect 32493 25987 32551 25993
rect 32674 25984 32680 25996
rect 32732 25984 32738 26036
rect 32766 25984 32772 26036
rect 32824 26024 32830 26036
rect 33778 26024 33784 26036
rect 32824 25996 33784 26024
rect 32824 25984 32830 25996
rect 33778 25984 33784 25996
rect 33836 26024 33842 26036
rect 36262 26024 36268 26036
rect 33836 25996 36268 26024
rect 33836 25984 33842 25996
rect 36262 25984 36268 25996
rect 36320 25984 36326 26036
rect 39022 25984 39028 26036
rect 39080 25984 39086 26036
rect 39853 26027 39911 26033
rect 39853 26024 39865 26027
rect 39500 25996 39865 26024
rect 25222 25956 25228 25968
rect 23584 25928 25228 25956
rect 25222 25916 25228 25928
rect 25280 25916 25286 25968
rect 31386 25956 31392 25968
rect 29118 25942 31392 25956
rect 29104 25928 31392 25942
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25857 23351 25891
rect 23293 25851 23351 25857
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25888 23535 25891
rect 23842 25888 23848 25900
rect 23523 25860 23848 25888
rect 23523 25857 23535 25860
rect 23477 25851 23535 25857
rect 23308 25820 23336 25851
rect 23842 25848 23848 25860
rect 23900 25848 23906 25900
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 25133 25891 25191 25897
rect 25133 25888 25145 25891
rect 25004 25860 25145 25888
rect 25004 25848 25010 25860
rect 25133 25857 25145 25860
rect 25179 25857 25191 25891
rect 25133 25851 25191 25857
rect 25409 25891 25467 25897
rect 25409 25857 25421 25891
rect 25455 25888 25467 25891
rect 25498 25888 25504 25900
rect 25455 25860 25504 25888
rect 25455 25857 25467 25860
rect 25409 25851 25467 25857
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 23658 25820 23664 25832
rect 23308 25792 23664 25820
rect 23658 25780 23664 25792
rect 23716 25820 23722 25832
rect 23937 25823 23995 25829
rect 23937 25820 23949 25823
rect 23716 25792 23949 25820
rect 23716 25780 23722 25792
rect 23937 25789 23949 25792
rect 23983 25789 23995 25823
rect 23937 25783 23995 25789
rect 27614 25780 27620 25832
rect 27672 25780 27678 25832
rect 27890 25780 27896 25832
rect 27948 25780 27954 25832
rect 28442 25780 28448 25832
rect 28500 25820 28506 25832
rect 29104 25820 29132 25928
rect 31386 25916 31392 25928
rect 31444 25916 31450 25968
rect 37550 25916 37556 25968
rect 37608 25916 37614 25968
rect 39114 25956 39120 25968
rect 38778 25928 39120 25956
rect 39114 25916 39120 25928
rect 39172 25916 39178 25968
rect 39298 25916 39304 25968
rect 39356 25916 39362 25968
rect 39500 25965 39528 25996
rect 39853 25993 39865 25996
rect 39899 25993 39911 26027
rect 39853 25987 39911 25993
rect 40034 25984 40040 26036
rect 40092 26024 40098 26036
rect 40310 26024 40316 26036
rect 40092 25996 40316 26024
rect 40092 25984 40098 25996
rect 40310 25984 40316 25996
rect 40368 25984 40374 26036
rect 40497 26027 40555 26033
rect 40497 25993 40509 26027
rect 40543 26024 40555 26027
rect 40586 26024 40592 26036
rect 40543 25996 40592 26024
rect 40543 25993 40555 25996
rect 40497 25987 40555 25993
rect 40586 25984 40592 25996
rect 40644 25984 40650 26036
rect 42058 25984 42064 26036
rect 42116 25984 42122 26036
rect 39485 25959 39543 25965
rect 39485 25925 39497 25959
rect 39531 25925 39543 25959
rect 40770 25956 40776 25968
rect 40828 25965 40834 25968
rect 39485 25919 39543 25925
rect 39960 25928 40632 25956
rect 40735 25928 40776 25956
rect 39206 25848 39212 25900
rect 39264 25888 39270 25900
rect 39960 25888 39988 25928
rect 39264 25860 39988 25888
rect 39264 25848 39270 25860
rect 40034 25848 40040 25900
rect 40092 25848 40098 25900
rect 40126 25848 40132 25900
rect 40184 25848 40190 25900
rect 40218 25848 40224 25900
rect 40276 25848 40282 25900
rect 40405 25891 40463 25897
rect 40405 25857 40417 25891
rect 40451 25888 40463 25891
rect 40494 25888 40500 25900
rect 40451 25860 40500 25888
rect 40451 25857 40463 25860
rect 40405 25851 40463 25857
rect 40494 25848 40500 25860
rect 40552 25848 40558 25900
rect 40604 25888 40632 25928
rect 40770 25916 40776 25928
rect 40828 25919 40835 25965
rect 40828 25916 40834 25919
rect 40681 25891 40739 25897
rect 40681 25888 40693 25891
rect 40604 25860 40693 25888
rect 40681 25857 40693 25860
rect 40727 25857 40739 25891
rect 40681 25851 40739 25857
rect 40862 25848 40868 25900
rect 40920 25848 40926 25900
rect 41046 25848 41052 25900
rect 41104 25848 41110 25900
rect 41874 25848 41880 25900
rect 41932 25848 41938 25900
rect 28500 25792 29132 25820
rect 28500 25780 28506 25792
rect 32122 25780 32128 25832
rect 32180 25820 32186 25832
rect 32217 25823 32275 25829
rect 32217 25820 32229 25823
rect 32180 25792 32229 25820
rect 32180 25780 32186 25792
rect 32217 25789 32229 25792
rect 32263 25789 32275 25823
rect 32217 25783 32275 25789
rect 37274 25780 37280 25832
rect 37332 25780 37338 25832
rect 39390 25780 39396 25832
rect 39448 25820 39454 25832
rect 40144 25820 40172 25848
rect 40770 25820 40776 25832
rect 39448 25792 40776 25820
rect 39448 25780 39454 25792
rect 40770 25780 40776 25792
rect 40828 25780 40834 25832
rect 23290 25712 23296 25764
rect 23348 25752 23354 25764
rect 24213 25755 24271 25761
rect 24213 25752 24225 25755
rect 23348 25724 24225 25752
rect 23348 25712 23354 25724
rect 24213 25721 24225 25724
rect 24259 25721 24271 25755
rect 24213 25715 24271 25721
rect 38580 25724 39252 25752
rect 22060 25656 22968 25684
rect 22060 25644 22066 25656
rect 23014 25644 23020 25696
rect 23072 25644 23078 25696
rect 23750 25644 23756 25696
rect 23808 25684 23814 25696
rect 23845 25687 23903 25693
rect 23845 25684 23857 25687
rect 23808 25656 23857 25684
rect 23808 25644 23814 25656
rect 23845 25653 23857 25656
rect 23891 25653 23903 25687
rect 23845 25647 23903 25653
rect 25038 25644 25044 25696
rect 25096 25684 25102 25696
rect 25317 25687 25375 25693
rect 25317 25684 25329 25687
rect 25096 25656 25329 25684
rect 25096 25644 25102 25656
rect 25317 25653 25329 25656
rect 25363 25684 25375 25687
rect 28902 25684 28908 25696
rect 25363 25656 28908 25684
rect 25363 25653 25375 25656
rect 25317 25647 25375 25653
rect 28902 25644 28908 25656
rect 28960 25684 28966 25696
rect 30558 25684 30564 25696
rect 28960 25656 30564 25684
rect 28960 25644 28966 25656
rect 30558 25644 30564 25656
rect 30616 25644 30622 25696
rect 32858 25644 32864 25696
rect 32916 25644 32922 25696
rect 33778 25644 33784 25696
rect 33836 25684 33842 25696
rect 38580 25684 38608 25724
rect 33836 25656 38608 25684
rect 33836 25644 33842 25656
rect 39114 25644 39120 25696
rect 39172 25644 39178 25696
rect 39224 25684 39252 25724
rect 40218 25712 40224 25764
rect 40276 25752 40282 25764
rect 40862 25752 40868 25764
rect 40276 25724 40868 25752
rect 40276 25712 40282 25724
rect 40862 25712 40868 25724
rect 40920 25712 40926 25764
rect 40954 25684 40960 25696
rect 39224 25656 40960 25684
rect 40954 25644 40960 25656
rect 41012 25644 41018 25696
rect 1104 25594 42504 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 42504 25594
rect 1104 25520 42504 25542
rect 14737 25483 14795 25489
rect 14737 25449 14749 25483
rect 14783 25480 14795 25483
rect 14826 25480 14832 25492
rect 14783 25452 14832 25480
rect 14783 25449 14795 25452
rect 14737 25443 14795 25449
rect 14826 25440 14832 25452
rect 14884 25440 14890 25492
rect 14918 25440 14924 25492
rect 14976 25480 14982 25492
rect 15381 25483 15439 25489
rect 15381 25480 15393 25483
rect 14976 25452 15393 25480
rect 14976 25440 14982 25452
rect 15381 25449 15393 25452
rect 15427 25480 15439 25483
rect 17313 25483 17371 25489
rect 15427 25452 16896 25480
rect 15427 25449 15439 25452
rect 15381 25443 15439 25449
rect 4430 25372 4436 25424
rect 4488 25412 4494 25424
rect 5442 25412 5448 25424
rect 4488 25384 5448 25412
rect 4488 25372 4494 25384
rect 5442 25372 5448 25384
rect 5500 25412 5506 25424
rect 5810 25412 5816 25424
rect 5500 25384 5816 25412
rect 5500 25372 5506 25384
rect 5810 25372 5816 25384
rect 5868 25412 5874 25424
rect 16868 25412 16896 25452
rect 17313 25449 17325 25483
rect 17359 25480 17371 25483
rect 17770 25480 17776 25492
rect 17359 25452 17776 25480
rect 17359 25449 17371 25452
rect 17313 25443 17371 25449
rect 17770 25440 17776 25452
rect 17828 25440 17834 25492
rect 18138 25440 18144 25492
rect 18196 25440 18202 25492
rect 21174 25440 21180 25492
rect 21232 25480 21238 25492
rect 22094 25480 22100 25492
rect 21232 25452 22100 25480
rect 21232 25440 21238 25452
rect 22094 25440 22100 25452
rect 22152 25480 22158 25492
rect 23382 25480 23388 25492
rect 22152 25452 23388 25480
rect 22152 25440 22158 25452
rect 23382 25440 23388 25452
rect 23440 25440 23446 25492
rect 24946 25440 24952 25492
rect 25004 25440 25010 25492
rect 26234 25480 26240 25492
rect 25148 25452 26240 25480
rect 20806 25412 20812 25424
rect 5868 25384 15516 25412
rect 16868 25384 20812 25412
rect 5868 25372 5874 25384
rect 2866 25304 2872 25356
rect 2924 25304 2930 25356
rect 3145 25347 3203 25353
rect 3145 25313 3157 25347
rect 3191 25344 3203 25347
rect 3510 25344 3516 25356
rect 3191 25316 3516 25344
rect 3191 25313 3203 25316
rect 3145 25307 3203 25313
rect 3510 25304 3516 25316
rect 3568 25344 3574 25356
rect 6086 25344 6092 25356
rect 3568 25316 6092 25344
rect 3568 25304 3574 25316
rect 6086 25304 6092 25316
rect 6144 25304 6150 25356
rect 15102 25304 15108 25356
rect 15160 25304 15166 25356
rect 4522 25236 4528 25288
rect 4580 25276 4586 25288
rect 4985 25279 5043 25285
rect 4985 25276 4997 25279
rect 4580 25248 4997 25276
rect 4580 25236 4586 25248
rect 4985 25245 4997 25248
rect 5031 25245 5043 25279
rect 4985 25239 5043 25245
rect 7558 25236 7564 25288
rect 7616 25276 7622 25288
rect 7653 25279 7711 25285
rect 7653 25276 7665 25279
rect 7616 25248 7665 25276
rect 7616 25236 7622 25248
rect 7653 25245 7665 25248
rect 7699 25245 7711 25279
rect 7653 25239 7711 25245
rect 2958 25208 2964 25220
rect 2438 25180 2964 25208
rect 2958 25168 2964 25180
rect 3016 25168 3022 25220
rect 7668 25208 7696 25239
rect 7742 25236 7748 25288
rect 7800 25276 7806 25288
rect 7837 25279 7895 25285
rect 7837 25276 7849 25279
rect 7800 25248 7849 25276
rect 7800 25236 7806 25248
rect 7837 25245 7849 25248
rect 7883 25245 7895 25279
rect 7837 25239 7895 25245
rect 13446 25236 13452 25288
rect 13504 25236 13510 25288
rect 15010 25236 15016 25288
rect 15068 25236 15074 25288
rect 15488 25285 15516 25384
rect 20806 25372 20812 25384
rect 20864 25372 20870 25424
rect 15838 25304 15844 25356
rect 15896 25304 15902 25356
rect 18322 25344 18328 25356
rect 18064 25316 18328 25344
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 8294 25208 8300 25220
rect 7668 25180 8300 25208
rect 8294 25168 8300 25180
rect 8352 25168 8358 25220
rect 11422 25168 11428 25220
rect 11480 25208 11486 25220
rect 14366 25208 14372 25220
rect 11480 25180 14372 25208
rect 11480 25168 11486 25180
rect 14366 25168 14372 25180
rect 14424 25168 14430 25220
rect 14550 25168 14556 25220
rect 14608 25168 14614 25220
rect 1394 25100 1400 25152
rect 1452 25100 1458 25152
rect 5169 25143 5227 25149
rect 5169 25109 5181 25143
rect 5215 25140 5227 25143
rect 5718 25140 5724 25152
rect 5215 25112 5724 25140
rect 5215 25109 5227 25112
rect 5169 25103 5227 25109
rect 5718 25100 5724 25112
rect 5776 25140 5782 25152
rect 6454 25140 6460 25152
rect 5776 25112 6460 25140
rect 5776 25100 5782 25112
rect 6454 25100 6460 25112
rect 6512 25100 6518 25152
rect 7834 25100 7840 25152
rect 7892 25100 7898 25152
rect 13357 25143 13415 25149
rect 13357 25109 13369 25143
rect 13403 25140 13415 25143
rect 13630 25140 13636 25152
rect 13403 25112 13636 25140
rect 13403 25109 13415 25112
rect 13357 25103 13415 25109
rect 13630 25100 13636 25112
rect 13688 25100 13694 25152
rect 14829 25143 14887 25149
rect 14829 25109 14841 25143
rect 14875 25140 14887 25143
rect 14918 25140 14924 25152
rect 14875 25112 14924 25140
rect 14875 25109 14887 25112
rect 14829 25103 14887 25109
rect 14918 25100 14924 25112
rect 14976 25100 14982 25152
rect 15488 25140 15516 25239
rect 15562 25236 15568 25288
rect 15620 25236 15626 25288
rect 18064 25285 18092 25316
rect 18322 25304 18328 25316
rect 18380 25304 18386 25356
rect 23014 25344 23020 25356
rect 21744 25316 23020 25344
rect 18049 25279 18107 25285
rect 18049 25245 18061 25279
rect 18095 25245 18107 25279
rect 18049 25239 18107 25245
rect 18230 25236 18236 25288
rect 18288 25236 18294 25288
rect 20898 25236 20904 25288
rect 20956 25276 20962 25288
rect 21082 25276 21088 25288
rect 20956 25248 21088 25276
rect 20956 25236 20962 25248
rect 21082 25236 21088 25248
rect 21140 25276 21146 25288
rect 21269 25279 21327 25285
rect 21269 25276 21281 25279
rect 21140 25248 21281 25276
rect 21140 25236 21146 25248
rect 21269 25245 21281 25248
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 21634 25236 21640 25288
rect 21692 25236 21698 25288
rect 21744 25285 21772 25316
rect 23014 25304 23020 25316
rect 23072 25304 23078 25356
rect 23566 25344 23572 25356
rect 23216 25316 23572 25344
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25245 21787 25279
rect 22094 25276 22100 25288
rect 21729 25239 21787 25245
rect 21836 25248 22100 25276
rect 17126 25208 17132 25220
rect 17066 25180 17132 25208
rect 17126 25168 17132 25180
rect 17184 25208 17190 25220
rect 17497 25211 17555 25217
rect 17497 25208 17509 25211
rect 17184 25180 17509 25208
rect 17184 25168 17190 25180
rect 17497 25177 17509 25180
rect 17543 25177 17555 25211
rect 17497 25171 17555 25177
rect 17862 25168 17868 25220
rect 17920 25168 17926 25220
rect 17954 25168 17960 25220
rect 18012 25208 18018 25220
rect 18248 25208 18276 25236
rect 18012 25180 18276 25208
rect 21407 25211 21465 25217
rect 18012 25168 18018 25180
rect 21407 25177 21419 25211
rect 21453 25177 21465 25211
rect 21407 25171 21465 25177
rect 21545 25211 21603 25217
rect 21545 25177 21557 25211
rect 21591 25208 21603 25211
rect 21836 25208 21864 25248
rect 22094 25236 22100 25248
rect 22152 25236 22158 25288
rect 22278 25236 22284 25288
rect 22336 25276 22342 25288
rect 23216 25285 23244 25316
rect 23566 25304 23572 25316
rect 23624 25304 23630 25356
rect 23201 25279 23259 25285
rect 22336 25248 23152 25276
rect 22336 25236 22342 25248
rect 21591 25180 21864 25208
rect 21913 25211 21971 25217
rect 21591 25177 21603 25180
rect 21545 25171 21603 25177
rect 21913 25177 21925 25211
rect 21959 25208 21971 25211
rect 21959 25180 22324 25208
rect 21959 25177 21971 25180
rect 21913 25171 21971 25177
rect 16758 25140 16764 25152
rect 15488 25112 16764 25140
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 18414 25100 18420 25152
rect 18472 25100 18478 25152
rect 20438 25100 20444 25152
rect 20496 25140 20502 25152
rect 21422 25140 21450 25171
rect 22296 25152 22324 25180
rect 22094 25140 22100 25152
rect 20496 25112 22100 25140
rect 20496 25100 20502 25112
rect 22094 25100 22100 25112
rect 22152 25100 22158 25152
rect 22278 25100 22284 25152
rect 22336 25100 22342 25152
rect 23014 25100 23020 25152
rect 23072 25100 23078 25152
rect 23124 25140 23152 25248
rect 23201 25245 23213 25279
rect 23247 25245 23259 25279
rect 23201 25239 23259 25245
rect 23290 25236 23296 25288
rect 23348 25236 23354 25288
rect 23658 25236 23664 25288
rect 23716 25276 23722 25288
rect 23934 25276 23940 25288
rect 23716 25248 23940 25276
rect 23716 25236 23722 25248
rect 23934 25236 23940 25248
rect 23992 25236 23998 25288
rect 24578 25236 24584 25288
rect 24636 25276 24642 25288
rect 25148 25285 25176 25452
rect 26234 25440 26240 25452
rect 26292 25440 26298 25492
rect 27890 25440 27896 25492
rect 27948 25480 27954 25492
rect 28169 25483 28227 25489
rect 28169 25480 28181 25483
rect 27948 25452 28181 25480
rect 27948 25440 27954 25452
rect 28169 25449 28181 25452
rect 28215 25449 28227 25483
rect 40313 25483 40371 25489
rect 40313 25480 40325 25483
rect 28169 25443 28227 25449
rect 29196 25452 40325 25480
rect 25498 25372 25504 25424
rect 25556 25372 25562 25424
rect 26694 25372 26700 25424
rect 26752 25412 26758 25424
rect 29196 25412 29224 25452
rect 40313 25449 40325 25452
rect 40359 25449 40371 25483
rect 40313 25443 40371 25449
rect 26752 25384 29224 25412
rect 26752 25372 26758 25384
rect 29270 25372 29276 25424
rect 29328 25412 29334 25424
rect 30193 25415 30251 25421
rect 30193 25412 30205 25415
rect 29328 25384 30205 25412
rect 29328 25372 29334 25384
rect 30193 25381 30205 25384
rect 30239 25381 30251 25415
rect 30193 25375 30251 25381
rect 25516 25344 25544 25372
rect 28813 25347 28871 25353
rect 25516 25316 25820 25344
rect 25133 25279 25191 25285
rect 25133 25276 25145 25279
rect 24636 25248 25145 25276
rect 24636 25236 24642 25248
rect 25133 25245 25145 25248
rect 25179 25245 25191 25279
rect 25133 25239 25191 25245
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25276 25283 25279
rect 25406 25276 25412 25288
rect 25271 25248 25412 25276
rect 25271 25245 25283 25248
rect 25225 25239 25283 25245
rect 25406 25236 25412 25248
rect 25464 25236 25470 25288
rect 25792 25285 25820 25316
rect 28813 25313 28825 25347
rect 28859 25344 28871 25347
rect 28902 25344 28908 25356
rect 28859 25316 28908 25344
rect 28859 25313 28871 25316
rect 28813 25307 28871 25313
rect 28902 25304 28908 25316
rect 28960 25304 28966 25356
rect 29086 25304 29092 25356
rect 29144 25344 29150 25356
rect 30208 25344 30236 25375
rect 30466 25372 30472 25424
rect 30524 25412 30530 25424
rect 30561 25415 30619 25421
rect 30561 25412 30573 25415
rect 30524 25384 30573 25412
rect 30524 25372 30530 25384
rect 30561 25381 30573 25384
rect 30607 25381 30619 25415
rect 37274 25412 37280 25424
rect 30561 25375 30619 25381
rect 34532 25384 37280 25412
rect 34532 25356 34560 25384
rect 29144 25316 29684 25344
rect 30208 25316 31156 25344
rect 29144 25304 29150 25316
rect 25501 25279 25559 25285
rect 25501 25245 25513 25279
rect 25547 25276 25559 25279
rect 25593 25279 25651 25285
rect 25593 25276 25605 25279
rect 25547 25248 25605 25276
rect 25547 25245 25559 25248
rect 25501 25239 25559 25245
rect 25593 25245 25605 25248
rect 25639 25245 25651 25279
rect 25593 25239 25651 25245
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 26970 25236 26976 25288
rect 27028 25236 27034 25288
rect 27154 25236 27160 25288
rect 27212 25236 27218 25288
rect 29656 25285 29684 25316
rect 29641 25279 29699 25285
rect 29641 25245 29653 25279
rect 29687 25245 29699 25279
rect 29641 25239 29699 25245
rect 30282 25236 30288 25288
rect 30340 25236 30346 25288
rect 30377 25279 30435 25285
rect 30377 25245 30389 25279
rect 30423 25276 30435 25279
rect 30742 25276 30748 25288
rect 30423 25248 30748 25276
rect 30423 25245 30435 25248
rect 30377 25239 30435 25245
rect 30742 25236 30748 25248
rect 30800 25236 30806 25288
rect 30837 25279 30895 25285
rect 30837 25245 30849 25279
rect 30883 25276 30895 25279
rect 30926 25276 30932 25288
rect 30883 25248 30932 25276
rect 30883 25245 30895 25248
rect 30837 25239 30895 25245
rect 30926 25236 30932 25248
rect 30984 25236 30990 25288
rect 31128 25285 31156 25316
rect 34514 25304 34520 25356
rect 34572 25304 34578 25356
rect 34790 25304 34796 25356
rect 34848 25344 34854 25356
rect 36170 25344 36176 25356
rect 34848 25316 36176 25344
rect 34848 25304 34854 25316
rect 31113 25279 31171 25285
rect 31113 25245 31125 25279
rect 31159 25276 31171 25279
rect 32582 25276 32588 25288
rect 31159 25248 32588 25276
rect 31159 25245 31171 25248
rect 31113 25239 31171 25245
rect 32582 25236 32588 25248
rect 32640 25236 32646 25288
rect 35250 25236 35256 25288
rect 35308 25276 35314 25288
rect 35728 25285 35756 25316
rect 36170 25304 36176 25316
rect 36228 25304 36234 25356
rect 36446 25304 36452 25356
rect 36504 25344 36510 25356
rect 36504 25316 36676 25344
rect 36504 25304 36510 25316
rect 35437 25279 35495 25285
rect 35437 25276 35449 25279
rect 35308 25248 35449 25276
rect 35308 25236 35314 25248
rect 35437 25245 35449 25248
rect 35483 25245 35495 25279
rect 35437 25239 35495 25245
rect 35713 25279 35771 25285
rect 35713 25245 35725 25279
rect 35759 25245 35771 25279
rect 35713 25239 35771 25245
rect 35986 25236 35992 25288
rect 36044 25236 36050 25288
rect 36357 25279 36415 25285
rect 36357 25245 36369 25279
rect 36403 25276 36415 25279
rect 36538 25276 36544 25288
rect 36403 25248 36544 25276
rect 36403 25245 36415 25248
rect 36357 25239 36415 25245
rect 36538 25236 36544 25248
rect 36596 25236 36602 25288
rect 36648 25285 36676 25316
rect 37016 25285 37044 25384
rect 37274 25372 37280 25384
rect 37332 25372 37338 25424
rect 36633 25279 36691 25285
rect 36633 25245 36645 25279
rect 36679 25245 36691 25279
rect 36633 25239 36691 25245
rect 37001 25279 37059 25285
rect 37001 25245 37013 25279
rect 37047 25245 37059 25279
rect 37001 25239 37059 25245
rect 23382 25168 23388 25220
rect 23440 25168 23446 25220
rect 23566 25217 23572 25220
rect 23523 25211 23572 25217
rect 23523 25177 23535 25211
rect 23569 25177 23572 25211
rect 23523 25171 23572 25177
rect 23566 25168 23572 25171
rect 23624 25208 23630 25220
rect 24596 25208 24624 25236
rect 23624 25180 24624 25208
rect 23624 25168 23630 25180
rect 25314 25168 25320 25220
rect 25372 25168 25378 25220
rect 25866 25168 25872 25220
rect 25924 25208 25930 25220
rect 25961 25211 26019 25217
rect 25961 25208 25973 25211
rect 25924 25180 25973 25208
rect 25924 25168 25930 25180
rect 25961 25177 25973 25180
rect 26007 25177 26019 25211
rect 30009 25211 30067 25217
rect 30009 25208 30021 25211
rect 25961 25171 26019 25177
rect 26068 25180 30021 25208
rect 26068 25140 26096 25180
rect 30009 25177 30021 25180
rect 30055 25177 30067 25211
rect 30009 25171 30067 25177
rect 30561 25211 30619 25217
rect 30561 25177 30573 25211
rect 30607 25208 30619 25211
rect 30607 25180 30880 25208
rect 30607 25177 30619 25180
rect 30561 25171 30619 25177
rect 30852 25152 30880 25180
rect 32490 25168 32496 25220
rect 32548 25168 32554 25220
rect 33778 25168 33784 25220
rect 33836 25168 33842 25220
rect 34238 25168 34244 25220
rect 34296 25168 34302 25220
rect 34514 25168 34520 25220
rect 34572 25208 34578 25220
rect 35529 25211 35587 25217
rect 35529 25208 35541 25211
rect 34572 25180 35541 25208
rect 34572 25168 34578 25180
rect 35529 25177 35541 25180
rect 35575 25177 35587 25211
rect 35529 25171 35587 25177
rect 23124 25112 26096 25140
rect 27065 25143 27123 25149
rect 27065 25109 27077 25143
rect 27111 25140 27123 25143
rect 27430 25140 27436 25152
rect 27111 25112 27436 25140
rect 27111 25109 27123 25112
rect 27065 25103 27123 25109
rect 27430 25100 27436 25112
rect 27488 25100 27494 25152
rect 28534 25100 28540 25152
rect 28592 25100 28598 25152
rect 28626 25100 28632 25152
rect 28684 25100 28690 25152
rect 29086 25100 29092 25152
rect 29144 25140 29150 25152
rect 29730 25140 29736 25152
rect 29144 25112 29736 25140
rect 29144 25100 29150 25112
rect 29730 25100 29736 25112
rect 29788 25100 29794 25152
rect 30650 25100 30656 25152
rect 30708 25100 30714 25152
rect 30834 25100 30840 25152
rect 30892 25100 30898 25152
rect 31021 25143 31079 25149
rect 31021 25109 31033 25143
rect 31067 25140 31079 25143
rect 31570 25140 31576 25152
rect 31067 25112 31576 25140
rect 31067 25109 31079 25112
rect 31021 25103 31079 25109
rect 31570 25100 31576 25112
rect 31628 25100 31634 25152
rect 35342 25100 35348 25152
rect 35400 25140 35406 25152
rect 35437 25143 35495 25149
rect 35437 25140 35449 25143
rect 35400 25112 35449 25140
rect 35400 25100 35406 25112
rect 35437 25109 35449 25112
rect 35483 25109 35495 25143
rect 35544 25140 35572 25171
rect 35894 25168 35900 25220
rect 35952 25168 35958 25220
rect 36173 25211 36231 25217
rect 36173 25177 36185 25211
rect 36219 25208 36231 25211
rect 36262 25208 36268 25220
rect 36219 25180 36268 25208
rect 36219 25177 36231 25180
rect 36173 25171 36231 25177
rect 36262 25168 36268 25180
rect 36320 25168 36326 25220
rect 36541 25143 36599 25149
rect 36541 25140 36553 25143
rect 35544 25112 36553 25140
rect 35437 25103 35495 25109
rect 36541 25109 36553 25112
rect 36587 25140 36599 25143
rect 38562 25140 38568 25152
rect 36587 25112 38568 25140
rect 36587 25109 36599 25112
rect 36541 25103 36599 25109
rect 38562 25100 38568 25112
rect 38620 25100 38626 25152
rect 40328 25140 40356 25443
rect 41782 25440 41788 25492
rect 41840 25480 41846 25492
rect 41877 25483 41935 25489
rect 41877 25480 41889 25483
rect 41840 25452 41889 25480
rect 41840 25440 41846 25452
rect 41877 25449 41889 25452
rect 41923 25449 41935 25483
rect 41877 25443 41935 25449
rect 40586 25236 40592 25288
rect 40644 25276 40650 25288
rect 41325 25279 41383 25285
rect 41325 25276 41337 25279
rect 40644 25248 41337 25276
rect 40644 25236 40650 25248
rect 41325 25245 41337 25248
rect 41371 25245 41383 25279
rect 41800 25276 41828 25440
rect 41325 25239 41383 25245
rect 41708 25248 41828 25276
rect 40494 25168 40500 25220
rect 40552 25168 40558 25220
rect 40681 25211 40739 25217
rect 40681 25177 40693 25211
rect 40727 25177 40739 25211
rect 40681 25171 40739 25177
rect 40696 25140 40724 25171
rect 40954 25168 40960 25220
rect 41012 25208 41018 25220
rect 41708 25208 41736 25248
rect 41012 25180 41736 25208
rect 41785 25211 41843 25217
rect 41012 25168 41018 25180
rect 41785 25177 41797 25211
rect 41831 25208 41843 25211
rect 41966 25208 41972 25220
rect 41831 25180 41972 25208
rect 41831 25177 41843 25180
rect 41785 25171 41843 25177
rect 40328 25112 40724 25140
rect 40770 25100 40776 25152
rect 40828 25140 40834 25152
rect 40865 25143 40923 25149
rect 40865 25140 40877 25143
rect 40828 25112 40877 25140
rect 40828 25100 40834 25112
rect 40865 25109 40877 25112
rect 40911 25109 40923 25143
rect 40865 25103 40923 25109
rect 41506 25100 41512 25152
rect 41564 25100 41570 25152
rect 41598 25100 41604 25152
rect 41656 25140 41662 25152
rect 41800 25140 41828 25171
rect 41966 25168 41972 25180
rect 42024 25168 42030 25220
rect 41656 25112 41828 25140
rect 41656 25100 41662 25112
rect 1104 25050 42504 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 42504 25050
rect 1104 24976 42504 24998
rect 4706 24936 4712 24948
rect 3804 24908 4712 24936
rect 1394 24760 1400 24812
rect 1452 24760 1458 24812
rect 2682 24760 2688 24812
rect 2740 24800 2746 24812
rect 3804 24809 3832 24908
rect 4706 24896 4712 24908
rect 4764 24896 4770 24948
rect 7193 24939 7251 24945
rect 7193 24905 7205 24939
rect 7239 24936 7251 24939
rect 7282 24936 7288 24948
rect 7239 24908 7288 24936
rect 7239 24905 7251 24908
rect 7193 24899 7251 24905
rect 7282 24896 7288 24908
rect 7340 24896 7346 24948
rect 7561 24939 7619 24945
rect 7561 24905 7573 24939
rect 7607 24936 7619 24939
rect 7926 24936 7932 24948
rect 7607 24908 7932 24936
rect 7607 24905 7619 24908
rect 7561 24899 7619 24905
rect 7926 24896 7932 24908
rect 7984 24896 7990 24948
rect 8110 24896 8116 24948
rect 8168 24936 8174 24948
rect 8205 24939 8263 24945
rect 8205 24936 8217 24939
rect 8168 24908 8217 24936
rect 8168 24896 8174 24908
rect 8205 24905 8217 24908
rect 8251 24905 8263 24939
rect 8205 24899 8263 24905
rect 8386 24896 8392 24948
rect 8444 24936 8450 24948
rect 8849 24939 8907 24945
rect 8849 24936 8861 24939
rect 8444 24908 8861 24936
rect 8444 24896 8450 24908
rect 8849 24905 8861 24908
rect 8895 24905 8907 24939
rect 8849 24899 8907 24905
rect 12805 24939 12863 24945
rect 12805 24905 12817 24939
rect 12851 24936 12863 24939
rect 13630 24936 13636 24948
rect 12851 24908 13636 24936
rect 12851 24905 12863 24908
rect 12805 24899 12863 24905
rect 13630 24896 13636 24908
rect 13688 24896 13694 24948
rect 16114 24896 16120 24948
rect 16172 24936 16178 24948
rect 17218 24936 17224 24948
rect 16172 24908 17224 24936
rect 16172 24896 16178 24908
rect 17218 24896 17224 24908
rect 17276 24896 17282 24948
rect 19334 24936 19340 24948
rect 19168 24908 19340 24936
rect 5350 24868 5356 24880
rect 4724 24840 4936 24868
rect 3697 24803 3755 24809
rect 3697 24800 3709 24803
rect 2740 24772 3709 24800
rect 2740 24760 2746 24772
rect 3697 24769 3709 24772
rect 3743 24769 3755 24803
rect 3697 24763 3755 24769
rect 3789 24803 3847 24809
rect 3789 24769 3801 24803
rect 3835 24769 3847 24803
rect 3789 24763 3847 24769
rect 3878 24760 3884 24812
rect 3936 24760 3942 24812
rect 4430 24760 4436 24812
rect 4488 24760 4494 24812
rect 4522 24760 4528 24812
rect 4580 24760 4586 24812
rect 4614 24760 4620 24812
rect 4672 24760 4678 24812
rect 4065 24735 4123 24741
rect 4065 24701 4077 24735
rect 4111 24732 4123 24735
rect 4540 24732 4568 24760
rect 4111 24704 4568 24732
rect 4111 24701 4123 24704
rect 4065 24695 4123 24701
rect 1302 24624 1308 24676
rect 1360 24664 1366 24676
rect 1581 24667 1639 24673
rect 1581 24664 1593 24667
rect 1360 24636 1593 24664
rect 1360 24624 1366 24636
rect 1581 24633 1593 24636
rect 1627 24633 1639 24667
rect 4157 24667 4215 24673
rect 4157 24664 4169 24667
rect 1581 24627 1639 24633
rect 2746 24636 4169 24664
rect 2498 24556 2504 24608
rect 2556 24596 2562 24608
rect 2746 24596 2774 24636
rect 4157 24633 4169 24636
rect 4203 24633 4215 24667
rect 4157 24627 4215 24633
rect 2556 24568 2774 24596
rect 2556 24556 2562 24568
rect 3970 24556 3976 24608
rect 4028 24596 4034 24608
rect 4724 24596 4752 24840
rect 4908 24809 4936 24840
rect 5092 24840 5356 24868
rect 5092 24812 5120 24840
rect 5350 24828 5356 24840
rect 5408 24828 5414 24880
rect 7101 24871 7159 24877
rect 7101 24837 7113 24871
rect 7147 24868 7159 24871
rect 7374 24868 7380 24880
rect 7147 24840 7380 24868
rect 7147 24837 7159 24840
rect 7101 24831 7159 24837
rect 7374 24828 7380 24840
rect 7432 24828 7438 24880
rect 8174 24840 9352 24868
rect 8174 24812 8202 24840
rect 4801 24803 4859 24809
rect 4801 24769 4813 24803
rect 4847 24769 4859 24803
rect 4801 24763 4859 24769
rect 4893 24803 4951 24809
rect 4893 24769 4905 24803
rect 4939 24769 4951 24803
rect 4893 24763 4951 24769
rect 4816 24732 4844 24763
rect 5074 24760 5080 24812
rect 5132 24760 5138 24812
rect 5258 24760 5264 24812
rect 5316 24760 5322 24812
rect 6178 24760 6184 24812
rect 6236 24800 6242 24812
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 6236 24772 6561 24800
rect 6236 24760 6242 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 6733 24803 6791 24809
rect 6733 24769 6745 24803
rect 6779 24800 6791 24803
rect 6825 24803 6883 24809
rect 6825 24800 6837 24803
rect 6779 24772 6837 24800
rect 6779 24769 6791 24772
rect 6733 24763 6791 24769
rect 6825 24769 6837 24772
rect 6871 24798 6883 24803
rect 6914 24798 6920 24812
rect 6871 24770 6920 24798
rect 6871 24769 6883 24770
rect 6825 24763 6883 24769
rect 4985 24735 5043 24741
rect 4985 24732 4997 24735
rect 4816 24704 4997 24732
rect 4985 24701 4997 24704
rect 5031 24701 5043 24735
rect 4985 24695 5043 24701
rect 6086 24692 6092 24744
rect 6144 24692 6150 24744
rect 4028 24568 4752 24596
rect 6564 24596 6592 24763
rect 6914 24760 6920 24770
rect 6972 24760 6978 24812
rect 7193 24803 7251 24809
rect 7193 24800 7205 24803
rect 7024 24772 7205 24800
rect 6641 24735 6699 24741
rect 6641 24701 6653 24735
rect 6687 24732 6699 24735
rect 7024 24732 7052 24772
rect 7193 24769 7205 24772
rect 7239 24800 7251 24803
rect 7745 24803 7803 24809
rect 7745 24800 7757 24803
rect 7239 24772 7757 24800
rect 7239 24769 7251 24772
rect 7193 24763 7251 24769
rect 7745 24769 7757 24772
rect 7791 24769 7803 24803
rect 7745 24763 7803 24769
rect 7837 24803 7895 24809
rect 7837 24769 7849 24803
rect 7883 24769 7895 24803
rect 7837 24763 7895 24769
rect 7929 24806 7987 24809
rect 8174 24806 8208 24812
rect 7929 24803 8208 24806
rect 7929 24769 7941 24803
rect 7975 24778 8208 24803
rect 7975 24769 7987 24778
rect 7929 24763 7987 24769
rect 6687 24704 7052 24732
rect 6687 24701 6699 24704
rect 6641 24695 6699 24701
rect 7098 24692 7104 24744
rect 7156 24692 7162 24744
rect 7466 24692 7472 24744
rect 7524 24692 7530 24744
rect 7558 24692 7564 24744
rect 7616 24732 7622 24744
rect 7852 24732 7880 24763
rect 8202 24760 8208 24778
rect 8260 24760 8266 24812
rect 8294 24760 8300 24812
rect 8352 24800 8358 24812
rect 8588 24809 8616 24840
rect 8481 24803 8539 24809
rect 8481 24800 8493 24803
rect 8352 24772 8493 24800
rect 8352 24760 8358 24772
rect 8481 24769 8493 24772
rect 8527 24769 8539 24803
rect 8481 24763 8539 24769
rect 8573 24803 8631 24809
rect 8573 24769 8585 24803
rect 8619 24769 8631 24803
rect 8573 24763 8631 24769
rect 9030 24760 9036 24812
rect 9088 24760 9094 24812
rect 9214 24760 9220 24812
rect 9272 24760 9278 24812
rect 9324 24809 9352 24840
rect 9582 24828 9588 24880
rect 9640 24868 9646 24880
rect 13449 24871 13507 24877
rect 9640 24840 10088 24868
rect 9640 24828 9646 24840
rect 9309 24803 9367 24809
rect 9309 24769 9321 24803
rect 9355 24769 9367 24803
rect 9309 24763 9367 24769
rect 9490 24760 9496 24812
rect 9548 24800 9554 24812
rect 10060 24809 10088 24840
rect 13449 24837 13461 24871
rect 13495 24868 13507 24871
rect 13495 24840 14688 24868
rect 13495 24837 13507 24840
rect 13449 24831 13507 24837
rect 9677 24803 9735 24809
rect 9677 24800 9689 24803
rect 9548 24772 9689 24800
rect 9548 24760 9554 24772
rect 9677 24769 9689 24772
rect 9723 24769 9735 24803
rect 9677 24763 9735 24769
rect 9861 24803 9919 24809
rect 9861 24769 9873 24803
rect 9907 24769 9919 24803
rect 9861 24763 9919 24769
rect 9953 24803 10011 24809
rect 9953 24769 9965 24803
rect 9999 24769 10011 24803
rect 9953 24763 10011 24769
rect 10045 24803 10103 24809
rect 10045 24769 10057 24803
rect 10091 24800 10103 24803
rect 10091 24772 12434 24800
rect 10091 24769 10103 24772
rect 10045 24763 10103 24769
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 7616 24704 7880 24732
rect 7918 24704 8033 24732
rect 7616 24692 7622 24704
rect 6822 24624 6828 24676
rect 6880 24664 6886 24676
rect 7285 24667 7343 24673
rect 7285 24664 7297 24667
rect 6880 24636 7297 24664
rect 6880 24624 6886 24636
rect 7285 24633 7297 24636
rect 7331 24664 7343 24667
rect 7742 24664 7748 24676
rect 7331 24636 7748 24664
rect 7331 24633 7343 24636
rect 7285 24627 7343 24633
rect 7742 24624 7748 24636
rect 7800 24664 7806 24676
rect 7918 24664 7946 24704
rect 8021 24701 8033 24704
rect 8067 24701 8079 24735
rect 8021 24695 8079 24701
rect 8386 24692 8392 24744
rect 8444 24692 8450 24744
rect 8665 24735 8723 24741
rect 8665 24701 8677 24735
rect 8711 24732 8723 24735
rect 8846 24732 8852 24744
rect 8711 24704 8852 24732
rect 8711 24701 8723 24704
rect 8665 24695 8723 24701
rect 8846 24692 8852 24704
rect 8904 24692 8910 24744
rect 9232 24732 9260 24760
rect 9876 24732 9904 24763
rect 9232 24704 9904 24732
rect 9968 24732 9996 24763
rect 10318 24732 10324 24744
rect 9968 24704 10324 24732
rect 10318 24692 10324 24704
rect 10376 24692 10382 24744
rect 11149 24735 11207 24741
rect 11149 24701 11161 24735
rect 11195 24732 11207 24735
rect 11330 24732 11336 24744
rect 11195 24704 11336 24732
rect 11195 24701 11207 24704
rect 11149 24695 11207 24701
rect 11330 24692 11336 24704
rect 11388 24692 11394 24744
rect 12066 24692 12072 24744
rect 12124 24692 12130 24744
rect 12406 24732 12434 24772
rect 12710 24760 12716 24812
rect 12768 24760 12774 24812
rect 13725 24803 13783 24809
rect 13725 24769 13737 24803
rect 13771 24800 13783 24803
rect 13814 24800 13820 24812
rect 13771 24772 13820 24800
rect 13771 24769 13783 24772
rect 13725 24763 13783 24769
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 14366 24760 14372 24812
rect 14424 24760 14430 24812
rect 14660 24809 14688 24840
rect 15010 24828 15016 24880
rect 15068 24868 15074 24880
rect 17586 24868 17592 24880
rect 15068 24840 17592 24868
rect 15068 24828 15074 24840
rect 14645 24803 14703 24809
rect 14645 24769 14657 24803
rect 14691 24769 14703 24803
rect 14645 24763 14703 24769
rect 14734 24760 14740 24812
rect 14792 24760 14798 24812
rect 14918 24760 14924 24812
rect 14976 24760 14982 24812
rect 15654 24760 15660 24812
rect 15712 24760 15718 24812
rect 15856 24809 15884 24840
rect 17586 24828 17592 24840
rect 17644 24828 17650 24880
rect 15841 24803 15899 24809
rect 15841 24769 15853 24803
rect 15887 24769 15899 24803
rect 15841 24763 15899 24769
rect 15930 24760 15936 24812
rect 15988 24760 15994 24812
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24800 17187 24803
rect 18414 24800 18420 24812
rect 17175 24772 18420 24800
rect 17175 24769 17187 24772
rect 17129 24763 17187 24769
rect 18414 24760 18420 24772
rect 18472 24760 18478 24812
rect 19168 24809 19196 24908
rect 19334 24896 19340 24908
rect 19392 24896 19398 24948
rect 19610 24936 19616 24948
rect 19536 24908 19616 24936
rect 19153 24803 19211 24809
rect 19153 24769 19165 24803
rect 19199 24769 19211 24803
rect 19153 24763 19211 24769
rect 19337 24803 19395 24809
rect 19337 24769 19349 24803
rect 19383 24800 19395 24803
rect 19536 24800 19564 24908
rect 19610 24896 19616 24908
rect 19668 24896 19674 24948
rect 20165 24939 20223 24945
rect 20165 24905 20177 24939
rect 20211 24936 20223 24939
rect 21358 24936 21364 24948
rect 20211 24908 21364 24936
rect 20211 24905 20223 24908
rect 20165 24899 20223 24905
rect 21358 24896 21364 24908
rect 21416 24896 21422 24948
rect 22186 24896 22192 24948
rect 22244 24936 22250 24948
rect 22370 24936 22376 24948
rect 22244 24908 22376 24936
rect 22244 24896 22250 24908
rect 22370 24896 22376 24908
rect 22428 24896 22434 24948
rect 25041 24939 25099 24945
rect 25041 24905 25053 24939
rect 25087 24936 25099 24939
rect 25314 24936 25320 24948
rect 25087 24908 25320 24936
rect 25087 24905 25099 24908
rect 25041 24899 25099 24905
rect 25314 24896 25320 24908
rect 25372 24896 25378 24948
rect 25415 24908 27292 24936
rect 19797 24871 19855 24877
rect 19797 24837 19809 24871
rect 19843 24868 19855 24871
rect 19843 24840 20208 24868
rect 19843 24837 19855 24840
rect 19797 24831 19855 24837
rect 20180 24812 20208 24840
rect 21266 24828 21272 24880
rect 21324 24868 21330 24880
rect 21324 24840 23336 24868
rect 21324 24828 21330 24840
rect 19613 24803 19671 24809
rect 19613 24800 19625 24803
rect 19383 24772 19625 24800
rect 19383 24769 19395 24772
rect 19337 24763 19395 24769
rect 19613 24769 19625 24772
rect 19659 24769 19671 24803
rect 19613 24763 19671 24769
rect 19889 24803 19947 24809
rect 19889 24769 19901 24803
rect 19935 24769 19947 24803
rect 19889 24763 19947 24769
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24769 20131 24803
rect 20073 24763 20131 24769
rect 14553 24735 14611 24741
rect 12406 24704 13400 24732
rect 7800 24636 7946 24664
rect 7800 24624 7806 24636
rect 9582 24624 9588 24676
rect 9640 24664 9646 24676
rect 10505 24667 10563 24673
rect 10505 24664 10517 24667
rect 9640 24636 10517 24664
rect 9640 24624 9646 24636
rect 10505 24633 10517 24636
rect 10551 24633 10563 24667
rect 11348 24664 11376 24692
rect 12345 24667 12403 24673
rect 12345 24664 12357 24667
rect 11348 24636 12357 24664
rect 10505 24627 10563 24633
rect 12345 24633 12357 24636
rect 12391 24664 12403 24667
rect 12802 24664 12808 24676
rect 12391 24636 12808 24664
rect 12391 24633 12403 24636
rect 12345 24627 12403 24633
rect 12802 24624 12808 24636
rect 12860 24624 12866 24676
rect 6917 24599 6975 24605
rect 6917 24596 6929 24599
rect 6564 24568 6929 24596
rect 4028 24556 4034 24568
rect 6917 24565 6929 24568
rect 6963 24596 6975 24599
rect 7006 24596 7012 24608
rect 6963 24568 7012 24596
rect 6963 24565 6975 24568
rect 6917 24559 6975 24565
rect 7006 24556 7012 24568
rect 7064 24556 7070 24608
rect 7190 24556 7196 24608
rect 7248 24596 7254 24608
rect 7926 24596 7932 24608
rect 7248 24568 7932 24596
rect 7248 24556 7254 24568
rect 7926 24556 7932 24568
rect 7984 24556 7990 24608
rect 10226 24556 10232 24608
rect 10284 24556 10290 24608
rect 12526 24556 12532 24608
rect 12584 24556 12590 24608
rect 12986 24556 12992 24608
rect 13044 24556 13050 24608
rect 13078 24556 13084 24608
rect 13136 24556 13142 24608
rect 13170 24556 13176 24608
rect 13228 24556 13234 24608
rect 13372 24596 13400 24704
rect 14553 24701 14565 24735
rect 14599 24732 14611 24735
rect 14599 24704 14688 24732
rect 14599 24701 14611 24704
rect 14553 24695 14611 24701
rect 14660 24664 14688 24704
rect 18138 24692 18144 24744
rect 18196 24692 18202 24744
rect 19168 24732 19196 24763
rect 19429 24735 19487 24741
rect 19429 24732 19441 24735
rect 19168 24704 19441 24732
rect 19429 24701 19441 24704
rect 19475 24701 19487 24735
rect 19429 24695 19487 24701
rect 19518 24692 19524 24744
rect 19576 24732 19582 24744
rect 19904 24732 19932 24763
rect 19576 24704 19932 24732
rect 19576 24692 19582 24704
rect 15470 24664 15476 24676
rect 14660 24636 15476 24664
rect 15470 24624 15476 24636
rect 15528 24624 15534 24676
rect 15654 24624 15660 24676
rect 15712 24664 15718 24676
rect 18156 24664 18184 24692
rect 20088 24676 20116 24763
rect 20162 24760 20168 24812
rect 20220 24800 20226 24812
rect 20349 24803 20407 24809
rect 20349 24800 20361 24803
rect 20220 24772 20361 24800
rect 20220 24760 20226 24772
rect 20349 24769 20361 24772
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 22278 24760 22284 24812
rect 22336 24760 22342 24812
rect 22925 24803 22983 24809
rect 22925 24769 22937 24803
rect 22971 24800 22983 24803
rect 23106 24800 23112 24812
rect 22971 24772 23112 24800
rect 22971 24769 22983 24772
rect 22925 24763 22983 24769
rect 23106 24760 23112 24772
rect 23164 24760 23170 24812
rect 23308 24800 23336 24840
rect 23382 24828 23388 24880
rect 23440 24868 23446 24880
rect 25415 24868 25443 24908
rect 23440 24840 25443 24868
rect 23440 24828 23446 24840
rect 25682 24828 25688 24880
rect 25740 24828 25746 24880
rect 25866 24868 25872 24880
rect 25924 24877 25930 24880
rect 25924 24871 25943 24877
rect 25792 24840 25872 24868
rect 24670 24800 24676 24812
rect 23308 24772 24676 24800
rect 24670 24760 24676 24772
rect 24728 24800 24734 24812
rect 24765 24803 24823 24809
rect 24765 24800 24777 24803
rect 24728 24772 24777 24800
rect 24728 24760 24734 24772
rect 24765 24769 24777 24772
rect 24811 24769 24823 24803
rect 24765 24763 24823 24769
rect 25222 24760 25228 24812
rect 25280 24800 25286 24812
rect 25317 24803 25375 24809
rect 25317 24800 25329 24803
rect 25280 24772 25329 24800
rect 25280 24760 25286 24772
rect 25317 24769 25329 24772
rect 25363 24800 25375 24803
rect 25792 24800 25820 24840
rect 25866 24828 25872 24840
rect 25931 24837 25943 24871
rect 25924 24831 25943 24837
rect 25924 24828 25930 24831
rect 26050 24828 26056 24880
rect 26108 24868 26114 24880
rect 26513 24871 26571 24877
rect 26513 24868 26525 24871
rect 26108 24840 26525 24868
rect 26108 24828 26114 24840
rect 26513 24837 26525 24840
rect 26559 24837 26571 24871
rect 26513 24831 26571 24837
rect 26326 24800 26332 24812
rect 25363 24772 25820 24800
rect 25884 24772 26332 24800
rect 25363 24769 25375 24772
rect 25317 24763 25375 24769
rect 22465 24735 22523 24741
rect 22465 24701 22477 24735
rect 22511 24732 22523 24735
rect 25038 24732 25044 24744
rect 22511 24704 25044 24732
rect 22511 24701 22523 24704
rect 22465 24695 22523 24701
rect 25038 24692 25044 24704
rect 25096 24692 25102 24744
rect 25498 24692 25504 24744
rect 25556 24732 25562 24744
rect 25556 24704 25636 24732
rect 25556 24692 25562 24704
rect 15712 24636 18184 24664
rect 15712 24624 15718 24636
rect 18322 24624 18328 24676
rect 18380 24664 18386 24676
rect 18417 24667 18475 24673
rect 18417 24664 18429 24667
rect 18380 24636 18429 24664
rect 18380 24624 18386 24636
rect 18417 24633 18429 24636
rect 18463 24633 18475 24667
rect 18417 24627 18475 24633
rect 19337 24667 19395 24673
rect 19337 24633 19349 24667
rect 19383 24664 19395 24667
rect 20070 24664 20076 24676
rect 19383 24636 20076 24664
rect 19383 24633 19395 24636
rect 19337 24627 19395 24633
rect 20070 24624 20076 24636
rect 20128 24624 20134 24676
rect 22738 24624 22744 24676
rect 22796 24624 22802 24676
rect 24854 24624 24860 24676
rect 24912 24664 24918 24676
rect 25133 24667 25191 24673
rect 25133 24664 25145 24667
rect 24912 24636 25145 24664
rect 24912 24624 24918 24636
rect 25133 24633 25145 24636
rect 25179 24633 25191 24667
rect 25133 24627 25191 24633
rect 13998 24596 14004 24608
rect 13372 24568 14004 24596
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 14182 24556 14188 24608
rect 14240 24556 14246 24608
rect 15378 24556 15384 24608
rect 15436 24596 15442 24608
rect 15930 24596 15936 24608
rect 15436 24568 15936 24596
rect 15436 24556 15442 24568
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 17034 24556 17040 24608
rect 17092 24556 17098 24608
rect 18598 24556 18604 24608
rect 18656 24556 18662 24608
rect 21818 24556 21824 24608
rect 21876 24556 21882 24608
rect 25314 24556 25320 24608
rect 25372 24596 25378 24608
rect 25608 24596 25636 24704
rect 25682 24692 25688 24744
rect 25740 24732 25746 24744
rect 25884 24732 25912 24772
rect 26326 24760 26332 24772
rect 26384 24760 26390 24812
rect 27264 24809 27292 24908
rect 28626 24896 28632 24948
rect 28684 24936 28690 24948
rect 28721 24939 28779 24945
rect 28721 24936 28733 24939
rect 28684 24908 28733 24936
rect 28684 24896 28690 24908
rect 28721 24905 28733 24908
rect 28767 24905 28779 24939
rect 30282 24936 30288 24948
rect 28721 24899 28779 24905
rect 28920 24908 30288 24936
rect 27430 24828 27436 24880
rect 27488 24828 27494 24880
rect 27798 24868 27804 24880
rect 27540 24840 27804 24868
rect 27540 24812 27568 24840
rect 27798 24828 27804 24840
rect 27856 24828 27862 24880
rect 28810 24868 28816 24880
rect 27908 24840 28816 24868
rect 26421 24803 26479 24809
rect 26421 24769 26433 24803
rect 26467 24769 26479 24803
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 26421 24763 26479 24769
rect 26528 24772 27169 24800
rect 26436 24732 26464 24763
rect 26528 24744 26556 24772
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 27250 24803 27308 24809
rect 27250 24769 27262 24803
rect 27296 24769 27308 24803
rect 27250 24763 27308 24769
rect 27522 24760 27528 24812
rect 27580 24760 27586 24812
rect 27706 24809 27712 24812
rect 27663 24803 27712 24809
rect 27663 24769 27675 24803
rect 27709 24769 27712 24803
rect 27663 24763 27712 24769
rect 27706 24760 27712 24763
rect 27764 24800 27770 24812
rect 27908 24800 27936 24840
rect 28810 24828 28816 24840
rect 28868 24828 28874 24880
rect 27764 24772 27936 24800
rect 27764 24760 27770 24772
rect 27982 24760 27988 24812
rect 28040 24760 28046 24812
rect 28445 24803 28503 24809
rect 28445 24769 28457 24803
rect 28491 24769 28503 24803
rect 28445 24763 28503 24769
rect 25740 24704 25912 24732
rect 26068 24704 26464 24732
rect 25740 24692 25746 24704
rect 26068 24664 26096 24704
rect 26510 24692 26516 24744
rect 26568 24692 26574 24744
rect 26697 24735 26755 24741
rect 26697 24701 26709 24735
rect 26743 24732 26755 24735
rect 28460 24732 28488 24763
rect 28626 24760 28632 24812
rect 28684 24760 28690 24812
rect 28920 24809 28948 24908
rect 30282 24896 30288 24908
rect 30340 24896 30346 24948
rect 31846 24896 31852 24948
rect 31904 24936 31910 24948
rect 32674 24936 32680 24948
rect 31904 24908 32680 24936
rect 31904 24896 31910 24908
rect 32674 24896 32680 24908
rect 32732 24896 32738 24948
rect 33042 24896 33048 24948
rect 33100 24896 33106 24948
rect 33873 24939 33931 24945
rect 33873 24905 33885 24939
rect 33919 24936 33931 24939
rect 34238 24936 34244 24948
rect 33919 24908 34244 24936
rect 33919 24905 33931 24908
rect 33873 24899 33931 24905
rect 34238 24896 34244 24908
rect 34296 24896 34302 24948
rect 35250 24896 35256 24948
rect 35308 24936 35314 24948
rect 35308 24908 36584 24936
rect 35308 24896 35314 24908
rect 29012 24840 29408 24868
rect 29012 24809 29040 24840
rect 28905 24803 28963 24809
rect 28905 24769 28917 24803
rect 28951 24769 28963 24803
rect 28905 24763 28963 24769
rect 28997 24803 29055 24809
rect 28997 24769 29009 24803
rect 29043 24769 29055 24803
rect 28997 24763 29055 24769
rect 26743 24704 28488 24732
rect 26743 24701 26755 24704
rect 26697 24695 26755 24701
rect 27172 24676 27200 24704
rect 25884 24636 26096 24664
rect 26145 24667 26203 24673
rect 25884 24605 25912 24636
rect 26145 24633 26157 24667
rect 26191 24633 26203 24667
rect 26145 24627 26203 24633
rect 25869 24599 25927 24605
rect 25869 24596 25881 24599
rect 25372 24568 25881 24596
rect 25372 24556 25378 24568
rect 25869 24565 25881 24568
rect 25915 24565 25927 24599
rect 25869 24559 25927 24565
rect 26050 24556 26056 24608
rect 26108 24556 26114 24608
rect 26160 24596 26188 24627
rect 26234 24624 26240 24676
rect 26292 24664 26298 24676
rect 26292 24636 26832 24664
rect 26292 24624 26298 24636
rect 26694 24596 26700 24608
rect 26160 24568 26700 24596
rect 26694 24556 26700 24568
rect 26752 24556 26758 24608
rect 26804 24596 26832 24636
rect 27154 24624 27160 24676
rect 27212 24624 27218 24676
rect 27246 24624 27252 24676
rect 27304 24664 27310 24676
rect 28166 24664 28172 24676
rect 27304 24636 28172 24664
rect 27304 24624 27310 24636
rect 28166 24624 28172 24636
rect 28224 24624 28230 24676
rect 27706 24596 27712 24608
rect 26804 24568 27712 24596
rect 27706 24556 27712 24568
rect 27764 24556 27770 24608
rect 27798 24556 27804 24608
rect 27856 24556 27862 24608
rect 28460 24596 28488 24704
rect 28537 24735 28595 24741
rect 28537 24701 28549 24735
rect 28583 24732 28595 24735
rect 28920 24732 28948 24763
rect 29086 24760 29092 24812
rect 29144 24760 29150 24812
rect 29270 24809 29276 24812
rect 29227 24803 29276 24809
rect 29227 24769 29239 24803
rect 29273 24769 29276 24803
rect 29227 24763 29276 24769
rect 29270 24760 29276 24763
rect 29328 24760 29334 24812
rect 29380 24800 29408 24840
rect 29638 24828 29644 24880
rect 29696 24828 29702 24880
rect 31386 24828 31392 24880
rect 31444 24828 31450 24880
rect 32582 24828 32588 24880
rect 32640 24868 32646 24880
rect 33060 24868 33088 24896
rect 36556 24880 36584 24908
rect 40494 24896 40500 24948
rect 40552 24936 40558 24948
rect 40681 24939 40739 24945
rect 40681 24936 40693 24939
rect 40552 24908 40693 24936
rect 40552 24896 40558 24908
rect 40681 24905 40693 24908
rect 40727 24905 40739 24939
rect 40681 24899 40739 24905
rect 40862 24896 40868 24948
rect 40920 24936 40926 24948
rect 40920 24908 41092 24936
rect 40920 24896 40926 24908
rect 35805 24871 35863 24877
rect 35805 24868 35817 24871
rect 32640 24840 33180 24868
rect 32640 24828 32646 24840
rect 29457 24803 29515 24809
rect 29457 24800 29469 24803
rect 29380 24772 29469 24800
rect 29457 24769 29469 24772
rect 29503 24769 29515 24803
rect 29457 24763 29515 24769
rect 29822 24760 29828 24812
rect 29880 24760 29886 24812
rect 28583 24704 28948 24732
rect 29365 24735 29423 24741
rect 28583 24701 28595 24704
rect 28537 24695 28595 24701
rect 29365 24701 29377 24735
rect 29411 24732 29423 24735
rect 29546 24732 29552 24744
rect 29411 24704 29552 24732
rect 29411 24701 29423 24704
rect 29365 24695 29423 24701
rect 29546 24692 29552 24704
rect 29604 24692 29610 24744
rect 30101 24735 30159 24741
rect 30101 24701 30113 24735
rect 30147 24701 30159 24735
rect 30101 24695 30159 24701
rect 28902 24624 28908 24676
rect 28960 24664 28966 24676
rect 30116 24664 30144 24695
rect 30374 24692 30380 24744
rect 30432 24692 30438 24744
rect 31404 24732 31432 24828
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32677 24803 32735 24809
rect 32677 24769 32689 24803
rect 32723 24769 32735 24803
rect 32677 24763 32735 24769
rect 32125 24735 32183 24741
rect 32125 24732 32137 24735
rect 31404 24704 32137 24732
rect 32125 24701 32137 24704
rect 32171 24701 32183 24735
rect 32324 24732 32352 24763
rect 32582 24732 32588 24744
rect 32324 24704 32588 24732
rect 32125 24695 32183 24701
rect 32582 24692 32588 24704
rect 32640 24692 32646 24744
rect 32692 24664 32720 24763
rect 32766 24760 32772 24812
rect 32824 24800 32830 24812
rect 32824 24772 32869 24800
rect 32824 24760 32830 24772
rect 32950 24760 32956 24812
rect 33008 24760 33014 24812
rect 33152 24809 33180 24840
rect 33612 24840 33824 24868
rect 33045 24803 33103 24809
rect 33045 24769 33057 24803
rect 33091 24769 33103 24803
rect 33045 24763 33103 24769
rect 33142 24803 33200 24809
rect 33142 24769 33154 24803
rect 33188 24769 33200 24803
rect 33612 24800 33640 24840
rect 33142 24763 33200 24769
rect 33327 24772 33640 24800
rect 33060 24732 33088 24763
rect 33327 24732 33355 24772
rect 33686 24760 33692 24812
rect 33744 24760 33750 24812
rect 33796 24800 33824 24840
rect 35360 24840 35817 24868
rect 35360 24812 35388 24840
rect 35805 24837 35817 24840
rect 35851 24837 35863 24871
rect 36262 24868 36268 24880
rect 35805 24831 35863 24837
rect 35912 24840 36268 24868
rect 35069 24803 35127 24809
rect 35069 24800 35081 24803
rect 33796 24772 35081 24800
rect 35069 24769 35081 24772
rect 35115 24769 35127 24803
rect 35069 24763 35127 24769
rect 35158 24760 35164 24812
rect 35216 24800 35222 24812
rect 35253 24803 35311 24809
rect 35253 24800 35265 24803
rect 35216 24772 35265 24800
rect 35216 24760 35222 24772
rect 35253 24769 35265 24772
rect 35299 24769 35311 24803
rect 35253 24763 35311 24769
rect 35342 24760 35348 24812
rect 35400 24760 35406 24812
rect 35618 24809 35624 24812
rect 35437 24803 35495 24809
rect 35437 24802 35449 24803
rect 35483 24802 35495 24803
rect 35595 24803 35624 24809
rect 35434 24750 35440 24802
rect 35492 24750 35498 24802
rect 35595 24769 35607 24803
rect 35595 24763 35624 24769
rect 35618 24760 35624 24763
rect 35676 24760 35682 24812
rect 35912 24809 35940 24840
rect 36262 24828 36268 24840
rect 36320 24828 36326 24880
rect 36538 24828 36544 24880
rect 36596 24868 36602 24880
rect 36725 24871 36783 24877
rect 36725 24868 36737 24871
rect 36596 24840 36737 24868
rect 36596 24828 36602 24840
rect 36725 24837 36737 24840
rect 36771 24837 36783 24871
rect 36725 24831 36783 24837
rect 35713 24803 35771 24809
rect 35713 24769 35725 24803
rect 35759 24769 35771 24803
rect 35713 24763 35771 24769
rect 35897 24803 35955 24809
rect 35897 24769 35909 24803
rect 35943 24769 35955 24803
rect 35897 24763 35955 24769
rect 36081 24803 36139 24809
rect 36081 24769 36093 24803
rect 36127 24800 36139 24803
rect 36633 24803 36691 24809
rect 36633 24800 36645 24803
rect 36127 24772 36645 24800
rect 36127 24769 36139 24772
rect 36081 24763 36139 24769
rect 36633 24769 36645 24772
rect 36679 24769 36691 24803
rect 36633 24763 36691 24769
rect 33060 24704 33180 24732
rect 33152 24676 33180 24704
rect 33244 24704 33355 24732
rect 33413 24735 33471 24741
rect 28960 24636 30144 24664
rect 31404 24636 32720 24664
rect 28960 24624 28966 24636
rect 29822 24596 29828 24608
rect 28460 24568 29828 24596
rect 29822 24556 29828 24568
rect 29880 24556 29886 24608
rect 30926 24556 30932 24608
rect 30984 24596 30990 24608
rect 31404 24596 31432 24636
rect 33134 24624 33140 24676
rect 33192 24624 33198 24676
rect 30984 24568 31432 24596
rect 30984 24556 30990 24568
rect 31478 24556 31484 24608
rect 31536 24596 31542 24608
rect 33244 24596 33272 24704
rect 33413 24701 33425 24735
rect 33459 24732 33471 24735
rect 34514 24732 34520 24744
rect 33459 24704 34520 24732
rect 33459 24701 33471 24704
rect 33413 24695 33471 24701
rect 34514 24692 34520 24704
rect 34572 24692 34578 24744
rect 33321 24667 33379 24673
rect 33321 24633 33333 24667
rect 33367 24664 33379 24667
rect 33686 24664 33692 24676
rect 33367 24636 33692 24664
rect 33367 24633 33379 24636
rect 33321 24627 33379 24633
rect 33686 24624 33692 24636
rect 33744 24624 33750 24676
rect 35447 24664 35475 24750
rect 35728 24732 35756 24763
rect 36170 24732 36176 24744
rect 35728 24704 36176 24732
rect 36170 24692 36176 24704
rect 36228 24692 36234 24744
rect 36446 24692 36452 24744
rect 36504 24692 36510 24744
rect 36630 24664 36636 24676
rect 35447 24636 36636 24664
rect 36630 24624 36636 24636
rect 36688 24624 36694 24676
rect 36740 24664 36768 24831
rect 36998 24828 37004 24880
rect 37056 24868 37062 24880
rect 37274 24868 37280 24880
rect 37056 24840 37280 24868
rect 37056 24828 37062 24840
rect 37274 24828 37280 24840
rect 37332 24868 37338 24880
rect 37369 24871 37427 24877
rect 37369 24868 37381 24871
rect 37332 24840 37381 24868
rect 37332 24828 37338 24840
rect 37369 24837 37381 24840
rect 37415 24837 37427 24871
rect 37369 24831 37427 24837
rect 37384 24732 37412 24831
rect 39114 24828 39120 24880
rect 39172 24828 39178 24880
rect 39574 24828 39580 24880
rect 39632 24828 39638 24880
rect 41064 24877 41092 24908
rect 41049 24871 41107 24877
rect 41049 24837 41061 24871
rect 41095 24868 41107 24871
rect 41690 24868 41696 24880
rect 41095 24840 41696 24868
rect 41095 24837 41107 24840
rect 41049 24831 41107 24837
rect 41690 24828 41696 24840
rect 41748 24828 41754 24880
rect 41782 24828 41788 24880
rect 41840 24868 41846 24880
rect 42061 24871 42119 24877
rect 42061 24868 42073 24871
rect 41840 24840 42073 24868
rect 41840 24828 41846 24840
rect 42061 24837 42073 24840
rect 42107 24837 42119 24871
rect 42061 24831 42119 24837
rect 38197 24803 38255 24809
rect 38197 24769 38209 24803
rect 38243 24800 38255 24803
rect 38746 24800 38752 24812
rect 38243 24772 38752 24800
rect 38243 24769 38255 24772
rect 38197 24763 38255 24769
rect 38746 24760 38752 24772
rect 38804 24760 38810 24812
rect 40862 24760 40868 24812
rect 40920 24760 40926 24812
rect 40954 24760 40960 24812
rect 41012 24760 41018 24812
rect 41233 24803 41291 24809
rect 41233 24769 41245 24803
rect 41279 24800 41291 24803
rect 41322 24800 41328 24812
rect 41279 24772 41328 24800
rect 41279 24769 41291 24772
rect 41233 24763 41291 24769
rect 41322 24760 41328 24772
rect 41380 24760 41386 24812
rect 38841 24735 38899 24741
rect 38841 24732 38853 24735
rect 37384 24704 38853 24732
rect 38841 24701 38853 24704
rect 38887 24701 38899 24735
rect 38841 24695 38899 24701
rect 39574 24692 39580 24744
rect 39632 24732 39638 24744
rect 39632 24704 40163 24732
rect 39632 24692 39638 24704
rect 38746 24664 38752 24676
rect 36740 24636 38752 24664
rect 38746 24624 38752 24636
rect 38804 24624 38810 24676
rect 40135 24664 40163 24704
rect 40586 24692 40592 24744
rect 40644 24692 40650 24744
rect 41782 24664 41788 24676
rect 40135 24636 41788 24664
rect 41782 24624 41788 24636
rect 41840 24624 41846 24676
rect 31536 24568 33272 24596
rect 31536 24556 31542 24568
rect 33502 24556 33508 24608
rect 33560 24556 33566 24608
rect 34885 24599 34943 24605
rect 34885 24565 34897 24599
rect 34931 24596 34943 24599
rect 35618 24596 35624 24608
rect 34931 24568 35624 24596
rect 34931 24565 34943 24568
rect 34885 24559 34943 24565
rect 35618 24556 35624 24568
rect 35676 24556 35682 24608
rect 37093 24599 37151 24605
rect 37093 24565 37105 24599
rect 37139 24596 37151 24599
rect 37274 24596 37280 24608
rect 37139 24568 37280 24596
rect 37139 24565 37151 24568
rect 37093 24559 37151 24565
rect 37274 24556 37280 24568
rect 37332 24556 37338 24608
rect 38654 24556 38660 24608
rect 38712 24596 38718 24608
rect 39666 24596 39672 24608
rect 38712 24568 39672 24596
rect 38712 24556 38718 24568
rect 39666 24556 39672 24568
rect 39724 24596 39730 24608
rect 41414 24596 41420 24608
rect 39724 24568 41420 24596
rect 39724 24556 39730 24568
rect 41414 24556 41420 24568
rect 41472 24556 41478 24608
rect 41506 24556 41512 24608
rect 41564 24556 41570 24608
rect 1104 24506 42504 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 42504 24506
rect 1104 24432 42504 24454
rect 4893 24395 4951 24401
rect 4893 24392 4905 24395
rect 4356 24364 4905 24392
rect 1581 24259 1639 24265
rect 1581 24225 1593 24259
rect 1627 24256 1639 24259
rect 3510 24256 3516 24268
rect 1627 24228 3516 24256
rect 1627 24225 1639 24228
rect 1581 24219 1639 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 2958 24148 2964 24200
rect 3016 24148 3022 24200
rect 3605 24191 3663 24197
rect 3605 24157 3617 24191
rect 3651 24188 3663 24191
rect 3786 24188 3792 24200
rect 3651 24160 3792 24188
rect 3651 24157 3663 24160
rect 3605 24151 3663 24157
rect 3786 24148 3792 24160
rect 3844 24188 3850 24200
rect 4356 24197 4384 24364
rect 4893 24361 4905 24364
rect 4939 24361 4951 24395
rect 4893 24355 4951 24361
rect 5077 24395 5135 24401
rect 5077 24361 5089 24395
rect 5123 24392 5135 24395
rect 6546 24392 6552 24404
rect 5123 24364 6552 24392
rect 5123 24361 5135 24364
rect 5077 24355 5135 24361
rect 6546 24352 6552 24364
rect 6604 24352 6610 24404
rect 6733 24395 6791 24401
rect 6733 24361 6745 24395
rect 6779 24392 6791 24395
rect 7282 24392 7288 24404
rect 6779 24364 7288 24392
rect 6779 24361 6791 24364
rect 6733 24355 6791 24361
rect 7282 24352 7288 24364
rect 7340 24392 7346 24404
rect 7837 24395 7895 24401
rect 7837 24392 7849 24395
rect 7340 24364 7849 24392
rect 7340 24352 7346 24364
rect 7837 24361 7849 24364
rect 7883 24361 7895 24395
rect 7837 24355 7895 24361
rect 8018 24352 8024 24404
rect 8076 24352 8082 24404
rect 8386 24352 8392 24404
rect 8444 24392 8450 24404
rect 9217 24395 9275 24401
rect 9217 24392 9229 24395
rect 8444 24364 9229 24392
rect 8444 24352 8450 24364
rect 9217 24361 9229 24364
rect 9263 24392 9275 24395
rect 9306 24392 9312 24404
rect 9263 24364 9312 24392
rect 9263 24361 9275 24364
rect 9217 24355 9275 24361
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 11330 24352 11336 24404
rect 11388 24352 11394 24404
rect 12986 24352 12992 24404
rect 13044 24392 13050 24404
rect 13173 24395 13231 24401
rect 13173 24392 13185 24395
rect 13044 24364 13185 24392
rect 13044 24352 13050 24364
rect 13173 24361 13185 24364
rect 13219 24361 13231 24395
rect 13173 24355 13231 24361
rect 6273 24327 6331 24333
rect 6273 24324 6285 24327
rect 5368 24296 6285 24324
rect 4341 24191 4399 24197
rect 4341 24188 4353 24191
rect 3844 24160 4353 24188
rect 3844 24148 3850 24160
rect 4341 24157 4353 24160
rect 4387 24157 4399 24191
rect 4341 24151 4399 24157
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24188 4583 24191
rect 4798 24188 4804 24200
rect 4571 24160 4804 24188
rect 4571 24157 4583 24160
rect 4525 24151 4583 24157
rect 1857 24123 1915 24129
rect 1857 24089 1869 24123
rect 1903 24120 1915 24123
rect 2130 24120 2136 24132
rect 1903 24092 2136 24120
rect 1903 24089 1915 24092
rect 1857 24083 1915 24089
rect 2130 24080 2136 24092
rect 2188 24080 2194 24132
rect 4246 24080 4252 24132
rect 4304 24120 4310 24132
rect 4540 24120 4568 24151
rect 4798 24148 4804 24160
rect 4856 24148 4862 24200
rect 5166 24148 5172 24200
rect 5224 24148 5230 24200
rect 5368 24197 5396 24296
rect 6273 24293 6285 24296
rect 6319 24293 6331 24327
rect 6273 24287 6331 24293
rect 7009 24327 7067 24333
rect 7009 24293 7021 24327
rect 7055 24324 7067 24327
rect 7374 24324 7380 24336
rect 7055 24296 7380 24324
rect 7055 24293 7067 24296
rect 7009 24287 7067 24293
rect 7374 24284 7380 24296
rect 7432 24324 7438 24336
rect 8202 24324 8208 24336
rect 7432 24296 8208 24324
rect 7432 24284 7438 24296
rect 8202 24284 8208 24296
rect 8260 24284 8266 24336
rect 6178 24216 6184 24268
rect 6236 24256 6242 24268
rect 6236 24228 6684 24256
rect 6236 24216 6242 24228
rect 5353 24191 5411 24197
rect 5353 24157 5365 24191
rect 5399 24157 5411 24191
rect 5353 24151 5411 24157
rect 6086 24148 6092 24200
rect 6144 24148 6150 24200
rect 6454 24148 6460 24200
rect 6512 24190 6518 24200
rect 6656 24197 6684 24228
rect 7558 24216 7564 24268
rect 7616 24216 7622 24268
rect 7650 24216 7656 24268
rect 7708 24256 7714 24268
rect 13188 24256 13216 24355
rect 14734 24352 14740 24404
rect 14792 24392 14798 24404
rect 15013 24395 15071 24401
rect 15013 24392 15025 24395
rect 14792 24364 15025 24392
rect 14792 24352 14798 24364
rect 15013 24361 15025 24364
rect 15059 24361 15071 24395
rect 15013 24355 15071 24361
rect 13998 24284 14004 24336
rect 14056 24324 14062 24336
rect 14056 24296 14780 24324
rect 14056 24284 14062 24296
rect 13265 24259 13323 24265
rect 13265 24256 13277 24259
rect 7708 24228 9996 24256
rect 13188 24228 13277 24256
rect 7708 24216 7714 24228
rect 9968 24200 9996 24228
rect 13265 24225 13277 24228
rect 13311 24225 13323 24259
rect 13265 24219 13323 24225
rect 14090 24216 14096 24268
rect 14148 24256 14154 24268
rect 14645 24259 14703 24265
rect 14645 24256 14657 24259
rect 14148 24228 14657 24256
rect 14148 24216 14154 24228
rect 14645 24225 14657 24228
rect 14691 24225 14703 24259
rect 14645 24219 14703 24225
rect 6549 24191 6607 24197
rect 6549 24190 6561 24191
rect 6512 24162 6561 24190
rect 6512 24148 6518 24162
rect 6549 24157 6561 24162
rect 6595 24157 6607 24191
rect 6549 24151 6607 24157
rect 6641 24191 6699 24197
rect 6641 24157 6653 24191
rect 6687 24157 6699 24191
rect 6641 24151 6699 24157
rect 6822 24148 6828 24200
rect 6880 24148 6886 24200
rect 6917 24191 6975 24197
rect 6917 24157 6929 24191
rect 6963 24157 6975 24191
rect 6917 24151 6975 24157
rect 4304 24092 4568 24120
rect 4304 24080 4310 24092
rect 4614 24080 4620 24132
rect 4672 24120 4678 24132
rect 5261 24123 5319 24129
rect 5261 24120 5273 24123
rect 4672 24092 5273 24120
rect 4672 24080 4678 24092
rect 5261 24089 5273 24092
rect 5307 24089 5319 24123
rect 5261 24083 5319 24089
rect 5626 24080 5632 24132
rect 5684 24120 5690 24132
rect 6273 24123 6331 24129
rect 6273 24120 6285 24123
rect 5684 24092 6285 24120
rect 5684 24080 5690 24092
rect 6273 24089 6285 24092
rect 6319 24089 6331 24123
rect 6932 24120 6960 24151
rect 7098 24148 7104 24200
rect 7156 24148 7162 24200
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24188 7251 24191
rect 7466 24188 7472 24200
rect 7239 24160 7472 24188
rect 7239 24157 7251 24160
rect 7193 24151 7251 24157
rect 7208 24120 7236 24151
rect 7466 24148 7472 24160
rect 7524 24148 7530 24200
rect 8202 24148 8208 24200
rect 8260 24188 8266 24200
rect 8389 24191 8447 24197
rect 8389 24188 8401 24191
rect 8260 24160 8401 24188
rect 8260 24148 8266 24160
rect 8389 24157 8401 24160
rect 8435 24157 8447 24191
rect 8389 24151 8447 24157
rect 8481 24191 8539 24197
rect 8481 24157 8493 24191
rect 8527 24157 8539 24191
rect 8481 24151 8539 24157
rect 6932 24092 7236 24120
rect 7377 24123 7435 24129
rect 6273 24083 6331 24089
rect 7377 24089 7389 24123
rect 7423 24120 7435 24123
rect 7653 24123 7711 24129
rect 7423 24092 7604 24120
rect 7423 24089 7435 24092
rect 7377 24083 7435 24089
rect 7576 24064 7604 24092
rect 7653 24089 7665 24123
rect 7699 24120 7711 24123
rect 7742 24120 7748 24132
rect 7699 24092 7748 24120
rect 7699 24089 7711 24092
rect 7653 24083 7711 24089
rect 7742 24080 7748 24092
rect 7800 24080 7806 24132
rect 7834 24080 7840 24132
rect 7892 24129 7898 24132
rect 7892 24123 7911 24129
rect 7899 24089 7911 24123
rect 7892 24083 7911 24089
rect 7892 24080 7898 24083
rect 8018 24080 8024 24132
rect 8076 24120 8082 24132
rect 8496 24120 8524 24151
rect 8938 24148 8944 24200
rect 8996 24188 9002 24200
rect 9033 24191 9091 24197
rect 9033 24188 9045 24191
rect 8996 24160 9045 24188
rect 8996 24148 9002 24160
rect 9033 24157 9045 24160
rect 9079 24157 9091 24191
rect 9033 24151 9091 24157
rect 9214 24148 9220 24200
rect 9272 24148 9278 24200
rect 9306 24148 9312 24200
rect 9364 24148 9370 24200
rect 9490 24148 9496 24200
rect 9548 24148 9554 24200
rect 9582 24148 9588 24200
rect 9640 24148 9646 24200
rect 9677 24191 9735 24197
rect 9677 24157 9689 24191
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 8076 24092 8524 24120
rect 8665 24123 8723 24129
rect 8076 24080 8082 24092
rect 8665 24089 8677 24123
rect 8711 24120 8723 24123
rect 9122 24120 9128 24132
rect 8711 24092 9128 24120
rect 8711 24089 8723 24092
rect 8665 24083 8723 24089
rect 9122 24080 9128 24092
rect 9180 24120 9186 24132
rect 9692 24120 9720 24151
rect 9950 24148 9956 24200
rect 10008 24148 10014 24200
rect 11790 24148 11796 24200
rect 11848 24148 11854 24200
rect 12526 24148 12532 24200
rect 12584 24188 12590 24200
rect 14553 24191 14611 24197
rect 14553 24188 14565 24191
rect 12584 24160 14565 24188
rect 12584 24148 12590 24160
rect 14553 24157 14565 24160
rect 14599 24157 14611 24191
rect 14553 24151 14611 24157
rect 10198 24123 10256 24129
rect 10198 24120 10210 24123
rect 9180 24092 9720 24120
rect 9876 24092 10210 24120
rect 9180 24080 9186 24092
rect 2774 24012 2780 24064
rect 2832 24052 2838 24064
rect 3789 24055 3847 24061
rect 3789 24052 3801 24055
rect 2832 24024 3801 24052
rect 2832 24012 2838 24024
rect 3789 24021 3801 24024
rect 3835 24021 3847 24055
rect 3789 24015 3847 24021
rect 4154 24012 4160 24064
rect 4212 24052 4218 24064
rect 4706 24052 4712 24064
rect 4212 24024 4712 24052
rect 4212 24012 4218 24024
rect 4706 24012 4712 24024
rect 4764 24052 4770 24064
rect 4893 24055 4951 24061
rect 4893 24052 4905 24055
rect 4764 24024 4905 24052
rect 4764 24012 4770 24024
rect 4893 24021 4905 24024
rect 4939 24021 4951 24055
rect 4893 24015 4951 24021
rect 5074 24012 5080 24064
rect 5132 24052 5138 24064
rect 5442 24052 5448 24064
rect 5132 24024 5448 24052
rect 5132 24012 5138 24024
rect 5442 24012 5448 24024
rect 5500 24012 5506 24064
rect 6457 24055 6515 24061
rect 6457 24021 6469 24055
rect 6503 24052 6515 24055
rect 6914 24052 6920 24064
rect 6503 24024 6920 24052
rect 6503 24021 6515 24024
rect 6457 24015 6515 24021
rect 6914 24012 6920 24024
rect 6972 24052 6978 24064
rect 7098 24052 7104 24064
rect 6972 24024 7104 24052
rect 6972 24012 6978 24024
rect 7098 24012 7104 24024
rect 7156 24052 7162 24064
rect 7558 24052 7564 24064
rect 7156 24024 7564 24052
rect 7156 24012 7162 24024
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 8389 24055 8447 24061
rect 8389 24021 8401 24055
rect 8435 24052 8447 24055
rect 9398 24052 9404 24064
rect 8435 24024 9404 24052
rect 8435 24021 8447 24024
rect 8389 24015 8447 24021
rect 9398 24012 9404 24024
rect 9456 24012 9462 24064
rect 9876 24061 9904 24092
rect 10198 24089 10210 24092
rect 10244 24089 10256 24123
rect 10198 24083 10256 24089
rect 12060 24123 12118 24129
rect 12060 24089 12072 24123
rect 12106 24120 12118 24123
rect 13909 24123 13967 24129
rect 12106 24092 13308 24120
rect 12106 24089 12118 24092
rect 12060 24083 12118 24089
rect 9861 24055 9919 24061
rect 9861 24021 9873 24055
rect 9907 24021 9919 24055
rect 13280 24052 13308 24092
rect 13909 24089 13921 24123
rect 13955 24120 13967 24123
rect 14461 24123 14519 24129
rect 14461 24120 14473 24123
rect 13955 24092 14473 24120
rect 13955 24089 13967 24092
rect 13909 24083 13967 24089
rect 14461 24089 14473 24092
rect 14507 24089 14519 24123
rect 14461 24083 14519 24089
rect 14093 24055 14151 24061
rect 14093 24052 14105 24055
rect 13280 24024 14105 24052
rect 9861 24015 9919 24021
rect 14093 24021 14105 24024
rect 14139 24021 14151 24055
rect 14660 24052 14688 24219
rect 14752 24120 14780 24296
rect 14826 24148 14832 24200
rect 14884 24188 14890 24200
rect 14921 24191 14979 24197
rect 14921 24188 14933 24191
rect 14884 24160 14933 24188
rect 14884 24148 14890 24160
rect 14921 24157 14933 24160
rect 14967 24157 14979 24191
rect 15028 24188 15056 24355
rect 17954 24352 17960 24404
rect 18012 24392 18018 24404
rect 19150 24392 19156 24404
rect 18012 24364 19156 24392
rect 18012 24352 18018 24364
rect 19150 24352 19156 24364
rect 19208 24392 19214 24404
rect 19886 24392 19892 24404
rect 19208 24364 19892 24392
rect 19208 24352 19214 24364
rect 19886 24352 19892 24364
rect 19944 24352 19950 24404
rect 20349 24395 20407 24401
rect 20349 24361 20361 24395
rect 20395 24392 20407 24395
rect 20714 24392 20720 24404
rect 20395 24364 20720 24392
rect 20395 24361 20407 24364
rect 20349 24355 20407 24361
rect 20714 24352 20720 24364
rect 20772 24392 20778 24404
rect 22186 24392 22192 24404
rect 20772 24364 22192 24392
rect 20772 24352 20778 24364
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 25409 24395 25467 24401
rect 25409 24361 25421 24395
rect 25455 24392 25467 24395
rect 26329 24395 26387 24401
rect 26329 24392 26341 24395
rect 25455 24364 26341 24392
rect 25455 24361 25467 24364
rect 25409 24355 25467 24361
rect 26329 24361 26341 24364
rect 26375 24361 26387 24395
rect 26329 24355 26387 24361
rect 26605 24395 26663 24401
rect 26605 24361 26617 24395
rect 26651 24392 26663 24395
rect 26970 24392 26976 24404
rect 26651 24364 26976 24392
rect 26651 24361 26663 24364
rect 26605 24355 26663 24361
rect 26970 24352 26976 24364
rect 27028 24352 27034 24404
rect 27890 24352 27896 24404
rect 27948 24392 27954 24404
rect 28350 24392 28356 24404
rect 27948 24364 28356 24392
rect 27948 24352 27954 24364
rect 28350 24352 28356 24364
rect 28408 24392 28414 24404
rect 28810 24392 28816 24404
rect 28408 24364 28816 24392
rect 28408 24352 28414 24364
rect 28810 24352 28816 24364
rect 28868 24352 28874 24404
rect 29917 24395 29975 24401
rect 29917 24361 29929 24395
rect 29963 24361 29975 24395
rect 29917 24355 29975 24361
rect 30285 24395 30343 24401
rect 30285 24361 30297 24395
rect 30331 24392 30343 24395
rect 30374 24392 30380 24404
rect 30331 24364 30380 24392
rect 30331 24361 30343 24364
rect 30285 24355 30343 24361
rect 18322 24284 18328 24336
rect 18380 24324 18386 24336
rect 23937 24327 23995 24333
rect 18380 24296 19932 24324
rect 18380 24284 18386 24296
rect 16761 24259 16819 24265
rect 16761 24225 16773 24259
rect 16807 24256 16819 24259
rect 17034 24256 17040 24268
rect 16807 24228 17040 24256
rect 16807 24225 16819 24228
rect 16761 24219 16819 24225
rect 17034 24216 17040 24228
rect 17092 24256 17098 24268
rect 18138 24256 18144 24268
rect 17092 24228 18144 24256
rect 17092 24216 17098 24228
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 18598 24216 18604 24268
rect 18656 24256 18662 24268
rect 19518 24256 19524 24268
rect 18656 24228 19524 24256
rect 18656 24216 18662 24228
rect 15197 24191 15255 24197
rect 15197 24188 15209 24191
rect 15028 24160 15209 24188
rect 14921 24151 14979 24157
rect 15197 24157 15209 24160
rect 15243 24157 15255 24191
rect 15197 24151 15255 24157
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24157 15439 24191
rect 15381 24151 15439 24157
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 16942 24188 16948 24200
rect 16899 24160 16948 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 15396 24120 15424 24151
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 17218 24148 17224 24200
rect 17276 24148 17282 24200
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24188 18107 24191
rect 18506 24188 18512 24200
rect 18095 24160 18512 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 18708 24197 18736 24228
rect 19518 24216 19524 24228
rect 19576 24216 19582 24268
rect 18693 24191 18751 24197
rect 18693 24157 18705 24191
rect 18739 24157 18751 24191
rect 18693 24151 18751 24157
rect 18782 24148 18788 24200
rect 18840 24148 18846 24200
rect 18969 24191 19027 24197
rect 18969 24157 18981 24191
rect 19015 24157 19027 24191
rect 18969 24151 19027 24157
rect 14752 24092 15424 24120
rect 16666 24080 16672 24132
rect 16724 24120 16730 24132
rect 17129 24123 17187 24129
rect 17129 24120 17141 24123
rect 16724 24092 17141 24120
rect 16724 24080 16730 24092
rect 17129 24089 17141 24092
rect 17175 24089 17187 24123
rect 17129 24083 17187 24089
rect 18230 24080 18236 24132
rect 18288 24120 18294 24132
rect 18800 24120 18828 24148
rect 18288 24092 18828 24120
rect 18984 24120 19012 24151
rect 19058 24148 19064 24200
rect 19116 24188 19122 24200
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 19116 24160 19257 24188
rect 19116 24148 19122 24160
rect 19245 24157 19257 24160
rect 19291 24157 19303 24191
rect 19245 24151 19303 24157
rect 19426 24148 19432 24200
rect 19484 24148 19490 24200
rect 19702 24148 19708 24200
rect 19760 24148 19766 24200
rect 19904 24188 19932 24296
rect 23937 24293 23949 24327
rect 23983 24324 23995 24327
rect 24210 24324 24216 24336
rect 23983 24296 24216 24324
rect 23983 24293 23995 24296
rect 23937 24287 23995 24293
rect 24210 24284 24216 24296
rect 24268 24284 24274 24336
rect 25130 24284 25136 24336
rect 25188 24324 25194 24336
rect 25593 24327 25651 24333
rect 25593 24324 25605 24327
rect 25188 24296 25605 24324
rect 25188 24284 25194 24296
rect 25593 24293 25605 24296
rect 25639 24293 25651 24327
rect 25593 24287 25651 24293
rect 28626 24284 28632 24336
rect 28684 24324 28690 24336
rect 29638 24324 29644 24336
rect 28684 24296 29644 24324
rect 28684 24284 28690 24296
rect 29638 24284 29644 24296
rect 29696 24324 29702 24336
rect 29932 24324 29960 24355
rect 30374 24352 30380 24364
rect 30432 24352 30438 24404
rect 30558 24352 30564 24404
rect 30616 24392 30622 24404
rect 30745 24395 30803 24401
rect 30745 24392 30757 24395
rect 30616 24364 30757 24392
rect 30616 24352 30622 24364
rect 30745 24361 30757 24364
rect 30791 24361 30803 24395
rect 30745 24355 30803 24361
rect 30834 24352 30840 24404
rect 30892 24392 30898 24404
rect 30929 24395 30987 24401
rect 30929 24392 30941 24395
rect 30892 24364 30941 24392
rect 30892 24352 30898 24364
rect 30929 24361 30941 24364
rect 30975 24361 30987 24395
rect 31662 24392 31668 24404
rect 30929 24355 30987 24361
rect 31588 24364 31668 24392
rect 29696 24296 29960 24324
rect 30101 24327 30159 24333
rect 29696 24284 29702 24296
rect 30101 24293 30113 24327
rect 30147 24324 30159 24327
rect 31588 24324 31616 24364
rect 31662 24352 31668 24364
rect 31720 24352 31726 24404
rect 32950 24352 32956 24404
rect 33008 24352 33014 24404
rect 33134 24352 33140 24404
rect 33192 24392 33198 24404
rect 33594 24392 33600 24404
rect 33192 24364 33600 24392
rect 33192 24352 33198 24364
rect 33594 24352 33600 24364
rect 33652 24352 33658 24404
rect 34606 24352 34612 24404
rect 34664 24392 34670 24404
rect 38654 24392 38660 24404
rect 34664 24364 38660 24392
rect 34664 24352 34670 24364
rect 38654 24352 38660 24364
rect 38712 24352 38718 24404
rect 41322 24352 41328 24404
rect 41380 24392 41386 24404
rect 42153 24395 42211 24401
rect 42153 24392 42165 24395
rect 41380 24364 42165 24392
rect 41380 24352 41386 24364
rect 42153 24361 42165 24364
rect 42199 24361 42211 24395
rect 42153 24355 42211 24361
rect 33502 24324 33508 24336
rect 30147 24296 31616 24324
rect 32416 24296 33508 24324
rect 30147 24293 30159 24296
rect 30101 24287 30159 24293
rect 19978 24216 19984 24268
rect 20036 24256 20042 24268
rect 20165 24259 20223 24265
rect 20165 24256 20177 24259
rect 20036 24228 20177 24256
rect 20036 24216 20042 24228
rect 20165 24225 20177 24228
rect 20211 24225 20223 24259
rect 20165 24219 20223 24225
rect 21818 24216 21824 24268
rect 21876 24216 21882 24268
rect 22097 24259 22155 24265
rect 22097 24225 22109 24259
rect 22143 24256 22155 24259
rect 22189 24259 22247 24265
rect 22189 24256 22201 24259
rect 22143 24228 22201 24256
rect 22143 24225 22155 24228
rect 22097 24219 22155 24225
rect 22189 24225 22201 24228
rect 22235 24256 22247 24259
rect 23474 24256 23480 24268
rect 22235 24228 23480 24256
rect 22235 24225 22247 24228
rect 22189 24219 22247 24225
rect 23474 24216 23480 24228
rect 23532 24216 23538 24268
rect 24670 24216 24676 24268
rect 24728 24256 24734 24268
rect 25774 24256 25780 24268
rect 24728 24228 25780 24256
rect 24728 24216 24734 24228
rect 25774 24216 25780 24228
rect 25832 24216 25838 24268
rect 26881 24259 26939 24265
rect 26068 24228 26648 24256
rect 26068 24200 26096 24228
rect 19904 24160 20070 24188
rect 19797 24123 19855 24129
rect 18984 24092 19380 24120
rect 18288 24080 18294 24092
rect 19352 24064 19380 24092
rect 19797 24089 19809 24123
rect 19843 24089 19855 24123
rect 19797 24083 19855 24089
rect 15289 24055 15347 24061
rect 15289 24052 15301 24055
rect 14660 24024 15301 24052
rect 14093 24015 14151 24021
rect 15289 24021 15301 24024
rect 15335 24021 15347 24055
rect 15289 24015 15347 24021
rect 16390 24012 16396 24064
rect 16448 24052 16454 24064
rect 16577 24055 16635 24061
rect 16577 24052 16589 24055
rect 16448 24024 16589 24052
rect 16448 24012 16454 24024
rect 16577 24021 16589 24024
rect 16623 24021 16635 24055
rect 16577 24015 16635 24021
rect 16758 24012 16764 24064
rect 16816 24052 16822 24064
rect 16945 24055 17003 24061
rect 16945 24052 16957 24055
rect 16816 24024 16957 24052
rect 16816 24012 16822 24024
rect 16945 24021 16957 24024
rect 16991 24021 17003 24055
rect 16945 24015 17003 24021
rect 18414 24012 18420 24064
rect 18472 24012 18478 24064
rect 18509 24055 18567 24061
rect 18509 24021 18521 24055
rect 18555 24052 18567 24055
rect 18782 24052 18788 24064
rect 18555 24024 18788 24052
rect 18555 24021 18567 24024
rect 18509 24015 18567 24021
rect 18782 24012 18788 24024
rect 18840 24012 18846 24064
rect 18877 24055 18935 24061
rect 18877 24021 18889 24055
rect 18923 24052 18935 24055
rect 19150 24052 19156 24064
rect 18923 24024 19156 24052
rect 18923 24021 18935 24024
rect 18877 24015 18935 24021
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 19334 24012 19340 24064
rect 19392 24012 19398 24064
rect 19518 24012 19524 24064
rect 19576 24012 19582 24064
rect 19812 24052 19840 24083
rect 19886 24080 19892 24132
rect 19944 24080 19950 24132
rect 20042 24129 20070 24160
rect 24578 24148 24584 24200
rect 24636 24148 24642 24200
rect 24854 24148 24860 24200
rect 24912 24148 24918 24200
rect 24946 24148 24952 24200
rect 25004 24148 25010 24200
rect 25130 24148 25136 24200
rect 25188 24148 25194 24200
rect 25222 24148 25228 24200
rect 25280 24148 25286 24200
rect 25501 24191 25559 24197
rect 25501 24157 25513 24191
rect 25547 24188 25559 24191
rect 25682 24188 25688 24200
rect 25547 24160 25688 24188
rect 25547 24157 25559 24160
rect 25501 24151 25559 24157
rect 25682 24148 25688 24160
rect 25740 24148 25746 24200
rect 25869 24191 25927 24197
rect 25869 24157 25881 24191
rect 25915 24188 25927 24191
rect 26050 24188 26056 24200
rect 25915 24160 26056 24188
rect 25915 24157 25927 24160
rect 25869 24151 25927 24157
rect 26050 24148 26056 24160
rect 26108 24148 26114 24200
rect 26234 24148 26240 24200
rect 26292 24148 26298 24200
rect 26329 24191 26387 24197
rect 26329 24157 26341 24191
rect 26375 24157 26387 24191
rect 26329 24151 26387 24157
rect 20027 24123 20085 24129
rect 20027 24089 20039 24123
rect 20073 24120 20085 24123
rect 20438 24120 20444 24132
rect 20073 24092 20444 24120
rect 20073 24089 20085 24092
rect 20027 24083 20085 24089
rect 20438 24080 20444 24092
rect 20496 24080 20502 24132
rect 21910 24120 21916 24132
rect 21390 24092 21916 24120
rect 21910 24080 21916 24092
rect 21968 24080 21974 24132
rect 22462 24080 22468 24132
rect 22520 24080 22526 24132
rect 24673 24123 24731 24129
rect 23690 24092 24624 24120
rect 24596 24064 24624 24092
rect 24673 24089 24685 24123
rect 24719 24120 24731 24123
rect 25590 24120 25596 24132
rect 24719 24092 25596 24120
rect 24719 24089 24731 24092
rect 24673 24083 24731 24089
rect 25590 24080 25596 24092
rect 25648 24120 25654 24132
rect 26142 24120 26148 24132
rect 25648 24092 26148 24120
rect 25648 24080 25654 24092
rect 26142 24080 26148 24092
rect 26200 24080 26206 24132
rect 20254 24052 20260 24064
rect 19812 24024 20260 24052
rect 20254 24012 20260 24024
rect 20312 24012 20318 24064
rect 24578 24012 24584 24064
rect 24636 24012 24642 24064
rect 24758 24055 24816 24061
rect 24758 24021 24770 24055
rect 24804 24052 24816 24055
rect 26344 24052 26372 24151
rect 26510 24148 26516 24200
rect 26568 24148 26574 24200
rect 26620 24197 26648 24228
rect 26881 24225 26893 24259
rect 26927 24256 26939 24259
rect 27614 24256 27620 24268
rect 26927 24228 27620 24256
rect 26927 24225 26939 24228
rect 26881 24219 26939 24225
rect 27614 24216 27620 24228
rect 27672 24216 27678 24268
rect 28166 24216 28172 24268
rect 28224 24256 28230 24268
rect 32416 24256 32444 24296
rect 33502 24284 33508 24296
rect 33560 24324 33566 24336
rect 36446 24324 36452 24336
rect 33560 24296 36452 24324
rect 33560 24284 33566 24296
rect 28224 24228 32444 24256
rect 32493 24259 32551 24265
rect 28224 24216 28230 24228
rect 32493 24225 32505 24259
rect 32539 24225 32551 24259
rect 32950 24256 32956 24268
rect 32493 24219 32551 24225
rect 32600 24228 32956 24256
rect 26605 24191 26663 24197
rect 26605 24157 26617 24191
rect 26651 24157 26663 24191
rect 26605 24151 26663 24157
rect 26786 24148 26792 24200
rect 26844 24148 26850 24200
rect 28442 24188 28448 24200
rect 28290 24160 28448 24188
rect 28442 24148 28448 24160
rect 28500 24148 28506 24200
rect 28552 24160 30420 24188
rect 24804 24024 26372 24052
rect 26528 24052 26556 24148
rect 27154 24080 27160 24132
rect 27212 24080 27218 24132
rect 28552 24052 28580 24160
rect 29733 24123 29791 24129
rect 29733 24089 29745 24123
rect 29779 24089 29791 24123
rect 29733 24083 29791 24089
rect 26528 24024 28580 24052
rect 28629 24055 28687 24061
rect 24804 24021 24816 24024
rect 24758 24015 24816 24021
rect 28629 24021 28641 24055
rect 28675 24052 28687 24055
rect 28810 24052 28816 24064
rect 28675 24024 28816 24052
rect 28675 24021 28687 24024
rect 28629 24015 28687 24021
rect 28810 24012 28816 24024
rect 28868 24012 28874 24064
rect 29748 24052 29776 24083
rect 29822 24080 29828 24132
rect 29880 24120 29886 24132
rect 29933 24123 29991 24129
rect 29933 24120 29945 24123
rect 29880 24092 29945 24120
rect 29880 24080 29886 24092
rect 29933 24089 29945 24092
rect 29979 24089 29991 24123
rect 30392 24120 30420 24160
rect 30466 24148 30472 24200
rect 30524 24148 30530 24200
rect 30561 24191 30619 24197
rect 30561 24157 30573 24191
rect 30607 24188 30619 24191
rect 30650 24188 30656 24200
rect 30607 24160 30656 24188
rect 30607 24157 30619 24160
rect 30561 24151 30619 24157
rect 30650 24148 30656 24160
rect 30708 24148 30714 24200
rect 30834 24148 30840 24200
rect 30892 24188 30898 24200
rect 31202 24188 31208 24200
rect 30892 24160 31208 24188
rect 30892 24148 30898 24160
rect 31202 24148 31208 24160
rect 31260 24148 31266 24200
rect 31386 24148 31392 24200
rect 31444 24188 31450 24200
rect 31846 24188 31852 24200
rect 31444 24160 31852 24188
rect 31444 24148 31450 24160
rect 31846 24148 31852 24160
rect 31904 24148 31910 24200
rect 30926 24120 30932 24132
rect 30392 24092 30932 24120
rect 29933 24083 29991 24089
rect 30926 24080 30932 24092
rect 30984 24080 30990 24132
rect 31018 24080 31024 24132
rect 31076 24120 31082 24132
rect 31113 24123 31171 24129
rect 31113 24120 31125 24123
rect 31076 24092 31125 24120
rect 31076 24080 31082 24092
rect 31113 24089 31125 24092
rect 31159 24089 31171 24123
rect 31113 24083 31171 24089
rect 31297 24123 31355 24129
rect 31297 24089 31309 24123
rect 31343 24120 31355 24123
rect 31662 24120 31668 24132
rect 31343 24092 31668 24120
rect 31343 24089 31355 24092
rect 31297 24083 31355 24089
rect 30834 24052 30840 24064
rect 29748 24024 30840 24052
rect 30834 24012 30840 24024
rect 30892 24012 30898 24064
rect 31128 24052 31156 24083
rect 31662 24080 31668 24092
rect 31720 24120 31726 24132
rect 32508 24120 32536 24219
rect 32600 24197 32628 24228
rect 32950 24216 32956 24228
rect 33008 24216 33014 24268
rect 33042 24216 33048 24268
rect 33100 24256 33106 24268
rect 35894 24256 35900 24268
rect 33100 24228 35900 24256
rect 33100 24216 33106 24228
rect 35894 24216 35900 24228
rect 35952 24216 35958 24268
rect 35986 24216 35992 24268
rect 36044 24216 36050 24268
rect 36280 24265 36308 24296
rect 36446 24284 36452 24296
rect 36504 24284 36510 24336
rect 36265 24259 36323 24265
rect 36265 24225 36277 24259
rect 36311 24225 36323 24259
rect 36265 24219 36323 24225
rect 36998 24216 37004 24268
rect 37056 24216 37062 24268
rect 37274 24216 37280 24268
rect 37332 24216 37338 24268
rect 38746 24216 38752 24268
rect 38804 24256 38810 24268
rect 39025 24259 39083 24265
rect 39025 24256 39037 24259
rect 38804 24228 39037 24256
rect 38804 24216 38810 24228
rect 39025 24225 39037 24228
rect 39071 24256 39083 24259
rect 39758 24256 39764 24268
rect 39071 24228 39764 24256
rect 39071 24225 39083 24228
rect 39025 24219 39083 24225
rect 39758 24216 39764 24228
rect 39816 24216 39822 24268
rect 40681 24259 40739 24265
rect 40681 24225 40693 24259
rect 40727 24256 40739 24259
rect 40770 24256 40776 24268
rect 40727 24228 40776 24256
rect 40727 24225 40739 24228
rect 40681 24219 40739 24225
rect 40770 24216 40776 24228
rect 40828 24216 40834 24268
rect 32585 24191 32643 24197
rect 32585 24157 32597 24191
rect 32631 24157 32643 24191
rect 32585 24151 32643 24157
rect 32674 24148 32680 24200
rect 32732 24188 32738 24200
rect 34606 24188 34612 24200
rect 32732 24160 34612 24188
rect 32732 24148 32738 24160
rect 34606 24148 34612 24160
rect 34664 24148 34670 24200
rect 34701 24191 34759 24197
rect 34701 24157 34713 24191
rect 34747 24188 34759 24191
rect 34974 24188 34980 24200
rect 34747 24160 34980 24188
rect 34747 24157 34759 24160
rect 34701 24151 34759 24157
rect 34974 24148 34980 24160
rect 35032 24188 35038 24200
rect 35529 24191 35587 24197
rect 35529 24188 35541 24191
rect 35032 24160 35541 24188
rect 35032 24148 35038 24160
rect 35529 24157 35541 24160
rect 35575 24157 35587 24191
rect 35529 24151 35587 24157
rect 35618 24148 35624 24200
rect 35676 24148 35682 24200
rect 36004 24188 36032 24216
rect 39574 24188 39580 24200
rect 35912 24160 36584 24188
rect 38410 24160 39580 24188
rect 34790 24120 34796 24132
rect 31720 24092 34796 24120
rect 31720 24080 31726 24092
rect 34790 24080 34796 24092
rect 34848 24120 34854 24132
rect 34885 24123 34943 24129
rect 34885 24120 34897 24123
rect 34848 24092 34897 24120
rect 34848 24080 34854 24092
rect 34885 24089 34897 24092
rect 34931 24089 34943 24123
rect 34885 24083 34943 24089
rect 35069 24123 35127 24129
rect 35069 24089 35081 24123
rect 35115 24120 35127 24123
rect 35158 24120 35164 24132
rect 35115 24092 35164 24120
rect 35115 24089 35127 24092
rect 35069 24083 35127 24089
rect 35158 24080 35164 24092
rect 35216 24080 35222 24132
rect 35253 24123 35311 24129
rect 35253 24089 35265 24123
rect 35299 24120 35311 24123
rect 35912 24120 35940 24160
rect 35299 24092 35940 24120
rect 35989 24123 36047 24129
rect 35299 24089 35311 24092
rect 35253 24083 35311 24089
rect 35989 24089 36001 24123
rect 36035 24120 36047 24123
rect 36078 24120 36084 24132
rect 36035 24092 36084 24120
rect 36035 24089 36047 24092
rect 35989 24083 36047 24089
rect 36078 24080 36084 24092
rect 36136 24080 36142 24132
rect 36556 24120 36584 24160
rect 39574 24148 39580 24160
rect 39632 24148 39638 24200
rect 40034 24148 40040 24200
rect 40092 24148 40098 24200
rect 40402 24148 40408 24200
rect 40460 24148 40466 24200
rect 41782 24148 41788 24200
rect 41840 24148 41846 24200
rect 36556 24092 37688 24120
rect 31478 24052 31484 24064
rect 31128 24024 31484 24052
rect 31478 24012 31484 24024
rect 31536 24012 31542 24064
rect 32490 24012 32496 24064
rect 32548 24052 32554 24064
rect 32950 24052 32956 24064
rect 32548 24024 32956 24052
rect 32548 24012 32554 24024
rect 32950 24012 32956 24024
rect 33008 24052 33014 24064
rect 34514 24052 34520 24064
rect 33008 24024 34520 24052
rect 33008 24012 33014 24024
rect 34514 24012 34520 24024
rect 34572 24052 34578 24064
rect 36556 24061 36584 24092
rect 34977 24055 35035 24061
rect 34977 24052 34989 24055
rect 34572 24024 34989 24052
rect 34572 24012 34578 24024
rect 34977 24021 34989 24024
rect 35023 24021 35035 24055
rect 34977 24015 35035 24021
rect 35345 24055 35403 24061
rect 35345 24021 35357 24055
rect 35391 24052 35403 24055
rect 36449 24055 36507 24061
rect 36449 24052 36461 24055
rect 35391 24024 36461 24052
rect 35391 24021 35403 24024
rect 35345 24015 35403 24021
rect 36449 24021 36461 24024
rect 36495 24021 36507 24055
rect 36449 24015 36507 24021
rect 36541 24055 36599 24061
rect 36541 24021 36553 24055
rect 36587 24052 36599 24055
rect 36722 24052 36728 24064
rect 36587 24024 36728 24052
rect 36587 24021 36599 24024
rect 36541 24015 36599 24021
rect 36722 24012 36728 24024
rect 36780 24012 36786 24064
rect 36909 24055 36967 24061
rect 36909 24021 36921 24055
rect 36955 24052 36967 24055
rect 37550 24052 37556 24064
rect 36955 24024 37556 24052
rect 36955 24021 36967 24024
rect 36909 24015 36967 24021
rect 37550 24012 37556 24024
rect 37608 24012 37614 24064
rect 37660 24052 37688 24092
rect 39298 24080 39304 24132
rect 39356 24080 39362 24132
rect 39482 24080 39488 24132
rect 39540 24080 39546 24132
rect 40678 24120 40684 24132
rect 39592 24092 40684 24120
rect 39022 24052 39028 24064
rect 37660 24024 39028 24052
rect 39022 24012 39028 24024
rect 39080 24052 39086 24064
rect 39592 24052 39620 24092
rect 40678 24080 40684 24092
rect 40736 24080 40742 24132
rect 39080 24024 39620 24052
rect 39669 24055 39727 24061
rect 39080 24012 39086 24024
rect 39669 24021 39681 24055
rect 39715 24052 39727 24055
rect 39758 24052 39764 24064
rect 39715 24024 39764 24052
rect 39715 24021 39727 24024
rect 39669 24015 39727 24021
rect 39758 24012 39764 24024
rect 39816 24012 39822 24064
rect 40218 24012 40224 24064
rect 40276 24012 40282 24064
rect 1104 23962 42504 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 42504 23962
rect 1104 23888 42504 23910
rect 2317 23851 2375 23857
rect 2317 23817 2329 23851
rect 2363 23848 2375 23851
rect 2363 23820 2728 23848
rect 2363 23817 2375 23820
rect 2317 23811 2375 23817
rect 2700 23792 2728 23820
rect 3970 23808 3976 23860
rect 4028 23808 4034 23860
rect 7742 23848 7748 23860
rect 7208 23820 7748 23848
rect 2133 23783 2191 23789
rect 2133 23749 2145 23783
rect 2179 23780 2191 23783
rect 2498 23780 2504 23792
rect 2179 23752 2504 23780
rect 2179 23749 2191 23752
rect 2133 23743 2191 23749
rect 2498 23740 2504 23752
rect 2556 23740 2562 23792
rect 2682 23740 2688 23792
rect 2740 23780 2746 23792
rect 2740 23752 3740 23780
rect 2740 23740 2746 23752
rect 1394 23672 1400 23724
rect 1452 23672 1458 23724
rect 2409 23715 2467 23721
rect 2409 23681 2421 23715
rect 2455 23712 2467 23715
rect 2774 23712 2780 23724
rect 2455 23684 2780 23712
rect 2455 23681 2467 23684
rect 2409 23675 2467 23681
rect 2774 23672 2780 23684
rect 2832 23672 2838 23724
rect 3712 23721 3740 23752
rect 3697 23715 3755 23721
rect 3697 23681 3709 23715
rect 3743 23681 3755 23715
rect 3697 23675 3755 23681
rect 3605 23647 3663 23653
rect 3605 23613 3617 23647
rect 3651 23613 3663 23647
rect 3712 23644 3740 23675
rect 3786 23672 3792 23724
rect 3844 23672 3850 23724
rect 3988 23712 4016 23808
rect 4614 23740 4620 23792
rect 4672 23740 4678 23792
rect 7208 23724 7236 23820
rect 7742 23808 7748 23820
rect 7800 23808 7806 23860
rect 8938 23808 8944 23860
rect 8996 23848 9002 23860
rect 12986 23848 12992 23860
rect 8996 23820 9536 23848
rect 8996 23808 9002 23820
rect 7282 23740 7288 23792
rect 7340 23780 7346 23792
rect 9508 23789 9536 23820
rect 9692 23820 12992 23848
rect 9493 23783 9551 23789
rect 7340 23752 7512 23780
rect 7340 23740 7346 23752
rect 4065 23715 4123 23721
rect 4065 23712 4077 23715
rect 3988 23684 4077 23712
rect 4065 23681 4077 23684
rect 4111 23681 4123 23715
rect 4065 23675 4123 23681
rect 5718 23672 5724 23724
rect 5776 23672 5782 23724
rect 6546 23672 6552 23724
rect 6604 23712 6610 23724
rect 6641 23715 6699 23721
rect 6641 23712 6653 23715
rect 6604 23684 6653 23712
rect 6604 23672 6610 23684
rect 6641 23681 6653 23684
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 7190 23672 7196 23724
rect 7248 23672 7254 23724
rect 7374 23672 7380 23724
rect 7432 23672 7438 23724
rect 7484 23721 7512 23752
rect 9493 23749 9505 23783
rect 9539 23749 9551 23783
rect 9493 23743 9551 23749
rect 7469 23715 7527 23721
rect 7469 23681 7481 23715
rect 7515 23681 7527 23715
rect 7469 23675 7527 23681
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23712 7619 23715
rect 7650 23712 7656 23724
rect 7607 23684 7656 23712
rect 7607 23681 7619 23684
rect 7561 23675 7619 23681
rect 4246 23644 4252 23656
rect 3712 23616 4252 23644
rect 3605 23607 3663 23613
rect 2130 23536 2136 23588
rect 2188 23536 2194 23588
rect 3620 23576 3648 23607
rect 4246 23604 4252 23616
rect 4304 23604 4310 23656
rect 4341 23647 4399 23653
rect 4341 23613 4353 23647
rect 4387 23644 4399 23647
rect 5994 23644 6000 23656
rect 4387 23616 6000 23644
rect 4387 23613 4399 23616
rect 4341 23607 4399 23613
rect 5994 23604 6000 23616
rect 6052 23604 6058 23656
rect 6089 23647 6147 23653
rect 6089 23613 6101 23647
rect 6135 23644 6147 23647
rect 7576 23644 7604 23675
rect 7650 23672 7656 23684
rect 7708 23672 7714 23724
rect 8849 23715 8907 23721
rect 8849 23681 8861 23715
rect 8895 23712 8907 23715
rect 9030 23712 9036 23724
rect 8895 23684 9036 23712
rect 8895 23681 8907 23684
rect 8849 23675 8907 23681
rect 6135 23616 7604 23644
rect 6135 23613 6147 23616
rect 6089 23607 6147 23613
rect 4154 23576 4160 23588
rect 3620 23548 4160 23576
rect 4154 23536 4160 23548
rect 4212 23536 4218 23588
rect 6822 23536 6828 23588
rect 6880 23576 6886 23588
rect 8864 23576 8892 23675
rect 9030 23672 9036 23684
rect 9088 23672 9094 23724
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23712 9367 23715
rect 9398 23712 9404 23724
rect 9355 23684 9404 23712
rect 9355 23681 9367 23684
rect 9309 23675 9367 23681
rect 9398 23672 9404 23684
rect 9456 23672 9462 23724
rect 9692 23721 9720 23820
rect 12986 23808 12992 23820
rect 13044 23808 13050 23860
rect 13078 23808 13084 23860
rect 13136 23848 13142 23860
rect 13357 23851 13415 23857
rect 13357 23848 13369 23851
rect 13136 23820 13369 23848
rect 13136 23808 13142 23820
rect 13357 23817 13369 23820
rect 13403 23848 13415 23851
rect 18046 23848 18052 23860
rect 13403 23820 14412 23848
rect 13403 23817 13415 23820
rect 13357 23811 13415 23817
rect 10226 23789 10232 23792
rect 10220 23780 10232 23789
rect 10187 23752 10232 23780
rect 10220 23743 10232 23752
rect 10226 23740 10232 23743
rect 10284 23740 10290 23792
rect 14274 23780 14280 23792
rect 11992 23752 14280 23780
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23681 9643 23715
rect 9585 23675 9643 23681
rect 9677 23715 9735 23721
rect 9677 23681 9689 23715
rect 9723 23681 9735 23715
rect 9677 23675 9735 23681
rect 9600 23644 9628 23675
rect 9950 23672 9956 23724
rect 10008 23672 10014 23724
rect 11790 23672 11796 23724
rect 11848 23712 11854 23724
rect 11992 23721 12020 23752
rect 14274 23740 14280 23752
rect 14332 23740 14338 23792
rect 11977 23715 12035 23721
rect 11977 23712 11989 23715
rect 11848 23684 11989 23712
rect 11848 23672 11854 23684
rect 11977 23681 11989 23684
rect 12023 23681 12035 23715
rect 11977 23675 12035 23681
rect 12244 23715 12302 23721
rect 12244 23681 12256 23715
rect 12290 23712 12302 23715
rect 13817 23715 13875 23721
rect 12290 23684 13492 23712
rect 12290 23681 12302 23684
rect 12244 23675 12302 23681
rect 9858 23644 9864 23656
rect 9600 23616 9864 23644
rect 9858 23604 9864 23616
rect 9916 23604 9922 23656
rect 13262 23576 13268 23588
rect 6880 23548 8892 23576
rect 12912 23548 13268 23576
rect 6880 23536 6886 23548
rect 1578 23468 1584 23520
rect 1636 23468 1642 23520
rect 4249 23511 4307 23517
rect 4249 23477 4261 23511
rect 4295 23508 4307 23511
rect 5810 23508 5816 23520
rect 4295 23480 5816 23508
rect 4295 23477 4307 23480
rect 4249 23471 4307 23477
rect 5810 23468 5816 23480
rect 5868 23468 5874 23520
rect 6457 23511 6515 23517
rect 6457 23477 6469 23511
rect 6503 23508 6515 23511
rect 7190 23508 7196 23520
rect 6503 23480 7196 23508
rect 6503 23477 6515 23480
rect 6457 23471 6515 23477
rect 7190 23468 7196 23480
rect 7248 23468 7254 23520
rect 7282 23468 7288 23520
rect 7340 23508 7346 23520
rect 7837 23511 7895 23517
rect 7837 23508 7849 23511
rect 7340 23480 7849 23508
rect 7340 23468 7346 23480
rect 7837 23477 7849 23480
rect 7883 23477 7895 23511
rect 7837 23471 7895 23477
rect 9861 23511 9919 23517
rect 9861 23477 9873 23511
rect 9907 23508 9919 23511
rect 10226 23508 10232 23520
rect 9907 23480 10232 23508
rect 9907 23477 9919 23480
rect 9861 23471 9919 23477
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 10318 23468 10324 23520
rect 10376 23508 10382 23520
rect 11333 23511 11391 23517
rect 11333 23508 11345 23511
rect 10376 23480 11345 23508
rect 10376 23468 10382 23480
rect 11333 23477 11345 23480
rect 11379 23508 11391 23511
rect 12912 23508 12940 23548
rect 13262 23536 13268 23548
rect 13320 23536 13326 23588
rect 13464 23585 13492 23684
rect 13817 23681 13829 23715
rect 13863 23712 13875 23715
rect 14384 23712 14412 23820
rect 17788 23820 18052 23848
rect 17788 23789 17816 23820
rect 18046 23808 18052 23820
rect 18104 23808 18110 23860
rect 18414 23808 18420 23860
rect 18472 23848 18478 23860
rect 18472 23820 18644 23848
rect 18472 23808 18478 23820
rect 18616 23789 18644 23820
rect 19702 23808 19708 23860
rect 19760 23848 19766 23860
rect 19889 23851 19947 23857
rect 19889 23848 19901 23851
rect 19760 23820 19901 23848
rect 19760 23808 19766 23820
rect 19889 23817 19901 23820
rect 19935 23817 19947 23851
rect 19889 23811 19947 23817
rect 20254 23808 20260 23860
rect 20312 23848 20318 23860
rect 20349 23851 20407 23857
rect 20349 23848 20361 23851
rect 20312 23820 20361 23848
rect 20312 23808 20318 23820
rect 20349 23817 20361 23820
rect 20395 23817 20407 23851
rect 20349 23811 20407 23817
rect 20438 23808 20444 23860
rect 20496 23848 20502 23860
rect 21910 23848 21916 23860
rect 20496 23820 21916 23848
rect 20496 23808 20502 23820
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 22462 23808 22468 23860
rect 22520 23848 22526 23860
rect 22649 23851 22707 23857
rect 22649 23848 22661 23851
rect 22520 23820 22661 23848
rect 22520 23808 22526 23820
rect 22649 23817 22661 23820
rect 22695 23817 22707 23851
rect 22649 23811 22707 23817
rect 23014 23808 23020 23860
rect 23072 23848 23078 23860
rect 23109 23851 23167 23857
rect 23109 23848 23121 23851
rect 23072 23820 23121 23848
rect 23072 23808 23078 23820
rect 23109 23817 23121 23820
rect 23155 23817 23167 23851
rect 24946 23848 24952 23860
rect 23109 23811 23167 23817
rect 24596 23820 24952 23848
rect 17773 23783 17831 23789
rect 17773 23749 17785 23783
rect 17819 23749 17831 23783
rect 17773 23743 17831 23749
rect 18601 23783 18659 23789
rect 18601 23749 18613 23783
rect 18647 23749 18659 23783
rect 18601 23743 18659 23749
rect 19426 23740 19432 23792
rect 19484 23780 19490 23792
rect 19794 23780 19800 23792
rect 19484 23752 19800 23780
rect 19484 23740 19490 23752
rect 19794 23740 19800 23752
rect 19852 23740 19858 23792
rect 20162 23740 20168 23792
rect 20220 23780 20226 23792
rect 20220 23752 20668 23780
rect 20220 23740 20226 23752
rect 14829 23715 14887 23721
rect 14829 23712 14841 23715
rect 13863 23684 14320 23712
rect 14384 23684 14841 23712
rect 13863 23681 13875 23684
rect 13817 23675 13875 23681
rect 13906 23604 13912 23656
rect 13964 23604 13970 23656
rect 13998 23604 14004 23656
rect 14056 23604 14062 23656
rect 14292 23653 14320 23684
rect 14829 23681 14841 23684
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 16209 23715 16267 23721
rect 16209 23681 16221 23715
rect 16255 23681 16267 23715
rect 16209 23675 16267 23681
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23613 14335 23647
rect 14277 23607 14335 23613
rect 13449 23579 13507 23585
rect 13449 23545 13461 23579
rect 13495 23545 13507 23579
rect 16224 23576 16252 23675
rect 16390 23672 16396 23724
rect 16448 23672 16454 23724
rect 16485 23715 16543 23721
rect 16485 23681 16497 23715
rect 16531 23712 16543 23715
rect 16574 23712 16580 23724
rect 16531 23684 16580 23712
rect 16531 23681 16543 23684
rect 16485 23675 16543 23681
rect 16574 23672 16580 23684
rect 16632 23712 16638 23724
rect 17034 23712 17040 23724
rect 16632 23684 17040 23712
rect 16632 23672 16638 23684
rect 17034 23672 17040 23684
rect 17092 23672 17098 23724
rect 17586 23672 17592 23724
rect 17644 23721 17650 23724
rect 17644 23715 17693 23721
rect 17644 23681 17647 23715
rect 17681 23681 17693 23715
rect 17644 23675 17693 23681
rect 17865 23715 17923 23721
rect 17865 23681 17877 23715
rect 17911 23681 17923 23715
rect 17865 23675 17923 23681
rect 17644 23672 17650 23675
rect 17126 23604 17132 23656
rect 17184 23604 17190 23656
rect 17405 23647 17463 23653
rect 17405 23613 17417 23647
rect 17451 23644 17463 23647
rect 17880 23644 17908 23675
rect 17954 23672 17960 23724
rect 18012 23721 18018 23724
rect 18012 23715 18051 23721
rect 18039 23681 18051 23715
rect 18012 23675 18051 23681
rect 18141 23715 18199 23721
rect 18141 23681 18153 23715
rect 18187 23681 18199 23715
rect 18141 23675 18199 23681
rect 18012 23672 18018 23675
rect 17451 23616 17908 23644
rect 18156 23644 18184 23675
rect 18322 23672 18328 23724
rect 18380 23712 18386 23724
rect 18417 23715 18475 23721
rect 18417 23712 18429 23715
rect 18380 23684 18429 23712
rect 18380 23672 18386 23684
rect 18417 23681 18429 23684
rect 18463 23681 18475 23715
rect 18417 23675 18475 23681
rect 18509 23715 18567 23721
rect 18509 23681 18521 23715
rect 18555 23712 18567 23715
rect 18555 23684 18736 23712
rect 18555 23681 18567 23684
rect 18509 23675 18567 23681
rect 18598 23644 18604 23656
rect 18156 23616 18604 23644
rect 17451 23613 17463 23616
rect 17405 23607 17463 23613
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 18708 23644 18736 23684
rect 18782 23672 18788 23724
rect 18840 23672 18846 23724
rect 20070 23672 20076 23724
rect 20128 23712 20134 23724
rect 20640 23721 20668 23752
rect 22554 23740 22560 23792
rect 22612 23780 22618 23792
rect 24596 23789 24624 23820
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 26973 23851 27031 23857
rect 26973 23817 26985 23851
rect 27019 23848 27031 23851
rect 27154 23848 27160 23860
rect 27019 23820 27160 23848
rect 27019 23817 27031 23820
rect 26973 23811 27031 23817
rect 27154 23808 27160 23820
rect 27212 23808 27218 23860
rect 27525 23851 27583 23857
rect 27525 23817 27537 23851
rect 27571 23817 27583 23851
rect 27525 23811 27583 23817
rect 30285 23851 30343 23857
rect 30285 23817 30297 23851
rect 30331 23848 30343 23851
rect 30742 23848 30748 23860
rect 30331 23820 30748 23848
rect 30331 23817 30343 23820
rect 30285 23811 30343 23817
rect 24581 23783 24639 23789
rect 22612 23752 23060 23780
rect 22612 23740 22618 23752
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 20128 23684 20269 23712
rect 20128 23672 20134 23684
rect 20257 23681 20269 23684
rect 20303 23712 20315 23715
rect 20533 23715 20591 23721
rect 20533 23712 20545 23715
rect 20303 23684 20545 23712
rect 20303 23681 20315 23684
rect 20257 23675 20315 23681
rect 20533 23681 20545 23684
rect 20579 23681 20591 23715
rect 20533 23675 20591 23681
rect 20625 23715 20683 23721
rect 20625 23681 20637 23715
rect 20671 23681 20683 23715
rect 20625 23675 20683 23681
rect 22097 23715 22155 23721
rect 22097 23681 22109 23715
rect 22143 23712 22155 23715
rect 22738 23712 22744 23724
rect 22143 23684 22744 23712
rect 22143 23681 22155 23684
rect 22097 23675 22155 23681
rect 22738 23672 22744 23684
rect 22796 23672 22802 23724
rect 23032 23721 23060 23752
rect 24581 23749 24593 23783
rect 24627 23749 24639 23783
rect 26142 23780 26148 23792
rect 25806 23752 26148 23780
rect 24581 23743 24639 23749
rect 26142 23740 26148 23752
rect 26200 23740 26206 23792
rect 26234 23740 26240 23792
rect 26292 23780 26298 23792
rect 27338 23780 27344 23792
rect 26292 23752 27344 23780
rect 26292 23740 26298 23752
rect 27338 23740 27344 23752
rect 27396 23740 27402 23792
rect 27430 23740 27436 23792
rect 27488 23780 27494 23792
rect 27540 23780 27568 23811
rect 30742 23808 30748 23820
rect 30800 23808 30806 23860
rect 31662 23848 31668 23860
rect 31128 23820 31668 23848
rect 27488 23752 27568 23780
rect 27893 23783 27951 23789
rect 27488 23740 27494 23752
rect 27893 23749 27905 23783
rect 27939 23780 27951 23783
rect 27982 23780 27988 23792
rect 27939 23752 27988 23780
rect 27939 23749 27951 23752
rect 27893 23743 27951 23749
rect 27982 23740 27988 23752
rect 28040 23780 28046 23792
rect 28353 23783 28411 23789
rect 28353 23780 28365 23783
rect 28040 23752 28365 23780
rect 28040 23740 28046 23752
rect 28353 23749 28365 23752
rect 28399 23749 28411 23783
rect 28353 23743 28411 23749
rect 23017 23715 23075 23721
rect 23017 23681 23029 23715
rect 23063 23712 23075 23715
rect 24210 23712 24216 23724
rect 23063 23684 24216 23712
rect 23063 23681 23075 23684
rect 23017 23675 23075 23681
rect 24210 23672 24216 23684
rect 24268 23672 24274 23724
rect 24302 23672 24308 23724
rect 24360 23672 24366 23724
rect 26050 23672 26056 23724
rect 26108 23672 26114 23724
rect 27157 23715 27215 23721
rect 27157 23681 27169 23715
rect 27203 23712 27215 23715
rect 27798 23712 27804 23724
rect 27203 23684 27804 23712
rect 27203 23681 27215 23684
rect 27157 23675 27215 23681
rect 27798 23672 27804 23684
rect 27856 23672 27862 23724
rect 28718 23712 28724 23724
rect 28000 23684 28724 23712
rect 19242 23644 19248 23656
rect 18708 23616 19248 23644
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 20165 23647 20223 23653
rect 20165 23644 20177 23647
rect 19392 23616 20177 23644
rect 19392 23604 19398 23616
rect 20165 23613 20177 23616
rect 20211 23644 20223 23647
rect 20349 23647 20407 23653
rect 20349 23644 20361 23647
rect 20211 23616 20361 23644
rect 20211 23613 20223 23616
rect 20165 23607 20223 23613
rect 20349 23613 20361 23616
rect 20395 23613 20407 23647
rect 23293 23647 23351 23653
rect 23293 23644 23305 23647
rect 20349 23607 20407 23613
rect 22066 23616 23305 23644
rect 17497 23579 17555 23585
rect 17497 23576 17509 23579
rect 16224 23548 17509 23576
rect 13449 23539 13507 23545
rect 17497 23545 17509 23548
rect 17543 23545 17555 23579
rect 17497 23539 17555 23545
rect 18046 23536 18052 23588
rect 18104 23576 18110 23588
rect 18104 23548 18644 23576
rect 18104 23536 18110 23548
rect 18616 23520 18644 23548
rect 19886 23536 19892 23588
rect 19944 23576 19950 23588
rect 22066 23576 22094 23616
rect 23293 23613 23305 23616
rect 23339 23644 23351 23647
rect 25038 23644 25044 23656
rect 23339 23616 25044 23644
rect 23339 23613 23351 23616
rect 23293 23607 23351 23613
rect 25038 23604 25044 23616
rect 25096 23604 25102 23656
rect 26068 23644 26096 23672
rect 26786 23644 26792 23656
rect 26068 23616 26792 23644
rect 26786 23604 26792 23616
rect 26844 23644 26850 23656
rect 27433 23647 27491 23653
rect 27433 23644 27445 23647
rect 26844 23616 27445 23644
rect 26844 23604 26850 23616
rect 27433 23613 27445 23616
rect 27479 23644 27491 23647
rect 27479 23636 27844 23644
rect 27890 23636 27896 23656
rect 27479 23616 27896 23636
rect 27479 23613 27491 23616
rect 27433 23607 27491 23613
rect 27816 23608 27896 23616
rect 27890 23604 27896 23608
rect 27948 23604 27954 23656
rect 28000 23653 28028 23684
rect 28718 23672 28724 23684
rect 28776 23672 28782 23724
rect 30193 23715 30251 23721
rect 30193 23681 30205 23715
rect 30239 23712 30251 23715
rect 30650 23712 30656 23724
rect 30239 23684 30656 23712
rect 30239 23681 30251 23684
rect 30193 23675 30251 23681
rect 30650 23672 30656 23684
rect 30708 23672 30714 23724
rect 31018 23712 31024 23724
rect 30852 23684 31024 23712
rect 27985 23647 28043 23653
rect 27985 23613 27997 23647
rect 28031 23613 28043 23647
rect 27985 23607 28043 23613
rect 28074 23604 28080 23656
rect 28132 23604 28138 23656
rect 28350 23604 28356 23656
rect 28408 23644 28414 23656
rect 28905 23647 28963 23653
rect 28905 23644 28917 23647
rect 28408 23616 28917 23644
rect 28408 23604 28414 23616
rect 28905 23613 28917 23616
rect 28951 23613 28963 23647
rect 30852 23644 30880 23684
rect 31018 23672 31024 23684
rect 31076 23672 31082 23724
rect 31128 23721 31156 23820
rect 31662 23808 31668 23820
rect 31720 23808 31726 23860
rect 34974 23808 34980 23860
rect 35032 23857 35038 23860
rect 35032 23851 35051 23857
rect 35039 23848 35051 23851
rect 40402 23848 40408 23860
rect 35039 23820 35388 23848
rect 35039 23817 35051 23820
rect 35032 23811 35051 23817
rect 35032 23808 35038 23811
rect 31294 23740 31300 23792
rect 31352 23740 31358 23792
rect 34698 23740 34704 23792
rect 34756 23780 34762 23792
rect 34793 23783 34851 23789
rect 34793 23780 34805 23783
rect 34756 23752 34805 23780
rect 34756 23740 34762 23752
rect 34793 23749 34805 23752
rect 34839 23749 34851 23783
rect 35158 23780 35164 23792
rect 34793 23743 34851 23749
rect 34900 23752 35164 23780
rect 31113 23715 31171 23721
rect 31113 23681 31125 23715
rect 31159 23681 31171 23715
rect 31665 23715 31723 23721
rect 31665 23712 31677 23715
rect 31113 23675 31171 23681
rect 31312 23684 31677 23712
rect 28905 23607 28963 23613
rect 29656 23616 30880 23644
rect 30929 23647 30987 23653
rect 19944 23548 22094 23576
rect 19944 23536 19950 23548
rect 25682 23536 25688 23588
rect 25740 23576 25746 23588
rect 25866 23576 25872 23588
rect 25740 23548 25872 23576
rect 25740 23536 25746 23548
rect 25866 23536 25872 23548
rect 25924 23576 25930 23588
rect 26053 23579 26111 23585
rect 26053 23576 26065 23579
rect 25924 23548 26065 23576
rect 25924 23536 25930 23548
rect 26053 23545 26065 23548
rect 26099 23545 26111 23579
rect 26053 23539 26111 23545
rect 27246 23536 27252 23588
rect 27304 23576 27310 23588
rect 27341 23579 27399 23585
rect 27341 23576 27353 23579
rect 27304 23548 27353 23576
rect 27304 23536 27310 23548
rect 27341 23545 27353 23548
rect 27387 23545 27399 23579
rect 27341 23539 27399 23545
rect 11379 23480 12940 23508
rect 11379 23477 11391 23480
rect 11333 23471 11391 23477
rect 12986 23468 12992 23520
rect 13044 23508 13050 23520
rect 13814 23508 13820 23520
rect 13044 23480 13820 23508
rect 13044 23468 13050 23480
rect 13814 23468 13820 23480
rect 13872 23508 13878 23520
rect 15654 23508 15660 23520
rect 13872 23480 15660 23508
rect 13872 23468 13878 23480
rect 15654 23468 15660 23480
rect 15712 23468 15718 23520
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 16025 23511 16083 23517
rect 16025 23508 16037 23511
rect 15988 23480 16037 23508
rect 15988 23468 15994 23480
rect 16025 23477 16037 23480
rect 16071 23477 16083 23511
rect 16025 23471 16083 23477
rect 17954 23468 17960 23520
rect 18012 23508 18018 23520
rect 18233 23511 18291 23517
rect 18233 23508 18245 23511
rect 18012 23480 18245 23508
rect 18012 23468 18018 23480
rect 18233 23477 18245 23480
rect 18279 23477 18291 23511
rect 18233 23471 18291 23477
rect 18598 23468 18604 23520
rect 18656 23468 18662 23520
rect 20162 23468 20168 23520
rect 20220 23468 20226 23520
rect 24302 23468 24308 23520
rect 24360 23508 24366 23520
rect 25130 23508 25136 23520
rect 24360 23480 25136 23508
rect 24360 23468 24366 23480
rect 25130 23468 25136 23480
rect 25188 23468 25194 23520
rect 25774 23468 25780 23520
rect 25832 23508 25838 23520
rect 29656 23508 29684 23616
rect 30929 23613 30941 23647
rect 30975 23644 30987 23647
rect 31312 23644 31340 23684
rect 31665 23681 31677 23684
rect 31711 23712 31723 23715
rect 31754 23712 31760 23724
rect 31711 23684 31760 23712
rect 31711 23681 31723 23684
rect 31665 23675 31723 23681
rect 31754 23672 31760 23684
rect 31812 23712 31818 23724
rect 32306 23712 32312 23724
rect 31812 23684 32312 23712
rect 31812 23672 31818 23684
rect 32306 23672 32312 23684
rect 32364 23672 32370 23724
rect 34606 23672 34612 23724
rect 34664 23712 34670 23724
rect 34900 23712 34928 23752
rect 35158 23740 35164 23752
rect 35216 23740 35222 23792
rect 35360 23780 35388 23820
rect 37292 23820 40408 23848
rect 35360 23752 35480 23780
rect 35452 23724 35480 23752
rect 34664 23684 34928 23712
rect 34664 23672 34670 23684
rect 34974 23672 34980 23724
rect 35032 23712 35038 23724
rect 35345 23715 35403 23721
rect 35345 23712 35357 23715
rect 35032 23684 35357 23712
rect 35032 23672 35038 23684
rect 35345 23681 35357 23684
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 35434 23672 35440 23724
rect 35492 23672 35498 23724
rect 36998 23672 37004 23724
rect 37056 23712 37062 23724
rect 37292 23721 37320 23820
rect 37550 23740 37556 23792
rect 37608 23740 37614 23792
rect 39500 23721 39528 23820
rect 40402 23808 40408 23820
rect 40460 23808 40466 23860
rect 39758 23740 39764 23792
rect 39816 23740 39822 23792
rect 41046 23780 41052 23792
rect 40986 23752 41052 23780
rect 41046 23740 41052 23752
rect 41104 23740 41110 23792
rect 41690 23740 41696 23792
rect 41748 23740 41754 23792
rect 37277 23715 37335 23721
rect 37277 23712 37289 23715
rect 37056 23684 37289 23712
rect 37056 23672 37062 23684
rect 37277 23681 37289 23684
rect 37323 23681 37335 23715
rect 39485 23715 39543 23721
rect 38686 23684 38792 23712
rect 37277 23675 37335 23681
rect 38764 23656 38792 23684
rect 39485 23681 39497 23715
rect 39531 23681 39543 23715
rect 39485 23675 39543 23681
rect 41138 23672 41144 23724
rect 41196 23712 41202 23724
rect 41196 23684 41276 23712
rect 41196 23672 41202 23684
rect 30975 23616 31340 23644
rect 31389 23647 31447 23653
rect 30975 23613 30987 23616
rect 30929 23607 30987 23613
rect 31389 23613 31401 23647
rect 31435 23644 31447 23647
rect 32766 23644 32772 23656
rect 31435 23616 32772 23644
rect 31435 23613 31447 23616
rect 31389 23607 31447 23613
rect 29730 23536 29736 23588
rect 29788 23576 29794 23588
rect 31404 23576 31432 23607
rect 32766 23604 32772 23616
rect 32824 23644 32830 23656
rect 34514 23644 34520 23656
rect 32824 23616 34520 23644
rect 32824 23604 32830 23616
rect 34514 23604 34520 23616
rect 34572 23644 34578 23656
rect 35621 23647 35679 23653
rect 35621 23644 35633 23647
rect 34572 23616 35633 23644
rect 34572 23604 34578 23616
rect 35621 23613 35633 23616
rect 35667 23644 35679 23647
rect 36170 23644 36176 23656
rect 35667 23616 36176 23644
rect 35667 23613 35679 23616
rect 35621 23607 35679 23613
rect 36170 23604 36176 23616
rect 36228 23604 36234 23656
rect 38746 23604 38752 23656
rect 38804 23604 38810 23656
rect 39022 23604 39028 23656
rect 39080 23604 39086 23656
rect 41248 23653 41276 23684
rect 41414 23672 41420 23724
rect 41472 23712 41478 23724
rect 41509 23715 41567 23721
rect 41509 23712 41521 23715
rect 41472 23684 41521 23712
rect 41472 23672 41478 23684
rect 41509 23681 41521 23684
rect 41555 23681 41567 23715
rect 41509 23675 41567 23681
rect 41598 23672 41604 23724
rect 41656 23672 41662 23724
rect 41877 23715 41935 23721
rect 41877 23681 41889 23715
rect 41923 23712 41935 23715
rect 42058 23712 42064 23724
rect 41923 23684 42064 23712
rect 41923 23681 41935 23684
rect 41877 23675 41935 23681
rect 42058 23672 42064 23684
rect 42116 23672 42122 23724
rect 41233 23647 41291 23653
rect 41233 23613 41245 23647
rect 41279 23613 41291 23647
rect 41233 23607 41291 23613
rect 29788 23548 31432 23576
rect 31573 23579 31631 23585
rect 29788 23536 29794 23548
rect 31573 23545 31585 23579
rect 31619 23576 31631 23579
rect 31662 23576 31668 23588
rect 31619 23548 31668 23576
rect 31619 23545 31631 23548
rect 31573 23539 31631 23545
rect 31662 23536 31668 23548
rect 31720 23576 31726 23588
rect 35161 23579 35219 23585
rect 35161 23576 35173 23579
rect 31720 23548 35173 23576
rect 31720 23536 31726 23548
rect 35161 23545 35173 23548
rect 35207 23576 35219 23579
rect 35710 23576 35716 23588
rect 35207 23548 35716 23576
rect 35207 23545 35219 23548
rect 35161 23539 35219 23545
rect 35710 23536 35716 23548
rect 35768 23536 35774 23588
rect 25832 23480 29684 23508
rect 25832 23468 25838 23480
rect 31478 23468 31484 23520
rect 31536 23468 31542 23520
rect 34790 23468 34796 23520
rect 34848 23508 34854 23520
rect 34974 23508 34980 23520
rect 34848 23480 34980 23508
rect 34848 23468 34854 23480
rect 34974 23468 34980 23480
rect 35032 23468 35038 23520
rect 35529 23511 35587 23517
rect 35529 23477 35541 23511
rect 35575 23508 35587 23511
rect 36538 23508 36544 23520
rect 35575 23480 36544 23508
rect 35575 23477 35587 23480
rect 35529 23471 35587 23477
rect 36538 23468 36544 23480
rect 36596 23468 36602 23520
rect 41322 23468 41328 23520
rect 41380 23468 41386 23520
rect 1104 23418 42504 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 42504 23418
rect 1104 23344 42504 23366
rect 1394 23264 1400 23316
rect 1452 23264 1458 23316
rect 5442 23264 5448 23316
rect 5500 23264 5506 23316
rect 5626 23264 5632 23316
rect 5684 23264 5690 23316
rect 6288 23276 20668 23304
rect 106 23128 112 23180
rect 164 23168 170 23180
rect 6288 23168 6316 23276
rect 7374 23196 7380 23248
rect 7432 23196 7438 23248
rect 11517 23239 11575 23245
rect 11517 23205 11529 23239
rect 11563 23236 11575 23239
rect 12434 23236 12440 23248
rect 11563 23208 12440 23236
rect 11563 23205 11575 23208
rect 11517 23199 11575 23205
rect 12434 23196 12440 23208
rect 12492 23196 12498 23248
rect 14369 23239 14427 23245
rect 14369 23236 14381 23239
rect 13648 23208 14381 23236
rect 164 23140 6316 23168
rect 164 23128 170 23140
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 13648 23168 13676 23208
rect 14369 23205 14381 23208
rect 14415 23236 14427 23239
rect 14829 23239 14887 23245
rect 14829 23236 14841 23239
rect 14415 23208 14841 23236
rect 14415 23205 14427 23208
rect 14369 23199 14427 23205
rect 14829 23205 14841 23208
rect 14875 23236 14887 23239
rect 15470 23236 15476 23248
rect 14875 23208 15476 23236
rect 14875 23205 14887 23208
rect 14829 23199 14887 23205
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 17405 23239 17463 23245
rect 17405 23236 17417 23239
rect 17092 23208 17417 23236
rect 17092 23196 17098 23208
rect 17405 23205 17417 23208
rect 17451 23205 17463 23239
rect 17405 23199 17463 23205
rect 12216 23140 13676 23168
rect 13725 23171 13783 23177
rect 12216 23128 12222 23140
rect 13725 23137 13737 23171
rect 13771 23168 13783 23171
rect 13906 23168 13912 23180
rect 13771 23140 13912 23168
rect 13771 23137 13783 23140
rect 13725 23131 13783 23137
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 14182 23128 14188 23180
rect 14240 23128 14246 23180
rect 14550 23128 14556 23180
rect 14608 23168 14614 23180
rect 15197 23171 15255 23177
rect 15197 23168 15209 23171
rect 14608 23140 15209 23168
rect 14608 23128 14614 23140
rect 3145 23103 3203 23109
rect 3145 23069 3157 23103
rect 3191 23100 3203 23103
rect 3234 23100 3240 23112
rect 3191 23072 3240 23100
rect 3191 23069 3203 23072
rect 3145 23063 3203 23069
rect 3234 23060 3240 23072
rect 3292 23060 3298 23112
rect 7098 23060 7104 23112
rect 7156 23060 7162 23112
rect 7190 23060 7196 23112
rect 7248 23100 7254 23112
rect 7285 23103 7343 23109
rect 7285 23100 7297 23103
rect 7248 23072 7297 23100
rect 7248 23060 7254 23072
rect 7285 23069 7297 23072
rect 7331 23100 7343 23103
rect 7374 23100 7380 23112
rect 7331 23072 7380 23100
rect 7331 23069 7343 23072
rect 7285 23063 7343 23069
rect 7374 23060 7380 23072
rect 7432 23060 7438 23112
rect 7466 23060 7472 23112
rect 7524 23060 7530 23112
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23100 7619 23103
rect 7650 23100 7656 23112
rect 7607 23072 7656 23100
rect 7607 23069 7619 23072
rect 7561 23063 7619 23069
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 10134 23060 10140 23112
rect 10192 23060 10198 23112
rect 10226 23060 10232 23112
rect 10284 23100 10290 23112
rect 10393 23103 10451 23109
rect 10393 23100 10405 23103
rect 10284 23072 10405 23100
rect 10284 23060 10290 23072
rect 10393 23069 10405 23072
rect 10439 23069 10451 23103
rect 10393 23063 10451 23069
rect 12986 23060 12992 23112
rect 13044 23100 13050 23112
rect 13170 23100 13176 23112
rect 13044 23072 13176 23100
rect 13044 23060 13050 23072
rect 13170 23060 13176 23072
rect 13228 23100 13234 23112
rect 13449 23103 13507 23109
rect 13449 23100 13461 23103
rect 13228 23072 13461 23100
rect 13228 23060 13234 23072
rect 13449 23069 13461 23072
rect 13495 23069 13507 23103
rect 13449 23063 13507 23069
rect 13630 23060 13636 23112
rect 13688 23060 13694 23112
rect 13817 23103 13875 23109
rect 13817 23069 13829 23103
rect 13863 23069 13875 23103
rect 13817 23063 13875 23069
rect 2406 22992 2412 23044
rect 2464 22992 2470 23044
rect 2866 22992 2872 23044
rect 2924 22992 2930 23044
rect 5261 23035 5319 23041
rect 5261 23001 5273 23035
rect 5307 23032 5319 23035
rect 5350 23032 5356 23044
rect 5307 23004 5356 23032
rect 5307 23001 5319 23004
rect 5261 22995 5319 23001
rect 5350 22992 5356 23004
rect 5408 22992 5414 23044
rect 13722 22992 13728 23044
rect 13780 23032 13786 23044
rect 13832 23032 13860 23063
rect 14458 23060 14464 23112
rect 14516 23060 14522 23112
rect 14660 23109 14688 23140
rect 15197 23137 15209 23140
rect 15243 23137 15255 23171
rect 15197 23131 15255 23137
rect 16666 23128 16672 23180
rect 16724 23168 16730 23180
rect 16724 23140 17724 23168
rect 16724 23128 16730 23140
rect 14645 23103 14703 23109
rect 14645 23069 14657 23103
rect 14691 23069 14703 23103
rect 14645 23063 14703 23069
rect 14660 23032 14688 23063
rect 14826 23060 14832 23112
rect 14884 23060 14890 23112
rect 15102 23060 15108 23112
rect 15160 23060 15166 23112
rect 15286 23060 15292 23112
rect 15344 23060 15350 23112
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 13780 23004 14688 23032
rect 13780 22992 13786 23004
rect 5471 22967 5529 22973
rect 5471 22933 5483 22967
rect 5517 22964 5529 22967
rect 5994 22964 6000 22976
rect 5517 22936 6000 22964
rect 5517 22933 5529 22936
rect 5471 22927 5529 22933
rect 5994 22924 6000 22936
rect 6052 22924 6058 22976
rect 7742 22924 7748 22976
rect 7800 22924 7806 22976
rect 12618 22924 12624 22976
rect 12676 22964 12682 22976
rect 12897 22967 12955 22973
rect 12897 22964 12909 22967
rect 12676 22936 12909 22964
rect 12676 22924 12682 22936
rect 12897 22933 12909 22936
rect 12943 22933 12955 22967
rect 12897 22927 12955 22933
rect 14182 22924 14188 22976
rect 14240 22924 14246 22976
rect 14844 22964 14872 23060
rect 15396 22964 15424 23063
rect 15562 23060 15568 23112
rect 15620 23100 15626 23112
rect 17696 23109 17724 23140
rect 19518 23128 19524 23180
rect 19576 23168 19582 23180
rect 19705 23171 19763 23177
rect 19705 23168 19717 23171
rect 19576 23140 19717 23168
rect 19576 23128 19582 23140
rect 19705 23137 19717 23140
rect 19751 23137 19763 23171
rect 19705 23131 19763 23137
rect 19886 23128 19892 23180
rect 19944 23128 19950 23180
rect 15657 23103 15715 23109
rect 15657 23100 15669 23103
rect 15620 23072 15669 23100
rect 15620 23060 15626 23072
rect 15657 23069 15669 23072
rect 15703 23069 15715 23103
rect 15657 23063 15715 23069
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23069 17739 23103
rect 17681 23063 17739 23069
rect 18138 23060 18144 23112
rect 18196 23100 18202 23112
rect 19904 23100 19932 23128
rect 20640 23109 20668 23276
rect 21726 23264 21732 23316
rect 21784 23304 21790 23316
rect 21910 23304 21916 23316
rect 21784 23276 21916 23304
rect 21784 23264 21790 23276
rect 21910 23264 21916 23276
rect 21968 23264 21974 23316
rect 28718 23264 28724 23316
rect 28776 23304 28782 23316
rect 39117 23307 39175 23313
rect 28776 23276 38792 23304
rect 28776 23264 28782 23276
rect 28994 23196 29000 23248
rect 29052 23236 29058 23248
rect 34698 23236 34704 23248
rect 29052 23208 31800 23236
rect 29052 23196 29058 23208
rect 30558 23128 30564 23180
rect 30616 23168 30622 23180
rect 30929 23171 30987 23177
rect 30929 23168 30941 23171
rect 30616 23140 30941 23168
rect 30616 23128 30622 23140
rect 30929 23137 30941 23140
rect 30975 23137 30987 23171
rect 30929 23131 30987 23137
rect 31294 23128 31300 23180
rect 31352 23168 31358 23180
rect 31772 23177 31800 23208
rect 34256 23208 34704 23236
rect 31389 23171 31447 23177
rect 31389 23168 31401 23171
rect 31352 23140 31401 23168
rect 31352 23128 31358 23140
rect 31389 23137 31401 23140
rect 31435 23137 31447 23171
rect 31389 23131 31447 23137
rect 31757 23171 31815 23177
rect 31757 23137 31769 23171
rect 31803 23137 31815 23171
rect 31757 23131 31815 23137
rect 31849 23171 31907 23177
rect 31849 23137 31861 23171
rect 31895 23168 31907 23171
rect 32030 23168 32036 23180
rect 31895 23140 32036 23168
rect 31895 23137 31907 23140
rect 31849 23131 31907 23137
rect 32030 23128 32036 23140
rect 32088 23168 32094 23180
rect 32214 23168 32220 23180
rect 32088 23140 32220 23168
rect 32088 23128 32094 23140
rect 32214 23128 32220 23140
rect 32272 23128 32278 23180
rect 34256 23168 34284 23208
rect 34698 23196 34704 23208
rect 34756 23196 34762 23248
rect 35268 23208 35847 23236
rect 33428 23140 34284 23168
rect 33428 23112 33456 23140
rect 18196 23072 19932 23100
rect 20625 23103 20683 23109
rect 18196 23060 18202 23072
rect 20625 23069 20637 23103
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 22649 23103 22707 23109
rect 22649 23069 22661 23103
rect 22695 23100 22707 23103
rect 22830 23100 22836 23112
rect 22695 23072 22836 23100
rect 22695 23069 22707 23072
rect 22649 23063 22707 23069
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 24670 23060 24676 23112
rect 24728 23100 24734 23112
rect 25498 23100 25504 23112
rect 24728 23072 25504 23100
rect 24728 23060 24734 23072
rect 25498 23060 25504 23072
rect 25556 23060 25562 23112
rect 25590 23060 25596 23112
rect 25648 23060 25654 23112
rect 25866 23060 25872 23112
rect 25924 23060 25930 23112
rect 25958 23060 25964 23112
rect 26016 23060 26022 23112
rect 27706 23060 27712 23112
rect 27764 23100 27770 23112
rect 28902 23100 28908 23112
rect 27764 23072 28908 23100
rect 27764 23060 27770 23072
rect 28902 23060 28908 23072
rect 28960 23100 28966 23112
rect 28997 23103 29055 23109
rect 28997 23100 29009 23103
rect 28960 23072 29009 23100
rect 28960 23060 28966 23072
rect 28997 23069 29009 23072
rect 29043 23069 29055 23103
rect 28997 23063 29055 23069
rect 31478 23060 31484 23112
rect 31536 23060 31542 23112
rect 33410 23060 33416 23112
rect 33468 23060 33474 23112
rect 33502 23060 33508 23112
rect 33560 23060 33566 23112
rect 34256 23109 34284 23140
rect 34514 23128 34520 23180
rect 34572 23128 34578 23180
rect 35268 23112 35296 23208
rect 35345 23171 35403 23177
rect 35345 23137 35357 23171
rect 35391 23168 35403 23171
rect 35526 23168 35532 23180
rect 35391 23140 35532 23168
rect 35391 23137 35403 23140
rect 35345 23131 35403 23137
rect 35526 23128 35532 23140
rect 35584 23128 35590 23180
rect 35710 23128 35716 23180
rect 35768 23128 35774 23180
rect 35819 23168 35847 23208
rect 35819 23140 35940 23168
rect 34241 23103 34299 23109
rect 34241 23069 34253 23103
rect 34287 23069 34299 23103
rect 34241 23063 34299 23069
rect 34333 23103 34391 23109
rect 34333 23069 34345 23103
rect 34379 23100 34391 23103
rect 35250 23100 35256 23112
rect 34379 23072 35256 23100
rect 34379 23069 34391 23072
rect 34333 23063 34391 23069
rect 35250 23060 35256 23072
rect 35308 23060 35314 23112
rect 35805 23103 35863 23109
rect 35805 23069 35817 23103
rect 35851 23069 35863 23103
rect 35912 23100 35940 23140
rect 35986 23128 35992 23180
rect 36044 23168 36050 23180
rect 36081 23171 36139 23177
rect 36081 23168 36093 23171
rect 36044 23140 36093 23168
rect 36044 23128 36050 23140
rect 36081 23137 36093 23140
rect 36127 23168 36139 23171
rect 36817 23171 36875 23177
rect 36817 23168 36829 23171
rect 36127 23140 36829 23168
rect 36127 23137 36139 23140
rect 36081 23131 36139 23137
rect 36817 23137 36829 23140
rect 36863 23137 36875 23171
rect 36817 23131 36875 23137
rect 36449 23103 36507 23109
rect 36449 23100 36461 23103
rect 35912 23072 36461 23100
rect 35805 23063 35863 23069
rect 36449 23069 36461 23072
rect 36495 23069 36507 23103
rect 36449 23063 36507 23069
rect 15930 22992 15936 23044
rect 15988 22992 15994 23044
rect 18046 23032 18052 23044
rect 17158 23004 18052 23032
rect 18046 22992 18052 23004
rect 18104 22992 18110 23044
rect 19610 22992 19616 23044
rect 19668 22992 19674 23044
rect 25222 22992 25228 23044
rect 25280 23032 25286 23044
rect 25777 23035 25835 23041
rect 25777 23032 25789 23035
rect 25280 23004 25789 23032
rect 25280 22992 25286 23004
rect 25777 23001 25789 23004
rect 25823 23001 25835 23035
rect 25777 22995 25835 23001
rect 28752 23035 28810 23041
rect 28752 23001 28764 23035
rect 28798 23032 28810 23035
rect 29086 23032 29092 23044
rect 28798 23004 29092 23032
rect 28798 23001 28810 23004
rect 28752 22995 28810 23001
rect 29086 22992 29092 23004
rect 29144 22992 29150 23044
rect 30745 23035 30803 23041
rect 30745 23001 30757 23035
rect 30791 23032 30803 23035
rect 31754 23032 31760 23044
rect 30791 23004 31760 23032
rect 30791 23001 30803 23004
rect 30745 22995 30803 23001
rect 31754 22992 31760 23004
rect 31812 22992 31818 23044
rect 33260 23035 33318 23041
rect 33260 23001 33272 23035
rect 33306 23032 33318 23035
rect 34517 23035 34575 23041
rect 33306 23004 34468 23032
rect 33306 23001 33318 23004
rect 33260 22995 33318 23001
rect 14844 22936 15424 22964
rect 15565 22967 15623 22973
rect 15565 22933 15577 22967
rect 15611 22964 15623 22967
rect 16574 22964 16580 22976
rect 15611 22936 16580 22964
rect 15611 22933 15623 22936
rect 15565 22927 15623 22933
rect 16574 22924 16580 22936
rect 16632 22924 16638 22976
rect 18782 22924 18788 22976
rect 18840 22964 18846 22976
rect 19245 22967 19303 22973
rect 19245 22964 19257 22967
rect 18840 22936 19257 22964
rect 18840 22924 18846 22936
rect 19245 22933 19257 22936
rect 19291 22933 19303 22967
rect 19245 22927 19303 22933
rect 22462 22924 22468 22976
rect 22520 22964 22526 22976
rect 23201 22967 23259 22973
rect 23201 22964 23213 22967
rect 22520 22936 23213 22964
rect 22520 22924 22526 22936
rect 23201 22933 23213 22936
rect 23247 22964 23259 22967
rect 23382 22964 23388 22976
rect 23247 22936 23388 22964
rect 23247 22933 23259 22936
rect 23201 22927 23259 22933
rect 23382 22924 23388 22936
rect 23440 22924 23446 22976
rect 26145 22967 26203 22973
rect 26145 22933 26157 22967
rect 26191 22964 26203 22967
rect 26418 22964 26424 22976
rect 26191 22936 26424 22964
rect 26191 22933 26203 22936
rect 26145 22927 26203 22933
rect 26418 22924 26424 22936
rect 26476 22924 26482 22976
rect 27154 22924 27160 22976
rect 27212 22964 27218 22976
rect 27617 22967 27675 22973
rect 27617 22964 27629 22967
rect 27212 22936 27629 22964
rect 27212 22924 27218 22936
rect 27617 22933 27629 22936
rect 27663 22933 27675 22967
rect 27617 22927 27675 22933
rect 30282 22924 30288 22976
rect 30340 22964 30346 22976
rect 30377 22967 30435 22973
rect 30377 22964 30389 22967
rect 30340 22936 30389 22964
rect 30340 22924 30346 22936
rect 30377 22933 30389 22936
rect 30423 22933 30435 22967
rect 30377 22927 30435 22933
rect 30837 22967 30895 22973
rect 30837 22933 30849 22967
rect 30883 22964 30895 22967
rect 31205 22967 31263 22973
rect 31205 22964 31217 22967
rect 30883 22936 31217 22964
rect 30883 22933 30895 22936
rect 30837 22927 30895 22933
rect 31205 22933 31217 22936
rect 31251 22933 31263 22967
rect 31205 22927 31263 22933
rect 32122 22924 32128 22976
rect 32180 22924 32186 22976
rect 34440 22964 34468 23004
rect 34517 23001 34529 23035
rect 34563 23032 34575 23035
rect 35820 23032 35848 23063
rect 36538 23059 36544 23111
rect 36596 23100 36602 23111
rect 36596 23072 36640 23100
rect 36596 23059 36602 23072
rect 38654 23060 38660 23112
rect 38712 23060 38718 23112
rect 38764 23100 38792 23276
rect 39117 23273 39129 23307
rect 39163 23304 39175 23307
rect 39298 23304 39304 23316
rect 39163 23276 39304 23304
rect 39163 23273 39175 23276
rect 39117 23267 39175 23273
rect 39298 23264 39304 23276
rect 39356 23264 39362 23316
rect 41690 23304 41696 23316
rect 39500 23276 41696 23304
rect 39301 23103 39359 23109
rect 39301 23100 39313 23103
rect 38764 23072 39313 23100
rect 39301 23069 39313 23072
rect 39347 23069 39359 23103
rect 39301 23063 39359 23069
rect 39390 23060 39396 23112
rect 39448 23060 39454 23112
rect 39500 23109 39528 23276
rect 41690 23264 41696 23276
rect 41748 23264 41754 23316
rect 39945 23171 40003 23177
rect 39945 23137 39957 23171
rect 39991 23168 40003 23171
rect 40681 23171 40739 23177
rect 40681 23168 40693 23171
rect 39991 23140 40693 23168
rect 39991 23137 40003 23140
rect 39945 23131 40003 23137
rect 40681 23137 40693 23140
rect 40727 23137 40739 23171
rect 40681 23131 40739 23137
rect 39485 23103 39543 23109
rect 39485 23069 39497 23103
rect 39531 23069 39543 23103
rect 39485 23063 39543 23069
rect 39669 23103 39727 23109
rect 39669 23069 39681 23103
rect 39715 23100 39727 23103
rect 40034 23100 40040 23112
rect 39715 23072 40040 23100
rect 39715 23069 39727 23072
rect 39669 23063 39727 23069
rect 40034 23060 40040 23072
rect 40092 23060 40098 23112
rect 40402 23060 40408 23112
rect 40460 23060 40466 23112
rect 34563 23004 35848 23032
rect 36173 23035 36231 23041
rect 34563 23001 34575 23004
rect 34517 22995 34575 23001
rect 36173 23001 36185 23035
rect 36219 23032 36231 23035
rect 36909 23035 36967 23041
rect 36219 23004 36492 23032
rect 36219 23001 36231 23004
rect 36173 22995 36231 23001
rect 34606 22964 34612 22976
rect 34440 22936 34612 22964
rect 34606 22924 34612 22936
rect 34664 22924 34670 22976
rect 34701 22967 34759 22973
rect 34701 22933 34713 22967
rect 34747 22964 34759 22967
rect 34882 22964 34888 22976
rect 34747 22936 34888 22964
rect 34747 22933 34759 22936
rect 34701 22927 34759 22933
rect 34882 22924 34888 22936
rect 34940 22924 34946 22976
rect 34974 22924 34980 22976
rect 35032 22964 35038 22976
rect 35069 22967 35127 22973
rect 35069 22964 35081 22967
rect 35032 22936 35081 22964
rect 35032 22924 35038 22936
rect 35069 22933 35081 22936
rect 35115 22933 35127 22967
rect 35069 22927 35127 22933
rect 35161 22967 35219 22973
rect 35161 22933 35173 22967
rect 35207 22964 35219 22967
rect 35529 22967 35587 22973
rect 35529 22964 35541 22967
rect 35207 22936 35541 22964
rect 35207 22933 35219 22936
rect 35161 22927 35219 22933
rect 35529 22933 35541 22936
rect 35575 22933 35587 22967
rect 35529 22927 35587 22933
rect 36262 22924 36268 22976
rect 36320 22924 36326 22976
rect 36464 22964 36492 23004
rect 36909 23001 36921 23035
rect 36955 23032 36967 23035
rect 36998 23032 37004 23044
rect 36955 23004 37004 23032
rect 36955 23001 36967 23004
rect 36909 22995 36967 23001
rect 36998 22992 37004 23004
rect 37056 22992 37062 23044
rect 37090 22992 37096 23044
rect 37148 23032 37154 23044
rect 40129 23035 40187 23041
rect 37148 23004 39344 23032
rect 37148 22992 37154 23004
rect 36814 22964 36820 22976
rect 36464 22936 36820 22964
rect 36814 22924 36820 22936
rect 36872 22924 36878 22976
rect 37734 22924 37740 22976
rect 37792 22964 37798 22976
rect 38013 22967 38071 22973
rect 38013 22964 38025 22967
rect 37792 22936 38025 22964
rect 37792 22924 37798 22936
rect 38013 22933 38025 22936
rect 38059 22933 38071 22967
rect 39316 22964 39344 23004
rect 40129 23001 40141 23035
rect 40175 23001 40187 23035
rect 40129 22995 40187 23001
rect 40313 23035 40371 23041
rect 40313 23001 40325 23035
rect 40359 23001 40371 23035
rect 40313 22995 40371 23001
rect 40144 22964 40172 22995
rect 39316 22936 40172 22964
rect 40328 22964 40356 22995
rect 41138 22992 41144 23044
rect 41196 22992 41202 23044
rect 41322 22964 41328 22976
rect 40328 22936 41328 22964
rect 38013 22927 38071 22933
rect 41322 22924 41328 22936
rect 41380 22924 41386 22976
rect 42058 22924 42064 22976
rect 42116 22964 42122 22976
rect 42153 22967 42211 22973
rect 42153 22964 42165 22967
rect 42116 22936 42165 22964
rect 42116 22924 42122 22936
rect 42153 22933 42165 22936
rect 42199 22933 42211 22967
rect 42153 22927 42211 22933
rect 1104 22874 42504 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 42504 22874
rect 1104 22800 42504 22822
rect 5718 22760 5724 22772
rect 2746 22732 4936 22760
rect 2406 22652 2412 22704
rect 2464 22692 2470 22704
rect 2746 22692 2774 22732
rect 4908 22692 4936 22732
rect 5552 22732 5724 22760
rect 5552 22704 5580 22732
rect 5718 22720 5724 22732
rect 5776 22720 5782 22772
rect 7098 22720 7104 22772
rect 7156 22760 7162 22772
rect 7926 22760 7932 22772
rect 7156 22732 7932 22760
rect 7156 22720 7162 22732
rect 7926 22720 7932 22732
rect 7984 22720 7990 22772
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 10597 22763 10655 22769
rect 10597 22760 10609 22763
rect 9916 22732 10609 22760
rect 9916 22720 9922 22732
rect 10597 22729 10609 22732
rect 10643 22729 10655 22763
rect 10597 22723 10655 22729
rect 12618 22720 12624 22772
rect 12676 22720 12682 22772
rect 13817 22763 13875 22769
rect 13817 22729 13829 22763
rect 13863 22760 13875 22763
rect 14458 22760 14464 22772
rect 13863 22732 14464 22760
rect 13863 22729 13875 22732
rect 13817 22723 13875 22729
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 15286 22720 15292 22772
rect 15344 22760 15350 22772
rect 16025 22763 16083 22769
rect 15344 22732 15884 22760
rect 15344 22720 15350 22732
rect 5534 22692 5540 22704
rect 2464 22664 2774 22692
rect 4830 22664 5540 22692
rect 2464 22652 2470 22664
rect 5534 22652 5540 22664
rect 5592 22652 5598 22704
rect 5626 22652 5632 22704
rect 5684 22692 5690 22704
rect 8018 22692 8024 22704
rect 5684 22664 8024 22692
rect 5684 22652 5690 22664
rect 8018 22652 8024 22664
rect 8076 22652 8082 22704
rect 10134 22692 10140 22704
rect 8128 22664 10140 22692
rect 7742 22584 7748 22636
rect 7800 22584 7806 22636
rect 8128 22633 8156 22664
rect 10134 22652 10140 22664
rect 10192 22652 10198 22704
rect 11146 22652 11152 22704
rect 11204 22692 11210 22704
rect 11701 22695 11759 22701
rect 11701 22692 11713 22695
rect 11204 22664 11713 22692
rect 11204 22652 11210 22664
rect 11701 22661 11713 22664
rect 11747 22692 11759 22695
rect 12066 22692 12072 22704
rect 11747 22664 12072 22692
rect 11747 22661 11759 22664
rect 11701 22655 11759 22661
rect 12066 22652 12072 22664
rect 12124 22692 12130 22704
rect 13722 22692 13728 22704
rect 12124 22664 13728 22692
rect 12124 22652 12130 22664
rect 13722 22652 13728 22664
rect 13780 22692 13786 22704
rect 13909 22695 13967 22701
rect 13909 22692 13921 22695
rect 13780 22664 13921 22692
rect 13780 22652 13786 22664
rect 13909 22661 13921 22664
rect 13955 22661 13967 22695
rect 13909 22655 13967 22661
rect 14182 22652 14188 22704
rect 14240 22692 14246 22704
rect 14553 22695 14611 22701
rect 14553 22692 14565 22695
rect 14240 22664 14565 22692
rect 14240 22652 14246 22664
rect 14553 22661 14565 22664
rect 14599 22661 14611 22695
rect 15856 22692 15884 22732
rect 16025 22729 16037 22763
rect 16071 22760 16083 22763
rect 16482 22760 16488 22772
rect 16071 22732 16488 22760
rect 16071 22729 16083 22732
rect 16025 22723 16083 22729
rect 16482 22720 16488 22732
rect 16540 22720 16546 22772
rect 18046 22760 18052 22772
rect 16592 22732 18052 22760
rect 16592 22692 16620 22732
rect 18046 22720 18052 22732
rect 18104 22760 18110 22772
rect 18104 22732 18920 22760
rect 18104 22720 18110 22732
rect 15778 22664 16620 22692
rect 14553 22655 14611 22661
rect 17586 22652 17592 22704
rect 17644 22652 17650 22704
rect 18782 22652 18788 22704
rect 18840 22652 18846 22704
rect 18892 22692 18920 22732
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 19794 22760 19800 22772
rect 19668 22732 19800 22760
rect 19668 22720 19674 22732
rect 19794 22720 19800 22732
rect 19852 22760 19858 22772
rect 20257 22763 20315 22769
rect 20257 22760 20269 22763
rect 19852 22732 20269 22760
rect 19852 22720 19858 22732
rect 20257 22729 20269 22732
rect 20303 22729 20315 22763
rect 22554 22760 22560 22772
rect 20257 22723 20315 22729
rect 21100 22732 22560 22760
rect 18892 22664 19274 22692
rect 20714 22652 20720 22704
rect 20772 22652 20778 22704
rect 8113 22627 8171 22633
rect 8113 22593 8125 22627
rect 8159 22593 8171 22627
rect 8369 22627 8427 22633
rect 8369 22624 8381 22627
rect 8113 22587 8171 22593
rect 8220 22596 8381 22624
rect 2774 22516 2780 22568
rect 2832 22556 2838 22568
rect 2869 22559 2927 22565
rect 2869 22556 2881 22559
rect 2832 22528 2881 22556
rect 2832 22516 2838 22528
rect 2869 22525 2881 22528
rect 2915 22525 2927 22559
rect 2869 22519 2927 22525
rect 3145 22559 3203 22565
rect 3145 22525 3157 22559
rect 3191 22556 3203 22559
rect 3234 22556 3240 22568
rect 3191 22528 3240 22556
rect 3191 22525 3203 22528
rect 3145 22519 3203 22525
rect 3234 22516 3240 22528
rect 3292 22556 3298 22568
rect 3421 22559 3479 22565
rect 3421 22556 3433 22559
rect 3292 22528 3433 22556
rect 3292 22516 3298 22528
rect 3421 22525 3433 22528
rect 3467 22525 3479 22559
rect 3421 22519 3479 22525
rect 3789 22559 3847 22565
rect 3789 22525 3801 22559
rect 3835 22556 3847 22559
rect 4706 22556 4712 22568
rect 3835 22528 4712 22556
rect 3835 22525 3847 22528
rect 3789 22519 3847 22525
rect 4706 22516 4712 22528
rect 4764 22516 4770 22568
rect 7650 22516 7656 22568
rect 7708 22516 7714 22568
rect 8220 22556 8248 22596
rect 8369 22593 8381 22596
rect 8415 22593 8427 22627
rect 8369 22587 8427 22593
rect 10229 22627 10287 22633
rect 10229 22593 10241 22627
rect 10275 22624 10287 22627
rect 11422 22624 11428 22636
rect 10275 22596 11428 22624
rect 10275 22593 10287 22596
rect 10229 22587 10287 22593
rect 7944 22528 8248 22556
rect 7561 22491 7619 22497
rect 7561 22457 7573 22491
rect 7607 22488 7619 22491
rect 7944 22488 7972 22528
rect 9585 22491 9643 22497
rect 9585 22488 9597 22491
rect 7607 22460 7972 22488
rect 9048 22460 9597 22488
rect 7607 22457 7619 22460
rect 7561 22451 7619 22457
rect 1394 22380 1400 22432
rect 1452 22380 1458 22432
rect 4798 22380 4804 22432
rect 4856 22420 4862 22432
rect 5169 22423 5227 22429
rect 5169 22420 5181 22423
rect 4856 22392 5181 22420
rect 4856 22380 4862 22392
rect 5169 22389 5181 22392
rect 5215 22420 5227 22423
rect 6822 22420 6828 22432
rect 5215 22392 6828 22420
rect 5215 22389 5227 22392
rect 5169 22383 5227 22389
rect 6822 22380 6828 22392
rect 6880 22380 6886 22432
rect 7742 22380 7748 22432
rect 7800 22420 7806 22432
rect 9048 22420 9076 22460
rect 9585 22457 9597 22460
rect 9631 22457 9643 22491
rect 9585 22451 9643 22457
rect 7800 22392 9076 22420
rect 9493 22423 9551 22429
rect 7800 22380 7806 22392
rect 9493 22389 9505 22423
rect 9539 22420 9551 22423
rect 10244 22420 10272 22587
rect 11422 22584 11428 22596
rect 11480 22584 11486 22636
rect 14274 22584 14280 22636
rect 14332 22584 14338 22636
rect 16206 22584 16212 22636
rect 16264 22584 16270 22636
rect 17954 22584 17960 22636
rect 18012 22584 18018 22636
rect 18138 22584 18144 22636
rect 18196 22584 18202 22636
rect 18230 22584 18236 22636
rect 18288 22584 18294 22636
rect 20622 22584 20628 22636
rect 20680 22584 20686 22636
rect 21100 22633 21128 22732
rect 22554 22720 22560 22732
rect 22612 22720 22618 22772
rect 24210 22720 24216 22772
rect 24268 22720 24274 22772
rect 24596 22732 25544 22760
rect 22462 22692 22468 22704
rect 21376 22664 22468 22692
rect 21376 22633 21404 22664
rect 22462 22652 22468 22664
rect 22520 22652 22526 22704
rect 24596 22692 24624 22732
rect 22756 22664 24624 22692
rect 20809 22627 20867 22633
rect 20809 22593 20821 22627
rect 20855 22593 20867 22627
rect 20809 22587 20867 22593
rect 20993 22627 21051 22633
rect 20993 22593 21005 22627
rect 21039 22593 21051 22627
rect 20993 22587 21051 22593
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 21361 22627 21419 22633
rect 21361 22593 21373 22627
rect 21407 22593 21419 22627
rect 21361 22587 21419 22593
rect 11241 22559 11299 22565
rect 11241 22525 11253 22559
rect 11287 22525 11299 22559
rect 11241 22519 11299 22525
rect 12161 22559 12219 22565
rect 12161 22525 12173 22559
rect 12207 22556 12219 22559
rect 12713 22559 12771 22565
rect 12713 22556 12725 22559
rect 12207 22528 12725 22556
rect 12207 22525 12219 22528
rect 12161 22519 12219 22525
rect 12713 22525 12725 22528
rect 12759 22525 12771 22559
rect 12713 22519 12771 22525
rect 12897 22559 12955 22565
rect 12897 22525 12909 22559
rect 12943 22556 12955 22559
rect 13998 22556 14004 22568
rect 12943 22528 14004 22556
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 11256 22488 11284 22519
rect 13998 22516 14004 22528
rect 14056 22516 14062 22568
rect 14292 22556 14320 22584
rect 15562 22556 15568 22568
rect 14292 22528 15568 22556
rect 15562 22516 15568 22528
rect 15620 22556 15626 22568
rect 16666 22556 16672 22568
rect 15620 22528 16672 22556
rect 15620 22516 15626 22528
rect 16666 22516 16672 22528
rect 16724 22556 16730 22568
rect 16761 22559 16819 22565
rect 16761 22556 16773 22559
rect 16724 22528 16773 22556
rect 16724 22516 16730 22528
rect 16761 22525 16773 22528
rect 16807 22556 16819 22559
rect 18509 22559 18567 22565
rect 18509 22556 18521 22559
rect 16807 22528 18521 22556
rect 16807 22525 16819 22528
rect 16761 22519 16819 22525
rect 18509 22525 18521 22528
rect 18555 22525 18567 22559
rect 18509 22519 18567 22525
rect 11977 22491 12035 22497
rect 11977 22488 11989 22491
rect 11256 22460 11989 22488
rect 11977 22457 11989 22460
rect 12023 22488 12035 22491
rect 12434 22488 12440 22500
rect 12023 22460 12440 22488
rect 12023 22457 12035 22460
rect 11977 22451 12035 22457
rect 12434 22448 12440 22460
rect 12492 22448 12498 22500
rect 20824 22488 20852 22587
rect 21008 22556 21036 22587
rect 21450 22584 21456 22636
rect 21508 22624 21514 22636
rect 22756 22624 22784 22664
rect 24670 22652 24676 22704
rect 24728 22652 24734 22704
rect 24762 22652 24768 22704
rect 24820 22652 24826 22704
rect 24854 22652 24860 22704
rect 24912 22692 24918 22704
rect 25516 22692 25544 22732
rect 25590 22720 25596 22772
rect 25648 22760 25654 22772
rect 26142 22760 26148 22772
rect 25648 22732 26148 22760
rect 25648 22720 25654 22732
rect 26142 22720 26148 22732
rect 26200 22720 26206 22772
rect 26234 22720 26240 22772
rect 26292 22760 26298 22772
rect 26292 22732 30420 22760
rect 26292 22720 26298 22732
rect 27890 22692 27896 22704
rect 24912 22664 25176 22692
rect 25516 22664 27896 22692
rect 24912 22652 24918 22664
rect 21508 22596 22784 22624
rect 22824 22627 22882 22633
rect 21508 22584 21514 22596
rect 22824 22593 22836 22627
rect 22870 22624 22882 22627
rect 23106 22624 23112 22636
rect 22870 22596 23112 22624
rect 22870 22593 22882 22596
rect 22824 22587 22882 22593
rect 23106 22584 23112 22596
rect 23164 22584 23170 22636
rect 24581 22627 24639 22633
rect 24581 22593 24593 22627
rect 24627 22624 24639 22627
rect 24780 22624 24808 22652
rect 25041 22627 25099 22633
rect 25041 22624 25053 22627
rect 24627 22596 25053 22624
rect 24627 22593 24639 22596
rect 24581 22587 24639 22593
rect 25041 22593 25053 22596
rect 25087 22593 25099 22627
rect 25148 22624 25176 22664
rect 27890 22652 27896 22664
rect 27948 22652 27954 22704
rect 30282 22652 30288 22704
rect 30340 22652 30346 22704
rect 30392 22692 30420 22732
rect 31754 22720 31760 22772
rect 31812 22760 31818 22772
rect 32490 22760 32496 22772
rect 31812 22732 32496 22760
rect 31812 22720 31818 22732
rect 32490 22720 32496 22732
rect 32548 22720 32554 22772
rect 33410 22720 33416 22772
rect 33468 22720 33474 22772
rect 33502 22720 33508 22772
rect 33560 22760 33566 22772
rect 33560 22732 35204 22760
rect 33560 22720 33566 22732
rect 30392 22664 30774 22692
rect 33226 22652 33232 22704
rect 33284 22692 33290 22704
rect 33284 22664 33718 22692
rect 33284 22652 33290 22664
rect 34882 22652 34888 22704
rect 34940 22652 34946 22704
rect 35176 22692 35204 22732
rect 35250 22720 35256 22772
rect 35308 22720 35314 22772
rect 36170 22720 36176 22772
rect 36228 22760 36234 22772
rect 36449 22763 36507 22769
rect 36449 22760 36461 22763
rect 36228 22732 36461 22760
rect 36228 22720 36234 22732
rect 36449 22729 36461 22732
rect 36495 22729 36507 22763
rect 36449 22723 36507 22729
rect 36541 22763 36599 22769
rect 36541 22729 36553 22763
rect 36587 22760 36599 22763
rect 37182 22760 37188 22772
rect 36587 22732 37188 22760
rect 36587 22729 36599 22732
rect 36541 22723 36599 22729
rect 36262 22692 36268 22704
rect 35176 22664 36268 22692
rect 25498 22624 25504 22636
rect 25148 22596 25504 22624
rect 25041 22587 25099 22593
rect 25498 22584 25504 22596
rect 25556 22624 25562 22636
rect 25556 22596 25728 22624
rect 25556 22584 25562 22596
rect 21008 22528 21588 22556
rect 21082 22488 21088 22500
rect 20824 22460 21088 22488
rect 21082 22448 21088 22460
rect 21140 22448 21146 22500
rect 21560 22488 21588 22528
rect 21818 22516 21824 22568
rect 21876 22516 21882 22568
rect 22370 22516 22376 22568
rect 22428 22556 22434 22568
rect 22557 22559 22615 22565
rect 22557 22556 22569 22559
rect 22428 22528 22569 22556
rect 22428 22516 22434 22528
rect 22557 22525 22569 22528
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 23750 22516 23756 22568
rect 23808 22556 23814 22568
rect 24765 22559 24823 22565
rect 24765 22556 24777 22559
rect 23808 22528 24777 22556
rect 23808 22516 23814 22528
rect 24765 22525 24777 22528
rect 24811 22525 24823 22559
rect 24765 22519 24823 22525
rect 22465 22491 22523 22497
rect 22465 22488 22477 22491
rect 21560 22460 22477 22488
rect 22465 22457 22477 22460
rect 22511 22488 22523 22491
rect 23937 22491 23995 22497
rect 22511 22460 22600 22488
rect 22511 22457 22523 22460
rect 22465 22451 22523 22457
rect 22572 22432 22600 22460
rect 23937 22457 23949 22491
rect 23983 22488 23995 22491
rect 24118 22488 24124 22500
rect 23983 22460 24124 22488
rect 23983 22457 23995 22460
rect 23937 22451 23995 22457
rect 24118 22448 24124 22460
rect 24176 22448 24182 22500
rect 24780 22488 24808 22519
rect 24854 22516 24860 22568
rect 24912 22556 24918 22568
rect 25593 22559 25651 22565
rect 25593 22556 25605 22559
rect 24912 22528 25605 22556
rect 24912 22516 24918 22528
rect 25593 22525 25605 22528
rect 25639 22525 25651 22559
rect 25700 22556 25728 22596
rect 25774 22584 25780 22636
rect 25832 22584 25838 22636
rect 27154 22584 27160 22636
rect 27212 22584 27218 22636
rect 27706 22584 27712 22636
rect 27764 22624 27770 22636
rect 27801 22627 27859 22633
rect 27801 22624 27813 22627
rect 27764 22596 27813 22624
rect 27764 22584 27770 22596
rect 27801 22593 27813 22596
rect 27847 22624 27859 22627
rect 28166 22624 28172 22636
rect 27847 22596 28172 22624
rect 27847 22593 27859 22596
rect 27801 22587 27859 22593
rect 28166 22584 28172 22596
rect 28224 22624 28230 22636
rect 30009 22627 30067 22633
rect 30009 22624 30021 22627
rect 28224 22596 30021 22624
rect 28224 22584 28230 22596
rect 30009 22593 30021 22596
rect 30055 22593 30067 22627
rect 30009 22587 30067 22593
rect 32122 22584 32128 22636
rect 32180 22624 32186 22636
rect 32674 22624 32680 22636
rect 32180 22596 32680 22624
rect 32180 22584 32186 22596
rect 32674 22584 32680 22596
rect 32732 22584 32738 22636
rect 35176 22633 35204 22664
rect 36262 22652 36268 22664
rect 36320 22652 36326 22704
rect 35161 22627 35219 22633
rect 35161 22593 35173 22627
rect 35207 22593 35219 22627
rect 35161 22587 35219 22593
rect 35434 22584 35440 22636
rect 35492 22584 35498 22636
rect 35621 22627 35679 22633
rect 35621 22593 35633 22627
rect 35667 22624 35679 22627
rect 36556 22624 36584 22723
rect 37182 22720 37188 22732
rect 37240 22760 37246 22772
rect 38010 22760 38016 22772
rect 37240 22732 38016 22760
rect 37240 22720 37246 22732
rect 38010 22720 38016 22732
rect 38068 22720 38074 22772
rect 38194 22720 38200 22772
rect 38252 22760 38258 22772
rect 38657 22763 38715 22769
rect 38657 22760 38669 22763
rect 38252 22732 38669 22760
rect 38252 22720 38258 22732
rect 38657 22729 38669 22732
rect 38703 22729 38715 22763
rect 38657 22723 38715 22729
rect 40310 22720 40316 22772
rect 40368 22720 40374 22772
rect 41141 22763 41199 22769
rect 41141 22729 41153 22763
rect 41187 22760 41199 22763
rect 41230 22760 41236 22772
rect 41187 22732 41236 22760
rect 41187 22729 41199 22732
rect 41141 22723 41199 22729
rect 41230 22720 41236 22732
rect 41288 22720 41294 22772
rect 42058 22692 42064 22704
rect 39776 22664 42064 22692
rect 35667 22596 36584 22624
rect 35667 22593 35679 22596
rect 35621 22587 35679 22593
rect 26234 22556 26240 22568
rect 25700 22528 26240 22556
rect 25593 22519 25651 22525
rect 26234 22516 26240 22528
rect 26292 22516 26298 22568
rect 26789 22559 26847 22565
rect 26789 22525 26801 22559
rect 26835 22556 26847 22559
rect 26970 22556 26976 22568
rect 26835 22528 26976 22556
rect 26835 22525 26847 22528
rect 26789 22519 26847 22525
rect 26970 22516 26976 22528
rect 27028 22516 27034 22568
rect 33321 22559 33379 22565
rect 33321 22525 33333 22559
rect 33367 22556 33379 22559
rect 34790 22556 34796 22568
rect 33367 22528 34796 22556
rect 33367 22525 33379 22528
rect 33321 22519 33379 22525
rect 34790 22516 34796 22528
rect 34848 22516 34854 22568
rect 35342 22516 35348 22568
rect 35400 22556 35406 22568
rect 35636 22556 35664 22587
rect 37734 22584 37740 22636
rect 37792 22624 37798 22636
rect 39776 22633 39804 22664
rect 42058 22652 42064 22664
rect 42116 22652 42122 22704
rect 38565 22627 38623 22633
rect 38565 22624 38577 22627
rect 37792 22596 38577 22624
rect 37792 22584 37798 22596
rect 38565 22593 38577 22596
rect 38611 22593 38623 22627
rect 38565 22587 38623 22593
rect 39761 22627 39819 22633
rect 39761 22593 39773 22627
rect 39807 22593 39819 22627
rect 39761 22587 39819 22593
rect 40221 22627 40279 22633
rect 40221 22593 40233 22627
rect 40267 22624 40279 22627
rect 40954 22624 40960 22636
rect 40267 22596 40960 22624
rect 40267 22593 40279 22596
rect 40221 22587 40279 22593
rect 40954 22584 40960 22596
rect 41012 22584 41018 22636
rect 41049 22627 41107 22633
rect 41049 22593 41061 22627
rect 41095 22624 41107 22627
rect 41966 22624 41972 22636
rect 41095 22596 41972 22624
rect 41095 22593 41107 22596
rect 41049 22587 41107 22593
rect 41966 22584 41972 22596
rect 42024 22584 42030 22636
rect 35400 22528 35664 22556
rect 36265 22559 36323 22565
rect 35400 22516 35406 22528
rect 36265 22525 36277 22559
rect 36311 22556 36323 22559
rect 36446 22556 36452 22568
rect 36311 22528 36452 22556
rect 36311 22525 36323 22528
rect 36265 22519 36323 22525
rect 36446 22516 36452 22528
rect 36504 22516 36510 22568
rect 38749 22559 38807 22565
rect 38749 22525 38761 22559
rect 38795 22556 38807 22559
rect 40405 22559 40463 22565
rect 40405 22556 40417 22559
rect 38795 22528 38829 22556
rect 39408 22528 40417 22556
rect 38795 22525 38807 22528
rect 38749 22519 38807 22525
rect 26510 22488 26516 22500
rect 24780 22460 26516 22488
rect 26510 22448 26516 22460
rect 26568 22488 26574 22500
rect 28074 22488 28080 22500
rect 26568 22460 28080 22488
rect 26568 22448 26574 22460
rect 28074 22448 28080 22460
rect 28132 22448 28138 22500
rect 31846 22448 31852 22500
rect 31904 22488 31910 22500
rect 38764 22488 38792 22519
rect 39408 22500 39436 22528
rect 40405 22525 40417 22528
rect 40451 22556 40463 22559
rect 41233 22559 41291 22565
rect 41233 22556 41245 22559
rect 40451 22528 41245 22556
rect 40451 22525 40463 22528
rect 40405 22519 40463 22525
rect 41233 22525 41245 22528
rect 41279 22525 41291 22559
rect 41233 22519 41291 22525
rect 41322 22516 41328 22568
rect 41380 22556 41386 22568
rect 42061 22559 42119 22565
rect 42061 22556 42073 22559
rect 41380 22528 42073 22556
rect 41380 22516 41386 22528
rect 42061 22525 42073 22528
rect 42107 22525 42119 22559
rect 42061 22519 42119 22525
rect 39390 22488 39396 22500
rect 31904 22460 33916 22488
rect 31904 22448 31910 22460
rect 9539 22392 10272 22420
rect 9539 22389 9551 22392
rect 9493 22383 9551 22389
rect 12250 22380 12256 22432
rect 12308 22380 12314 22432
rect 12802 22380 12808 22432
rect 12860 22420 12866 22432
rect 13449 22423 13507 22429
rect 13449 22420 13461 22423
rect 12860 22392 13461 22420
rect 12860 22380 12866 22392
rect 13449 22389 13461 22392
rect 13495 22389 13507 22423
rect 13449 22383 13507 22389
rect 16390 22380 16396 22432
rect 16448 22380 16454 22432
rect 17494 22380 17500 22432
rect 17552 22420 17558 22432
rect 17773 22423 17831 22429
rect 17773 22420 17785 22423
rect 17552 22392 17785 22420
rect 17552 22380 17558 22392
rect 17773 22389 17785 22392
rect 17819 22389 17831 22423
rect 17773 22383 17831 22389
rect 20438 22380 20444 22432
rect 20496 22380 20502 22432
rect 20530 22380 20536 22432
rect 20588 22420 20594 22432
rect 21177 22423 21235 22429
rect 21177 22420 21189 22423
rect 20588 22392 21189 22420
rect 20588 22380 20594 22392
rect 21177 22389 21189 22392
rect 21223 22389 21235 22423
rect 21177 22383 21235 22389
rect 21637 22423 21695 22429
rect 21637 22389 21649 22423
rect 21683 22420 21695 22423
rect 21726 22420 21732 22432
rect 21683 22392 21732 22420
rect 21683 22389 21695 22392
rect 21637 22383 21695 22389
rect 21726 22380 21732 22392
rect 21784 22380 21790 22432
rect 22554 22380 22560 22432
rect 22612 22380 22618 22432
rect 25958 22380 25964 22432
rect 26016 22380 26022 22432
rect 27709 22423 27767 22429
rect 27709 22389 27721 22423
rect 27755 22420 27767 22423
rect 28534 22420 28540 22432
rect 27755 22392 28540 22420
rect 27755 22389 27767 22392
rect 27709 22383 27767 22389
rect 28534 22380 28540 22392
rect 28592 22380 28598 22432
rect 33888 22420 33916 22460
rect 36832 22460 39396 22488
rect 36832 22420 36860 22460
rect 39390 22448 39396 22460
rect 39448 22448 39454 22500
rect 39577 22491 39635 22497
rect 39577 22457 39589 22491
rect 39623 22488 39635 22491
rect 42150 22488 42156 22500
rect 39623 22460 42156 22488
rect 39623 22457 39635 22460
rect 39577 22451 39635 22457
rect 42150 22448 42156 22460
rect 42208 22448 42214 22500
rect 33888 22392 36860 22420
rect 36906 22380 36912 22432
rect 36964 22380 36970 22432
rect 37550 22380 37556 22432
rect 37608 22420 37614 22432
rect 38197 22423 38255 22429
rect 38197 22420 38209 22423
rect 37608 22392 38209 22420
rect 37608 22380 37614 22392
rect 38197 22389 38209 22392
rect 38243 22389 38255 22423
rect 38197 22383 38255 22389
rect 39853 22423 39911 22429
rect 39853 22389 39865 22423
rect 39899 22420 39911 22423
rect 40126 22420 40132 22432
rect 39899 22392 40132 22420
rect 39899 22389 39911 22392
rect 39853 22383 39911 22389
rect 40126 22380 40132 22392
rect 40184 22380 40190 22432
rect 40678 22380 40684 22432
rect 40736 22380 40742 22432
rect 40954 22380 40960 22432
rect 41012 22420 41018 22432
rect 41138 22420 41144 22432
rect 41012 22392 41144 22420
rect 41012 22380 41018 22392
rect 41138 22380 41144 22392
rect 41196 22420 41202 22432
rect 41509 22423 41567 22429
rect 41509 22420 41521 22423
rect 41196 22392 41521 22420
rect 41196 22380 41202 22392
rect 41509 22389 41521 22392
rect 41555 22389 41567 22423
rect 41509 22383 41567 22389
rect 1104 22330 42504 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 42504 22330
rect 1104 22256 42504 22278
rect 5534 22176 5540 22228
rect 5592 22176 5598 22228
rect 7650 22176 7656 22228
rect 7708 22216 7714 22228
rect 7745 22219 7803 22225
rect 7745 22216 7757 22219
rect 7708 22188 7757 22216
rect 7708 22176 7714 22188
rect 7745 22185 7757 22188
rect 7791 22185 7803 22219
rect 7745 22179 7803 22185
rect 14458 22176 14464 22228
rect 14516 22216 14522 22228
rect 14737 22219 14795 22225
rect 14737 22216 14749 22219
rect 14516 22188 14749 22216
rect 14516 22176 14522 22188
rect 14737 22185 14749 22188
rect 14783 22185 14795 22219
rect 14737 22179 14795 22185
rect 15102 22176 15108 22228
rect 15160 22216 15166 22228
rect 16390 22216 16396 22228
rect 15160 22188 16396 22216
rect 15160 22176 15166 22188
rect 5552 22148 5580 22176
rect 7098 22148 7104 22160
rect 5368 22120 7104 22148
rect 3234 22040 3240 22092
rect 3292 22080 3298 22092
rect 3881 22083 3939 22089
rect 3881 22080 3893 22083
rect 3292 22052 3893 22080
rect 3292 22040 3298 22052
rect 3881 22049 3893 22052
rect 3927 22049 3939 22083
rect 3881 22043 3939 22049
rect 1394 21972 1400 22024
rect 1452 21972 1458 22024
rect 4246 21972 4252 22024
rect 4304 21972 4310 22024
rect 5368 21944 5396 22120
rect 7098 22108 7104 22120
rect 7156 22108 7162 22160
rect 7377 22083 7435 22089
rect 6748 22052 7144 22080
rect 6362 21972 6368 22024
rect 6420 22012 6426 22024
rect 6748 22012 6776 22052
rect 6420 21984 6776 22012
rect 6420 21972 6426 21984
rect 6822 21972 6828 22024
rect 6880 21972 6886 22024
rect 7116 22021 7144 22052
rect 7377 22049 7389 22083
rect 7423 22080 7435 22083
rect 7837 22083 7895 22089
rect 7837 22080 7849 22083
rect 7423 22052 7849 22080
rect 7423 22049 7435 22052
rect 7377 22043 7435 22049
rect 7837 22049 7849 22052
rect 7883 22049 7895 22083
rect 7837 22043 7895 22049
rect 9125 22083 9183 22089
rect 9125 22049 9137 22083
rect 9171 22080 9183 22083
rect 10134 22080 10140 22092
rect 9171 22052 10140 22080
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 7282 21972 7288 22024
rect 7340 21972 7346 22024
rect 7466 21972 7472 22024
rect 7524 21972 7530 22024
rect 7742 21972 7748 22024
rect 7800 21972 7806 22024
rect 8481 22015 8539 22021
rect 8481 21981 8493 22015
rect 8527 22012 8539 22015
rect 8846 22012 8852 22024
rect 8527 21984 8852 22012
rect 8527 21981 8539 21984
rect 8481 21975 8539 21981
rect 8846 21972 8852 21984
rect 8904 21972 8910 22024
rect 11606 21972 11612 22024
rect 11664 22012 11670 22024
rect 12802 22021 12808 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 11664 21984 12541 22012
rect 11664 21972 11670 21984
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 12796 21975 12808 22021
rect 12802 21972 12808 21975
rect 12860 21972 12866 22024
rect 15212 22021 15240 22188
rect 16390 22176 16396 22188
rect 16448 22176 16454 22228
rect 17494 22225 17500 22228
rect 17484 22219 17500 22225
rect 17484 22185 17496 22219
rect 17484 22179 17500 22185
rect 17494 22176 17500 22179
rect 17552 22176 17558 22228
rect 18230 22176 18236 22228
rect 18288 22216 18294 22228
rect 18969 22219 19027 22225
rect 18969 22216 18981 22219
rect 18288 22188 18981 22216
rect 18288 22176 18294 22188
rect 18969 22185 18981 22188
rect 19015 22185 19027 22219
rect 18969 22179 19027 22185
rect 20622 22176 20628 22228
rect 20680 22216 20686 22228
rect 20680 22188 23060 22216
rect 20680 22176 20686 22188
rect 16117 22151 16175 22157
rect 16117 22117 16129 22151
rect 16163 22148 16175 22151
rect 16942 22148 16948 22160
rect 16163 22120 16948 22148
rect 16163 22117 16175 22120
rect 16117 22111 16175 22117
rect 16942 22108 16948 22120
rect 17000 22108 17006 22160
rect 23032 22148 23060 22188
rect 23106 22176 23112 22228
rect 23164 22176 23170 22228
rect 25774 22216 25780 22228
rect 23216 22188 25780 22216
rect 23216 22148 23244 22188
rect 25774 22176 25780 22188
rect 25832 22216 25838 22228
rect 34054 22216 34060 22228
rect 25832 22188 34060 22216
rect 25832 22176 25838 22188
rect 34054 22176 34060 22188
rect 34112 22176 34118 22228
rect 34606 22176 34612 22228
rect 34664 22216 34670 22228
rect 34701 22219 34759 22225
rect 34701 22216 34713 22219
rect 34664 22188 34713 22216
rect 34664 22176 34670 22188
rect 34701 22185 34713 22188
rect 34747 22185 34759 22219
rect 34701 22179 34759 22185
rect 36528 22219 36586 22225
rect 36528 22185 36540 22219
rect 36574 22216 36586 22219
rect 36906 22216 36912 22228
rect 36574 22188 36912 22216
rect 36574 22185 36586 22188
rect 36528 22179 36586 22185
rect 36906 22176 36912 22188
rect 36964 22176 36970 22228
rect 41233 22219 41291 22225
rect 41233 22185 41245 22219
rect 41279 22216 41291 22219
rect 41322 22216 41328 22228
rect 41279 22188 41328 22216
rect 41279 22185 41291 22188
rect 41233 22179 41291 22185
rect 41322 22176 41328 22188
rect 41380 22176 41386 22228
rect 24026 22148 24032 22160
rect 23032 22120 23244 22148
rect 23584 22120 24032 22148
rect 15470 22040 15476 22092
rect 15528 22080 15534 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 15528 22052 15761 22080
rect 15528 22040 15534 22052
rect 15749 22049 15761 22052
rect 15795 22049 15807 22083
rect 16298 22080 16304 22092
rect 15749 22043 15807 22049
rect 15948 22052 16304 22080
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 15197 22015 15255 22021
rect 15197 21981 15209 22015
rect 15243 21981 15255 22015
rect 15197 21975 15255 21981
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 22012 15347 22015
rect 15335 21984 15516 22012
rect 15335 21981 15347 21984
rect 15289 21975 15347 21981
rect 5290 21916 5396 21944
rect 5902 21904 5908 21956
rect 5960 21944 5966 21956
rect 6454 21944 6460 21956
rect 5960 21916 6460 21944
rect 5960 21904 5966 21916
rect 6454 21904 6460 21916
rect 6512 21904 6518 21956
rect 6733 21947 6791 21953
rect 6733 21913 6745 21947
rect 6779 21944 6791 21947
rect 9030 21944 9036 21956
rect 6779 21916 9036 21944
rect 6779 21913 6791 21916
rect 6733 21907 6791 21913
rect 9030 21904 9036 21916
rect 9088 21904 9094 21956
rect 9398 21904 9404 21956
rect 9456 21904 9462 21956
rect 9508 21916 9890 21944
rect 1302 21836 1308 21888
rect 1360 21876 1366 21888
rect 5718 21885 5724 21888
rect 1581 21879 1639 21885
rect 1581 21876 1593 21879
rect 1360 21848 1593 21876
rect 1360 21836 1366 21848
rect 1581 21845 1593 21848
rect 1627 21845 1639 21879
rect 1581 21839 1639 21845
rect 5675 21879 5724 21885
rect 5675 21845 5687 21879
rect 5721 21845 5724 21879
rect 5675 21839 5724 21845
rect 5718 21836 5724 21839
rect 5776 21876 5782 21888
rect 6178 21876 6184 21888
rect 5776 21848 6184 21876
rect 5776 21836 5782 21848
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 6914 21836 6920 21888
rect 6972 21836 6978 21888
rect 7006 21836 7012 21888
rect 7064 21876 7070 21888
rect 7561 21879 7619 21885
rect 7561 21876 7573 21879
rect 7064 21848 7573 21876
rect 7064 21836 7070 21848
rect 7561 21845 7573 21848
rect 7607 21876 7619 21879
rect 7926 21876 7932 21888
rect 7607 21848 7932 21876
rect 7607 21845 7619 21848
rect 7561 21839 7619 21845
rect 7926 21836 7932 21848
rect 7984 21876 7990 21888
rect 9508 21876 9536 21916
rect 11146 21904 11152 21956
rect 11204 21904 11210 21956
rect 7984 21848 9536 21876
rect 13909 21879 13967 21885
rect 7984 21836 7990 21848
rect 13909 21845 13921 21879
rect 13955 21876 13967 21879
rect 14108 21876 14136 21975
rect 15378 21904 15384 21956
rect 15436 21904 15442 21956
rect 15488 21944 15516 21984
rect 15562 21972 15568 22024
rect 15620 21972 15626 22024
rect 15654 21972 15660 22024
rect 15712 21972 15718 22024
rect 15948 22021 15976 22052
rect 16298 22040 16304 22052
rect 16356 22040 16362 22092
rect 16666 22040 16672 22092
rect 16724 22080 16730 22092
rect 23584 22089 23612 22120
rect 24026 22108 24032 22120
rect 24084 22108 24090 22160
rect 27890 22108 27896 22160
rect 27948 22148 27954 22160
rect 31754 22148 31760 22160
rect 27948 22120 31760 22148
rect 27948 22108 27954 22120
rect 17221 22083 17279 22089
rect 17221 22080 17233 22083
rect 16724 22052 17233 22080
rect 16724 22040 16730 22052
rect 17221 22049 17233 22052
rect 17267 22080 17279 22083
rect 23569 22083 23627 22089
rect 17267 22052 18920 22080
rect 17267 22049 17279 22052
rect 17221 22043 17279 22049
rect 18892 22024 18920 22052
rect 23569 22049 23581 22083
rect 23615 22080 23627 22083
rect 23615 22052 23649 22080
rect 23615 22049 23627 22052
rect 23569 22043 23627 22049
rect 23750 22040 23756 22092
rect 23808 22040 23814 22092
rect 24118 22040 24124 22092
rect 24176 22080 24182 22092
rect 24949 22083 25007 22089
rect 24949 22080 24961 22083
rect 24176 22052 24961 22080
rect 24176 22040 24182 22052
rect 24949 22049 24961 22052
rect 24995 22049 25007 22083
rect 30116 22080 30144 22120
rect 31754 22108 31760 22120
rect 31812 22108 31818 22160
rect 30193 22083 30251 22089
rect 30193 22080 30205 22083
rect 30116 22052 30205 22080
rect 24949 22043 25007 22049
rect 30193 22049 30205 22052
rect 30239 22049 30251 22083
rect 30193 22043 30251 22049
rect 31202 22040 31208 22092
rect 31260 22080 31266 22092
rect 31260 22052 31708 22080
rect 31260 22040 31266 22052
rect 15933 22015 15991 22021
rect 15933 21981 15945 22015
rect 15979 21981 15991 22015
rect 15933 21975 15991 21981
rect 16209 22015 16267 22021
rect 16209 21981 16221 22015
rect 16255 22012 16267 22015
rect 16390 22012 16396 22024
rect 16255 21984 16396 22012
rect 16255 21981 16267 21984
rect 16209 21975 16267 21981
rect 16390 21972 16396 21984
rect 16448 22012 16454 22024
rect 16448 21984 16988 22012
rect 16448 21972 16454 21984
rect 16850 21944 16856 21956
rect 15488 21916 16856 21944
rect 16850 21904 16856 21916
rect 16908 21904 16914 21956
rect 13955 21848 14136 21876
rect 13955 21845 13967 21848
rect 13909 21839 13967 21845
rect 15010 21836 15016 21888
rect 15068 21836 15074 21888
rect 16298 21836 16304 21888
rect 16356 21836 16362 21888
rect 16960 21876 16988 21984
rect 18874 21972 18880 22024
rect 18932 22012 18938 22024
rect 19981 22015 20039 22021
rect 19981 22012 19993 22015
rect 18932 21984 19993 22012
rect 18932 21972 18938 21984
rect 19981 21981 19993 21984
rect 20027 21981 20039 22015
rect 19981 21975 20039 21981
rect 21450 21972 21456 22024
rect 21508 21972 21514 22024
rect 21726 22021 21732 22024
rect 21720 21975 21732 22021
rect 21726 21972 21732 21975
rect 21784 21972 21790 22024
rect 23198 21972 23204 22024
rect 23256 22012 23262 22024
rect 23937 22015 23995 22021
rect 23937 22012 23949 22015
rect 23256 21984 23949 22012
rect 23256 21972 23262 21984
rect 23937 21981 23949 21984
rect 23983 22012 23995 22015
rect 23983 21984 25084 22012
rect 23983 21981 23995 21984
rect 23937 21975 23995 21981
rect 18506 21904 18512 21956
rect 18564 21904 18570 21956
rect 20248 21947 20306 21953
rect 20248 21913 20260 21947
rect 20294 21944 20306 21947
rect 20438 21944 20444 21956
rect 20294 21916 20444 21944
rect 20294 21913 20306 21916
rect 20248 21907 20306 21913
rect 20438 21904 20444 21916
rect 20496 21904 20502 21956
rect 24397 21947 24455 21953
rect 24397 21944 24409 21947
rect 23492 21916 24409 21944
rect 18138 21876 18144 21888
rect 16960 21848 18144 21876
rect 18138 21836 18144 21848
rect 18196 21876 18202 21888
rect 20622 21876 20628 21888
rect 18196 21848 20628 21876
rect 18196 21836 18202 21848
rect 20622 21836 20628 21848
rect 20680 21836 20686 21888
rect 20990 21836 20996 21888
rect 21048 21876 21054 21888
rect 21361 21879 21419 21885
rect 21361 21876 21373 21879
rect 21048 21848 21373 21876
rect 21048 21836 21054 21848
rect 21361 21845 21373 21848
rect 21407 21876 21419 21879
rect 21818 21876 21824 21888
rect 21407 21848 21824 21876
rect 21407 21845 21419 21848
rect 21361 21839 21419 21845
rect 21818 21836 21824 21848
rect 21876 21836 21882 21888
rect 22830 21836 22836 21888
rect 22888 21836 22894 21888
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 23492 21885 23520 21916
rect 24397 21913 24409 21916
rect 24443 21913 24455 21947
rect 24397 21907 24455 21913
rect 23477 21879 23535 21885
rect 23477 21876 23489 21879
rect 23348 21848 23489 21876
rect 23348 21836 23354 21848
rect 23477 21845 23489 21848
rect 23523 21845 23535 21879
rect 23477 21839 23535 21845
rect 24121 21879 24179 21885
rect 24121 21845 24133 21879
rect 24167 21876 24179 21879
rect 24946 21876 24952 21888
rect 24167 21848 24952 21876
rect 24167 21845 24179 21848
rect 24121 21839 24179 21845
rect 24946 21836 24952 21848
rect 25004 21836 25010 21888
rect 25056 21876 25084 21984
rect 25130 21972 25136 22024
rect 25188 22012 25194 22024
rect 26605 22015 26663 22021
rect 26605 22012 26617 22015
rect 25188 21984 26617 22012
rect 25188 21972 25194 21984
rect 26605 21981 26617 21984
rect 26651 22012 26663 22015
rect 26651 21984 28212 22012
rect 26651 21981 26663 21984
rect 26605 21975 26663 21981
rect 26988 21956 27016 21984
rect 28184 21956 28212 21984
rect 28810 21972 28816 22024
rect 28868 22012 28874 22024
rect 28868 21984 30236 22012
rect 28868 21972 28874 21984
rect 25400 21947 25458 21953
rect 25400 21913 25412 21947
rect 25446 21944 25458 21947
rect 25590 21944 25596 21956
rect 25446 21916 25596 21944
rect 25446 21913 25458 21916
rect 25400 21907 25458 21913
rect 25590 21904 25596 21916
rect 25648 21904 25654 21956
rect 26418 21904 26424 21956
rect 26476 21944 26482 21956
rect 26850 21947 26908 21953
rect 26850 21944 26862 21947
rect 26476 21916 26862 21944
rect 26476 21904 26482 21916
rect 26850 21913 26862 21916
rect 26896 21913 26908 21947
rect 26850 21907 26908 21913
rect 26970 21904 26976 21956
rect 27028 21904 27034 21956
rect 28166 21904 28172 21956
rect 28224 21944 28230 21956
rect 28261 21947 28319 21953
rect 28261 21944 28273 21947
rect 28224 21916 28273 21944
rect 28224 21904 28230 21916
rect 28261 21913 28273 21916
rect 28307 21944 28319 21947
rect 28442 21944 28448 21956
rect 28307 21916 28448 21944
rect 28307 21913 28319 21916
rect 28261 21907 28319 21913
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 28994 21904 29000 21956
rect 29052 21904 29058 21956
rect 30009 21947 30067 21953
rect 30009 21913 30021 21947
rect 30055 21944 30067 21947
rect 30098 21944 30104 21956
rect 30055 21916 30104 21944
rect 30055 21913 30067 21916
rect 30009 21907 30067 21913
rect 30098 21904 30104 21916
rect 30156 21904 30162 21956
rect 30208 21944 30236 21984
rect 30926 21972 30932 22024
rect 30984 21972 30990 22024
rect 31297 22015 31355 22021
rect 31297 21981 31309 22015
rect 31343 21981 31355 22015
rect 31297 21975 31355 21981
rect 31312 21944 31340 21975
rect 31386 21972 31392 22024
rect 31444 21972 31450 22024
rect 31680 22021 31708 22052
rect 34790 22040 34796 22092
rect 34848 22080 34854 22092
rect 34848 22052 35296 22080
rect 34848 22040 34854 22052
rect 31665 22015 31723 22021
rect 31665 21981 31677 22015
rect 31711 21981 31723 22015
rect 31665 21975 31723 21981
rect 32122 21972 32128 22024
rect 32180 21972 32186 22024
rect 33134 22012 33140 22024
rect 32324 21984 33140 22012
rect 30208 21916 31340 21944
rect 25682 21876 25688 21888
rect 25056 21848 25688 21876
rect 25682 21836 25688 21848
rect 25740 21836 25746 21888
rect 26513 21879 26571 21885
rect 26513 21845 26525 21879
rect 26559 21876 26571 21879
rect 26602 21876 26608 21888
rect 26559 21848 26608 21876
rect 26559 21845 26571 21848
rect 26513 21839 26571 21845
rect 26602 21836 26608 21848
rect 26660 21836 26666 21888
rect 27062 21836 27068 21888
rect 27120 21876 27126 21888
rect 27985 21879 28043 21885
rect 27985 21876 27997 21879
rect 27120 21848 27997 21876
rect 27120 21836 27126 21848
rect 27985 21845 27997 21848
rect 28031 21845 28043 21879
rect 27985 21839 28043 21845
rect 29546 21836 29552 21888
rect 29604 21836 29610 21888
rect 29822 21836 29828 21888
rect 29880 21876 29886 21888
rect 29917 21879 29975 21885
rect 29917 21876 29929 21879
rect 29880 21848 29929 21876
rect 29880 21836 29886 21848
rect 29917 21845 29929 21848
rect 29963 21876 29975 21879
rect 30377 21879 30435 21885
rect 30377 21876 30389 21879
rect 29963 21848 30389 21876
rect 29963 21845 29975 21848
rect 29917 21839 29975 21845
rect 30377 21845 30389 21848
rect 30423 21845 30435 21879
rect 30377 21839 30435 21845
rect 31110 21836 31116 21888
rect 31168 21836 31174 21888
rect 31312 21876 31340 21916
rect 31478 21904 31484 21956
rect 31536 21904 31542 21956
rect 32324 21944 32352 21984
rect 33134 21972 33140 21984
rect 33192 21972 33198 22024
rect 34149 22015 34207 22021
rect 34149 21981 34161 22015
rect 34195 21981 34207 22015
rect 34149 21975 34207 21981
rect 32398 21953 32404 21956
rect 31726 21916 32352 21944
rect 31726 21876 31754 21916
rect 32392 21907 32404 21953
rect 32398 21904 32404 21907
rect 32456 21904 32462 21956
rect 33410 21904 33416 21956
rect 33468 21944 33474 21956
rect 33597 21947 33655 21953
rect 33597 21944 33609 21947
rect 33468 21916 33609 21944
rect 33468 21904 33474 21916
rect 33597 21913 33609 21916
rect 33643 21913 33655 21947
rect 33597 21907 33655 21913
rect 31312 21848 31754 21876
rect 32490 21836 32496 21888
rect 32548 21876 32554 21888
rect 33042 21876 33048 21888
rect 32548 21848 33048 21876
rect 32548 21836 32554 21848
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 33502 21836 33508 21888
rect 33560 21876 33566 21888
rect 34164 21876 34192 21975
rect 34422 21972 34428 22024
rect 34480 22012 34486 22024
rect 35268 22021 35296 22052
rect 36262 22040 36268 22092
rect 36320 22080 36326 22092
rect 36538 22080 36544 22092
rect 36320 22052 36544 22080
rect 36320 22040 36326 22052
rect 36538 22040 36544 22052
rect 36596 22040 36602 22092
rect 38010 22040 38016 22092
rect 38068 22040 38074 22092
rect 41966 22040 41972 22092
rect 42024 22040 42030 22092
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 34480 21984 34897 22012
rect 34480 21972 34486 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 35253 22015 35311 22021
rect 35253 21981 35265 22015
rect 35299 21981 35311 22015
rect 38746 22012 38752 22024
rect 37674 21984 38752 22012
rect 35253 21975 35311 21981
rect 38746 21972 38752 21984
rect 38804 21972 38810 22024
rect 39025 22015 39083 22021
rect 39025 21981 39037 22015
rect 39071 22012 39083 22015
rect 39853 22015 39911 22021
rect 39853 22012 39865 22015
rect 39071 21984 39865 22012
rect 39071 21981 39083 21984
rect 39025 21975 39083 21981
rect 39853 21981 39865 21984
rect 39899 22012 39911 22015
rect 40402 22012 40408 22024
rect 39899 21984 40408 22012
rect 39899 21981 39911 21984
rect 39853 21975 39911 21981
rect 40402 21972 40408 21984
rect 40460 21972 40466 22024
rect 41322 21972 41328 22024
rect 41380 21972 41386 22024
rect 34698 21904 34704 21956
rect 34756 21944 34762 21956
rect 34977 21947 35035 21953
rect 34977 21944 34989 21947
rect 34756 21916 34989 21944
rect 34756 21904 34762 21916
rect 34977 21913 34989 21916
rect 35023 21913 35035 21947
rect 34977 21907 35035 21913
rect 35066 21904 35072 21956
rect 35124 21904 35130 21956
rect 38194 21904 38200 21956
rect 38252 21904 38258 21956
rect 40126 21953 40132 21956
rect 40120 21907 40132 21953
rect 40126 21904 40132 21907
rect 40184 21904 40190 21956
rect 33560 21848 34192 21876
rect 33560 21836 33566 21848
rect 1104 21786 42504 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 42504 21786
rect 1104 21712 42504 21734
rect 4433 21675 4491 21681
rect 4433 21641 4445 21675
rect 4479 21672 4491 21675
rect 4706 21672 4712 21684
rect 4479 21644 4712 21672
rect 4479 21641 4491 21644
rect 4433 21635 4491 21641
rect 4706 21632 4712 21644
rect 4764 21632 4770 21684
rect 5810 21672 5816 21684
rect 5184 21644 5816 21672
rect 4246 21564 4252 21616
rect 4304 21604 4310 21616
rect 5077 21607 5135 21613
rect 5077 21604 5089 21607
rect 4304 21576 5089 21604
rect 4304 21564 4310 21576
rect 5077 21573 5089 21576
rect 5123 21573 5135 21607
rect 5077 21567 5135 21573
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21505 4675 21539
rect 4617 21499 4675 21505
rect 4709 21539 4767 21545
rect 4709 21505 4721 21539
rect 4755 21536 4767 21539
rect 4798 21536 4804 21548
rect 4755 21508 4804 21536
rect 4755 21505 4767 21508
rect 4709 21499 4767 21505
rect 3142 21428 3148 21480
rect 3200 21428 3206 21480
rect 4632 21468 4660 21499
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 4893 21539 4951 21545
rect 4893 21505 4905 21539
rect 4939 21505 4951 21539
rect 4893 21499 4951 21505
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21536 5043 21539
rect 5184 21536 5212 21644
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 6822 21632 6828 21684
rect 6880 21672 6886 21684
rect 8297 21675 8355 21681
rect 8297 21672 8309 21675
rect 6880 21644 8309 21672
rect 6880 21632 6886 21644
rect 8297 21641 8309 21644
rect 8343 21641 8355 21675
rect 8297 21635 8355 21641
rect 9398 21632 9404 21684
rect 9456 21672 9462 21684
rect 9585 21675 9643 21681
rect 9585 21672 9597 21675
rect 9456 21644 9597 21672
rect 9456 21632 9462 21644
rect 9585 21641 9597 21644
rect 9631 21641 9643 21675
rect 9585 21635 9643 21641
rect 12986 21632 12992 21684
rect 13044 21632 13050 21684
rect 15562 21632 15568 21684
rect 15620 21632 15626 21684
rect 17037 21675 17095 21681
rect 17037 21641 17049 21675
rect 17083 21672 17095 21675
rect 17218 21672 17224 21684
rect 17083 21644 17224 21672
rect 17083 21641 17095 21644
rect 17037 21635 17095 21641
rect 17218 21632 17224 21644
rect 17276 21672 17282 21684
rect 21358 21672 21364 21684
rect 17276 21644 21364 21672
rect 17276 21632 17282 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 22281 21675 22339 21681
rect 22281 21641 22293 21675
rect 22327 21672 22339 21675
rect 22646 21672 22652 21684
rect 22327 21644 22652 21672
rect 22327 21641 22339 21644
rect 22281 21635 22339 21641
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 24854 21632 24860 21684
rect 24912 21632 24918 21684
rect 25590 21632 25596 21684
rect 25648 21632 25654 21684
rect 25682 21632 25688 21684
rect 25740 21672 25746 21684
rect 25740 21644 27660 21672
rect 25740 21632 25746 21644
rect 5718 21604 5724 21616
rect 5368 21576 5724 21604
rect 5031 21508 5212 21536
rect 5031 21505 5043 21508
rect 4985 21499 5043 21505
rect 4908 21468 4936 21499
rect 5258 21496 5264 21548
rect 5316 21496 5322 21548
rect 5368 21545 5396 21576
rect 5718 21564 5724 21576
rect 5776 21564 5782 21616
rect 7098 21564 7104 21616
rect 7156 21564 7162 21616
rect 9217 21607 9275 21613
rect 9217 21604 9229 21607
rect 7852 21576 9229 21604
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21505 5411 21539
rect 5353 21499 5411 21505
rect 5534 21496 5540 21548
rect 5592 21496 5598 21548
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 5552 21468 5580 21496
rect 4632 21440 4752 21468
rect 4908 21440 5580 21468
rect 4724 21400 4752 21440
rect 5258 21400 5264 21412
rect 4724 21372 5264 21400
rect 5258 21360 5264 21372
rect 5316 21360 5322 21412
rect 5920 21400 5948 21499
rect 6181 21471 6239 21477
rect 6181 21437 6193 21471
rect 6227 21468 6239 21471
rect 6270 21468 6276 21480
rect 6227 21440 6276 21468
rect 6227 21437 6239 21440
rect 6181 21431 6239 21437
rect 6270 21428 6276 21440
rect 6328 21428 6334 21480
rect 6365 21471 6423 21477
rect 6365 21437 6377 21471
rect 6411 21468 6423 21471
rect 6638 21468 6644 21480
rect 6411 21440 6644 21468
rect 6411 21437 6423 21440
rect 6365 21431 6423 21437
rect 6638 21428 6644 21440
rect 6696 21428 6702 21480
rect 6730 21428 6736 21480
rect 6788 21428 6794 21480
rect 7282 21428 7288 21480
rect 7340 21468 7346 21480
rect 7852 21468 7880 21576
rect 9217 21573 9229 21576
rect 9263 21573 9275 21607
rect 9217 21567 9275 21573
rect 9309 21607 9367 21613
rect 9309 21573 9321 21607
rect 9355 21604 9367 21607
rect 11146 21604 11152 21616
rect 9355 21576 11152 21604
rect 9355 21573 9367 21576
rect 9309 21567 9367 21573
rect 11146 21564 11152 21576
rect 11204 21564 11210 21616
rect 11876 21607 11934 21613
rect 11876 21573 11888 21607
rect 11922 21604 11934 21607
rect 12250 21604 12256 21616
rect 11922 21576 12256 21604
rect 11922 21573 11934 21576
rect 11876 21567 11934 21573
rect 12250 21564 12256 21576
rect 12308 21564 12314 21616
rect 16574 21564 16580 21616
rect 16632 21604 16638 21616
rect 16761 21607 16819 21613
rect 16761 21604 16773 21607
rect 16632 21576 16773 21604
rect 16632 21564 16638 21576
rect 16761 21573 16773 21576
rect 16807 21573 16819 21607
rect 16761 21567 16819 21573
rect 16942 21564 16948 21616
rect 17000 21604 17006 21616
rect 17313 21607 17371 21613
rect 17313 21604 17325 21607
rect 17000 21576 17325 21604
rect 17000 21564 17006 21576
rect 17313 21573 17325 21576
rect 17359 21573 17371 21607
rect 20530 21604 20536 21616
rect 17313 21567 17371 21573
rect 17420 21576 20536 21604
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 9401 21539 9459 21545
rect 9401 21505 9413 21539
rect 9447 21505 9459 21539
rect 9401 21499 9459 21505
rect 7340 21440 7880 21468
rect 7340 21428 7346 21440
rect 8846 21428 8852 21480
rect 8904 21428 8910 21480
rect 8938 21428 8944 21480
rect 8996 21468 9002 21480
rect 9416 21468 9444 21499
rect 11606 21496 11612 21548
rect 11664 21496 11670 21548
rect 15010 21496 15016 21548
rect 15068 21536 15074 21548
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 15068 21508 15301 21536
rect 15068 21496 15074 21508
rect 15289 21505 15301 21508
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15378 21496 15384 21548
rect 15436 21536 15442 21548
rect 15436 21508 16252 21536
rect 15436 21496 15442 21508
rect 8996 21440 9444 21468
rect 8996 21428 9002 21440
rect 16114 21428 16120 21480
rect 16172 21428 16178 21480
rect 16224 21468 16252 21508
rect 16298 21496 16304 21548
rect 16356 21536 16362 21548
rect 17420 21536 17448 21576
rect 20530 21564 20536 21576
rect 20588 21564 20594 21616
rect 23198 21604 23204 21616
rect 21100 21576 23204 21604
rect 21100 21548 21128 21576
rect 23198 21564 23204 21576
rect 23256 21564 23262 21616
rect 23744 21607 23802 21613
rect 23744 21573 23756 21607
rect 23790 21604 23802 21607
rect 24210 21604 24216 21616
rect 23790 21576 24216 21604
rect 23790 21573 23802 21576
rect 23744 21567 23802 21573
rect 24210 21564 24216 21576
rect 24268 21564 24274 21616
rect 25314 21564 25320 21616
rect 25372 21564 25378 21616
rect 16356 21508 17448 21536
rect 16356 21496 16362 21508
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18506 21536 18512 21548
rect 18104 21508 18512 21536
rect 18104 21496 18110 21508
rect 18506 21496 18512 21508
rect 18564 21496 18570 21548
rect 18874 21496 18880 21548
rect 18932 21496 18938 21548
rect 19150 21545 19156 21548
rect 19144 21499 19156 21545
rect 19150 21496 19156 21499
rect 19208 21496 19214 21548
rect 21082 21536 21088 21548
rect 20180 21508 21088 21536
rect 17497 21471 17555 21477
rect 17497 21468 17509 21471
rect 16224 21440 17509 21468
rect 17497 21437 17509 21440
rect 17543 21468 17555 21471
rect 17954 21468 17960 21480
rect 17543 21440 17960 21468
rect 17543 21437 17555 21440
rect 17497 21431 17555 21437
rect 17954 21428 17960 21440
rect 18012 21428 18018 21480
rect 5920 21372 6408 21400
rect 2590 21292 2596 21344
rect 2648 21292 2654 21344
rect 5994 21292 6000 21344
rect 6052 21292 6058 21344
rect 6089 21335 6147 21341
rect 6089 21301 6101 21335
rect 6135 21332 6147 21335
rect 6178 21332 6184 21344
rect 6135 21304 6184 21332
rect 6135 21301 6147 21304
rect 6089 21295 6147 21301
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 6380 21332 6408 21372
rect 7558 21332 7564 21344
rect 6380 21304 7564 21332
rect 7558 21292 7564 21304
rect 7616 21332 7622 21344
rect 8159 21335 8217 21341
rect 8159 21332 8171 21335
rect 7616 21304 8171 21332
rect 7616 21292 7622 21304
rect 8159 21301 8171 21304
rect 8205 21301 8217 21335
rect 8159 21295 8217 21301
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 14737 21335 14795 21341
rect 14737 21332 14749 21335
rect 14424 21304 14749 21332
rect 14424 21292 14430 21304
rect 14737 21301 14749 21304
rect 14783 21301 14795 21335
rect 14737 21295 14795 21301
rect 17954 21292 17960 21344
rect 18012 21332 18018 21344
rect 20180 21332 20208 21508
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 22189 21539 22247 21545
rect 22189 21505 22201 21539
rect 22235 21536 22247 21539
rect 22278 21536 22284 21548
rect 22235 21508 22284 21536
rect 22235 21505 22247 21508
rect 22189 21499 22247 21505
rect 22278 21496 22284 21508
rect 22336 21536 22342 21548
rect 25041 21539 25099 21545
rect 22336 21508 22508 21536
rect 22336 21496 22342 21508
rect 20993 21471 21051 21477
rect 20993 21468 21005 21471
rect 20272 21440 21005 21468
rect 20272 21409 20300 21440
rect 20993 21437 21005 21440
rect 21039 21468 21051 21471
rect 21174 21468 21180 21480
rect 21039 21440 21180 21468
rect 21039 21437 21051 21440
rect 20993 21431 21051 21437
rect 21174 21428 21180 21440
rect 21232 21428 21238 21480
rect 22373 21471 22431 21477
rect 22373 21437 22385 21471
rect 22419 21437 22431 21471
rect 22480 21468 22508 21508
rect 25041 21505 25053 21539
rect 25087 21536 25099 21539
rect 25130 21536 25136 21548
rect 25087 21508 25136 21536
rect 25087 21505 25099 21508
rect 25041 21499 25099 21505
rect 25130 21496 25136 21508
rect 25188 21496 25194 21548
rect 25222 21496 25228 21548
rect 25280 21496 25286 21548
rect 25409 21539 25467 21545
rect 25409 21505 25421 21539
rect 25455 21536 25467 21539
rect 25958 21536 25964 21548
rect 25455 21508 25964 21536
rect 25455 21505 25467 21508
rect 25409 21499 25467 21505
rect 25958 21496 25964 21508
rect 26016 21496 26022 21548
rect 26970 21496 26976 21548
rect 27028 21496 27034 21548
rect 27240 21539 27298 21545
rect 27240 21505 27252 21539
rect 27286 21536 27298 21539
rect 27522 21536 27528 21548
rect 27286 21508 27528 21536
rect 27286 21505 27298 21508
rect 27240 21499 27298 21505
rect 27522 21496 27528 21508
rect 27580 21496 27586 21548
rect 27632 21536 27660 21644
rect 28350 21632 28356 21684
rect 28408 21632 28414 21684
rect 29825 21675 29883 21681
rect 29825 21641 29837 21675
rect 29871 21672 29883 21675
rect 30926 21672 30932 21684
rect 29871 21644 30932 21672
rect 29871 21641 29883 21644
rect 29825 21635 29883 21641
rect 30926 21632 30932 21644
rect 30984 21632 30990 21684
rect 32398 21632 32404 21684
rect 32456 21632 32462 21684
rect 35066 21672 35072 21684
rect 32508 21644 34284 21672
rect 28712 21607 28770 21613
rect 28712 21573 28724 21607
rect 28758 21604 28770 21607
rect 29546 21604 29552 21616
rect 28758 21576 29552 21604
rect 28758 21573 28770 21576
rect 28712 21567 28770 21573
rect 29546 21564 29552 21576
rect 29604 21564 29610 21616
rect 31478 21564 31484 21616
rect 31536 21604 31542 21616
rect 32508 21604 32536 21644
rect 32784 21613 32812 21644
rect 31536 21576 32536 21604
rect 32769 21607 32827 21613
rect 31536 21564 31542 21576
rect 32769 21573 32781 21607
rect 32815 21573 32827 21607
rect 32769 21567 32827 21573
rect 33042 21564 33048 21616
rect 33100 21604 33106 21616
rect 34256 21613 34284 21644
rect 34716 21644 35072 21672
rect 34716 21613 34744 21644
rect 35066 21632 35072 21644
rect 35124 21672 35130 21684
rect 36446 21672 36452 21684
rect 35124 21644 36452 21672
rect 35124 21632 35130 21644
rect 36446 21632 36452 21644
rect 36504 21632 36510 21684
rect 41322 21632 41328 21684
rect 41380 21632 41386 21684
rect 34149 21607 34207 21613
rect 34149 21604 34161 21607
rect 33100 21576 34161 21604
rect 33100 21564 33106 21576
rect 34149 21573 34161 21576
rect 34195 21573 34207 21607
rect 34149 21567 34207 21573
rect 34241 21607 34299 21613
rect 34241 21573 34253 21607
rect 34287 21604 34299 21607
rect 34701 21607 34759 21613
rect 34701 21604 34713 21607
rect 34287 21576 34713 21604
rect 34287 21573 34299 21576
rect 34241 21567 34299 21573
rect 34701 21573 34713 21576
rect 34747 21573 34759 21607
rect 34701 21567 34759 21573
rect 34793 21607 34851 21613
rect 34793 21573 34805 21607
rect 34839 21604 34851 21607
rect 35342 21604 35348 21616
rect 34839 21576 35348 21604
rect 34839 21573 34851 21576
rect 34793 21567 34851 21573
rect 35342 21564 35348 21576
rect 35400 21564 35406 21616
rect 40402 21604 40408 21616
rect 39960 21576 40408 21604
rect 32490 21536 32496 21548
rect 27632 21508 32496 21536
rect 32490 21496 32496 21508
rect 32548 21496 32554 21548
rect 32585 21539 32643 21545
rect 32585 21505 32597 21539
rect 32631 21505 32643 21539
rect 32585 21499 32643 21505
rect 32677 21539 32735 21545
rect 32677 21505 32689 21539
rect 32723 21505 32735 21539
rect 32677 21499 32735 21505
rect 32953 21539 33011 21545
rect 32953 21505 32965 21539
rect 32999 21536 33011 21539
rect 33410 21536 33416 21548
rect 32999 21508 33416 21536
rect 32999 21505 33011 21508
rect 32953 21499 33011 21505
rect 22649 21471 22707 21477
rect 22649 21468 22661 21471
rect 22480 21440 22661 21468
rect 22373 21431 22431 21437
rect 22649 21437 22661 21440
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 20257 21403 20315 21409
rect 20257 21369 20269 21403
rect 20303 21369 20315 21403
rect 20257 21363 20315 21369
rect 20622 21360 20628 21412
rect 20680 21400 20686 21412
rect 22388 21400 22416 21431
rect 23198 21428 23204 21480
rect 23256 21428 23262 21480
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21437 23535 21471
rect 25148 21468 25176 21496
rect 25869 21471 25927 21477
rect 25869 21468 25881 21471
rect 25148 21440 25881 21468
rect 23477 21431 23535 21437
rect 25869 21437 25881 21440
rect 25915 21437 25927 21471
rect 25869 21431 25927 21437
rect 26513 21471 26571 21477
rect 26513 21437 26525 21471
rect 26559 21468 26571 21471
rect 26602 21468 26608 21480
rect 26559 21440 26608 21468
rect 26559 21437 26571 21440
rect 26513 21431 26571 21437
rect 20680 21372 22416 21400
rect 20680 21360 20686 21372
rect 18012 21304 20208 21332
rect 20349 21335 20407 21341
rect 18012 21292 18018 21304
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20438 21332 20444 21344
rect 20395 21304 20444 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21818 21292 21824 21344
rect 21876 21292 21882 21344
rect 22388 21332 22416 21372
rect 22462 21360 22468 21412
rect 22520 21400 22526 21412
rect 23492 21400 23520 21431
rect 26602 21428 26608 21440
rect 26660 21428 26666 21480
rect 28442 21428 28448 21480
rect 28500 21428 28506 21480
rect 30098 21428 30104 21480
rect 30156 21468 30162 21480
rect 30653 21471 30711 21477
rect 30653 21468 30665 21471
rect 30156 21440 30665 21468
rect 30156 21428 30162 21440
rect 30653 21437 30665 21440
rect 30699 21437 30711 21471
rect 30653 21431 30711 21437
rect 31846 21428 31852 21480
rect 31904 21428 31910 21480
rect 32600 21468 32628 21499
rect 32508 21440 32628 21468
rect 22520 21372 23520 21400
rect 22520 21360 22526 21372
rect 23750 21332 23756 21344
rect 22388 21304 23756 21332
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 25958 21292 25964 21344
rect 26016 21332 26022 21344
rect 28810 21332 28816 21344
rect 26016 21304 28816 21332
rect 26016 21292 26022 21304
rect 28810 21292 28816 21304
rect 28868 21292 28874 21344
rect 29914 21292 29920 21344
rect 29972 21332 29978 21344
rect 30101 21335 30159 21341
rect 30101 21332 30113 21335
rect 29972 21304 30113 21332
rect 29972 21292 29978 21304
rect 30101 21301 30113 21304
rect 30147 21301 30159 21335
rect 30101 21295 30159 21301
rect 31202 21292 31208 21344
rect 31260 21292 31266 21344
rect 32508 21332 32536 21440
rect 32582 21360 32588 21412
rect 32640 21400 32646 21412
rect 32692 21400 32720 21499
rect 33410 21496 33416 21508
rect 33468 21496 33474 21548
rect 34054 21496 34060 21548
rect 34112 21496 34118 21548
rect 34425 21539 34483 21545
rect 34425 21505 34437 21539
rect 34471 21505 34483 21539
rect 34425 21499 34483 21505
rect 34517 21539 34575 21545
rect 34517 21505 34529 21539
rect 34563 21505 34575 21539
rect 34517 21499 34575 21505
rect 33229 21471 33287 21477
rect 33229 21437 33241 21471
rect 33275 21468 33287 21471
rect 33686 21468 33692 21480
rect 33275 21440 33692 21468
rect 33275 21437 33287 21440
rect 33229 21431 33287 21437
rect 33686 21428 33692 21440
rect 33744 21428 33750 21480
rect 34440 21468 34468 21499
rect 33796 21440 34468 21468
rect 34532 21468 34560 21499
rect 34606 21496 34612 21548
rect 34664 21536 34670 21548
rect 39960 21545 39988 21576
rect 40402 21564 40408 21576
rect 40460 21564 40466 21616
rect 34885 21539 34943 21545
rect 34885 21536 34897 21539
rect 34664 21508 34897 21536
rect 34664 21496 34670 21508
rect 34885 21505 34897 21508
rect 34931 21505 34943 21539
rect 34885 21499 34943 21505
rect 37921 21539 37979 21545
rect 37921 21505 37933 21539
rect 37967 21536 37979 21539
rect 39945 21539 40003 21545
rect 39945 21536 39957 21539
rect 37967 21508 39957 21536
rect 37967 21505 37979 21508
rect 37921 21499 37979 21505
rect 39945 21505 39957 21508
rect 39991 21505 40003 21539
rect 39945 21499 40003 21505
rect 40212 21539 40270 21545
rect 40212 21505 40224 21539
rect 40258 21536 40270 21539
rect 40678 21536 40684 21548
rect 40258 21508 40684 21536
rect 40258 21505 40270 21508
rect 40212 21499 40270 21505
rect 40678 21496 40684 21508
rect 40736 21496 40742 21548
rect 34532 21440 35020 21468
rect 32640 21372 32720 21400
rect 32640 21360 32646 21372
rect 33796 21344 33824 21440
rect 34992 21400 35020 21440
rect 35618 21428 35624 21480
rect 35676 21428 35682 21480
rect 41969 21471 42027 21477
rect 41969 21468 41981 21471
rect 41386 21440 41981 21468
rect 41386 21400 41414 21440
rect 41969 21437 41981 21440
rect 42015 21437 42027 21471
rect 41969 21431 42027 21437
rect 34992 21372 36308 21400
rect 33134 21332 33140 21344
rect 32508 21304 33140 21332
rect 33134 21292 33140 21304
rect 33192 21292 33198 21344
rect 33778 21292 33784 21344
rect 33836 21292 33842 21344
rect 33870 21292 33876 21344
rect 33928 21292 33934 21344
rect 35069 21335 35127 21341
rect 35069 21301 35081 21335
rect 35115 21332 35127 21335
rect 35986 21332 35992 21344
rect 35115 21304 35992 21332
rect 35115 21301 35127 21304
rect 35069 21295 35127 21301
rect 35986 21292 35992 21304
rect 36044 21292 36050 21344
rect 36280 21341 36308 21372
rect 40880 21372 41414 21400
rect 36265 21335 36323 21341
rect 36265 21301 36277 21335
rect 36311 21332 36323 21335
rect 36722 21332 36728 21344
rect 36311 21304 36728 21332
rect 36311 21301 36323 21304
rect 36265 21295 36323 21301
rect 36722 21292 36728 21304
rect 36780 21292 36786 21344
rect 40218 21292 40224 21344
rect 40276 21332 40282 21344
rect 40880 21332 40908 21372
rect 40276 21304 40908 21332
rect 40276 21292 40282 21304
rect 40954 21292 40960 21344
rect 41012 21332 41018 21344
rect 41417 21335 41475 21341
rect 41417 21332 41429 21335
rect 41012 21304 41429 21332
rect 41012 21292 41018 21304
rect 41417 21301 41429 21304
rect 41463 21301 41475 21335
rect 41417 21295 41475 21301
rect 1104 21242 42504 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 42504 21242
rect 1104 21168 42504 21190
rect 5169 21131 5227 21137
rect 5169 21097 5181 21131
rect 5215 21128 5227 21131
rect 5626 21128 5632 21140
rect 5215 21100 5632 21128
rect 5215 21097 5227 21100
rect 5169 21091 5227 21097
rect 5626 21088 5632 21100
rect 5684 21088 5690 21140
rect 6089 21131 6147 21137
rect 6089 21097 6101 21131
rect 6135 21128 6147 21131
rect 6730 21128 6736 21140
rect 6135 21100 6736 21128
rect 6135 21097 6147 21100
rect 6089 21091 6147 21097
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 8113 21131 8171 21137
rect 8113 21097 8125 21131
rect 8159 21128 8171 21131
rect 8846 21128 8852 21140
rect 8159 21100 8852 21128
rect 8159 21097 8171 21100
rect 8113 21091 8171 21097
rect 8846 21088 8852 21100
rect 8904 21088 8910 21140
rect 15473 21131 15531 21137
rect 15473 21097 15485 21131
rect 15519 21128 15531 21131
rect 16114 21128 16120 21140
rect 15519 21100 16120 21128
rect 15519 21097 15531 21100
rect 15473 21091 15531 21097
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 17497 21131 17555 21137
rect 17497 21097 17509 21131
rect 17543 21128 17555 21131
rect 17543 21100 18460 21128
rect 17543 21097 17555 21100
rect 17497 21091 17555 21097
rect 3145 21063 3203 21069
rect 3145 21029 3157 21063
rect 3191 21060 3203 21063
rect 4525 21063 4583 21069
rect 3191 21032 4016 21060
rect 3191 21029 3203 21032
rect 3145 21023 3203 21029
rect 3988 20936 4016 21032
rect 4525 21029 4537 21063
rect 4571 21060 4583 21063
rect 4614 21060 4620 21072
rect 4571 21032 4620 21060
rect 4571 21029 4583 21032
rect 4525 21023 4583 21029
rect 4614 21020 4620 21032
rect 4672 21020 4678 21072
rect 10873 21063 10931 21069
rect 10873 21029 10885 21063
rect 10919 21029 10931 21063
rect 10873 21023 10931 21029
rect 5258 20992 5264 21004
rect 5000 20964 5264 20992
rect 1670 20884 1676 20936
rect 1728 20924 1734 20936
rect 1765 20927 1823 20933
rect 1765 20924 1777 20927
rect 1728 20896 1777 20924
rect 1728 20884 1734 20896
rect 1765 20893 1777 20896
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 2032 20927 2090 20933
rect 2032 20893 2044 20927
rect 2078 20924 2090 20927
rect 2590 20924 2596 20936
rect 2078 20896 2596 20924
rect 2078 20893 2090 20896
rect 2032 20887 2090 20893
rect 2590 20884 2596 20896
rect 2648 20884 2654 20936
rect 3050 20884 3056 20936
rect 3108 20924 3114 20936
rect 3237 20927 3295 20933
rect 3237 20924 3249 20927
rect 3108 20896 3249 20924
rect 3108 20884 3114 20896
rect 3237 20893 3249 20896
rect 3283 20893 3295 20927
rect 3237 20887 3295 20893
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20893 3479 20927
rect 3421 20887 3479 20893
rect 3436 20856 3464 20887
rect 3970 20884 3976 20936
rect 4028 20924 4034 20936
rect 4341 20927 4399 20933
rect 4341 20924 4353 20927
rect 4028 20896 4353 20924
rect 4028 20884 4034 20896
rect 4341 20893 4353 20896
rect 4387 20893 4399 20927
rect 4341 20887 4399 20893
rect 4798 20884 4804 20936
rect 4856 20884 4862 20936
rect 5000 20933 5028 20964
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 6365 20995 6423 21001
rect 6365 20961 6377 20995
rect 6411 20992 6423 20995
rect 6638 20992 6644 21004
rect 6411 20964 6644 20992
rect 6411 20961 6423 20964
rect 6365 20955 6423 20961
rect 6638 20952 6644 20964
rect 6696 20952 6702 21004
rect 10778 20952 10784 21004
rect 10836 20992 10842 21004
rect 10888 20992 10916 21023
rect 11517 20995 11575 21001
rect 11517 20992 11529 20995
rect 10836 20964 11529 20992
rect 10836 20952 10842 20964
rect 11517 20961 11529 20964
rect 11563 20961 11575 20995
rect 11517 20955 11575 20961
rect 11790 20952 11796 21004
rect 11848 20952 11854 21004
rect 16022 20952 16028 21004
rect 16080 20952 16086 21004
rect 16209 20995 16267 21001
rect 16209 20961 16221 20995
rect 16255 20992 16267 20995
rect 17402 20992 17408 21004
rect 16255 20964 17408 20992
rect 16255 20961 16267 20964
rect 16209 20955 16267 20961
rect 17402 20952 17408 20964
rect 17460 20992 17466 21004
rect 17512 20992 17540 21091
rect 18325 21063 18383 21069
rect 18325 21029 18337 21063
rect 18371 21029 18383 21063
rect 18432 21060 18460 21100
rect 19150 21088 19156 21140
rect 19208 21128 19214 21140
rect 19245 21131 19303 21137
rect 19245 21128 19257 21131
rect 19208 21100 19257 21128
rect 19208 21088 19214 21100
rect 19245 21097 19257 21100
rect 19291 21097 19303 21131
rect 19245 21091 19303 21097
rect 22281 21131 22339 21137
rect 22281 21097 22293 21131
rect 22327 21128 22339 21131
rect 23198 21128 23204 21140
rect 22327 21100 23204 21128
rect 22327 21097 22339 21100
rect 22281 21091 22339 21097
rect 23198 21088 23204 21100
rect 23256 21088 23262 21140
rect 28997 21131 29055 21137
rect 28997 21097 29009 21131
rect 29043 21128 29055 21131
rect 29086 21128 29092 21140
rect 29043 21100 29092 21128
rect 29043 21097 29055 21100
rect 28997 21091 29055 21097
rect 29086 21088 29092 21100
rect 29144 21088 29150 21140
rect 38654 21088 38660 21140
rect 38712 21088 38718 21140
rect 20622 21060 20628 21072
rect 18432 21032 20628 21060
rect 18325 21023 18383 21029
rect 17460 20964 17540 20992
rect 18340 20992 18368 21023
rect 20622 21020 20628 21032
rect 20680 21020 20686 21072
rect 27617 21063 27675 21069
rect 27617 21029 27629 21063
rect 27663 21060 27675 21063
rect 27890 21060 27896 21072
rect 27663 21032 27896 21060
rect 27663 21029 27675 21032
rect 27617 21023 27675 21029
rect 27890 21020 27896 21032
rect 27948 21060 27954 21072
rect 27948 21032 28304 21060
rect 27948 21020 27954 21032
rect 18417 20995 18475 21001
rect 18417 20992 18429 20995
rect 18340 20964 18429 20992
rect 17460 20952 17466 20964
rect 18417 20961 18429 20964
rect 18463 20961 18475 20995
rect 18417 20955 18475 20961
rect 24762 20952 24768 21004
rect 24820 20992 24826 21004
rect 24857 20995 24915 21001
rect 24857 20992 24869 20995
rect 24820 20964 24869 20992
rect 24820 20952 24826 20964
rect 24857 20961 24869 20964
rect 24903 20961 24915 20995
rect 24857 20955 24915 20961
rect 24946 20952 24952 21004
rect 25004 20952 25010 21004
rect 28276 21001 28304 21032
rect 28442 21020 28448 21072
rect 28500 21060 28506 21072
rect 28500 21032 30512 21060
rect 28500 21020 28506 21032
rect 28261 20995 28319 21001
rect 28261 20961 28273 20995
rect 28307 20961 28319 20995
rect 28261 20955 28319 20961
rect 29822 20952 29828 21004
rect 29880 20992 29886 21004
rect 30484 21001 30512 21032
rect 30009 20995 30067 21001
rect 30009 20992 30021 20995
rect 29880 20964 30021 20992
rect 29880 20952 29886 20964
rect 30009 20961 30021 20964
rect 30055 20961 30067 20995
rect 30009 20955 30067 20961
rect 30193 20995 30251 21001
rect 30193 20961 30205 20995
rect 30239 20961 30251 20995
rect 30193 20955 30251 20961
rect 30469 20995 30527 21001
rect 30469 20961 30481 20995
rect 30515 20961 30527 20995
rect 30469 20955 30527 20961
rect 4985 20927 5043 20933
rect 4985 20893 4997 20927
rect 5031 20893 5043 20927
rect 4985 20887 5043 20893
rect 5169 20927 5227 20933
rect 5169 20893 5181 20927
rect 5215 20924 5227 20927
rect 5350 20924 5356 20936
rect 5215 20896 5356 20924
rect 5215 20893 5227 20896
rect 5169 20887 5227 20893
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20893 6055 20927
rect 5997 20887 6055 20893
rect 4154 20856 4160 20868
rect 3436 20828 4160 20856
rect 4154 20816 4160 20828
rect 4212 20816 4218 20868
rect 4522 20816 4528 20868
rect 4580 20816 4586 20868
rect 6012 20856 6040 20887
rect 6178 20884 6184 20936
rect 6236 20884 6242 20936
rect 8386 20884 8392 20936
rect 8444 20924 8450 20936
rect 8665 20927 8723 20933
rect 8665 20924 8677 20927
rect 8444 20896 8677 20924
rect 8444 20884 8450 20896
rect 8665 20893 8677 20896
rect 8711 20924 8723 20927
rect 9493 20927 9551 20933
rect 9493 20924 9505 20927
rect 8711 20896 9505 20924
rect 8711 20893 8723 20896
rect 8665 20887 8723 20893
rect 9493 20893 9505 20896
rect 9539 20924 9551 20927
rect 10134 20924 10140 20936
rect 9539 20896 10140 20924
rect 9539 20893 9551 20896
rect 9493 20887 9551 20893
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20924 11943 20927
rect 12529 20927 12587 20933
rect 12529 20924 12541 20927
rect 11931 20896 12541 20924
rect 11931 20893 11943 20896
rect 11885 20887 11943 20893
rect 12529 20893 12541 20896
rect 12575 20893 12587 20927
rect 12529 20887 12587 20893
rect 13170 20884 13176 20936
rect 13228 20884 13234 20936
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20924 14151 20927
rect 14139 20896 14504 20924
rect 14139 20893 14151 20896
rect 14093 20887 14151 20893
rect 14476 20868 14504 20896
rect 16574 20884 16580 20936
rect 16632 20924 16638 20936
rect 16945 20927 17003 20933
rect 16945 20924 16957 20927
rect 16632 20896 16957 20924
rect 16632 20884 16638 20896
rect 16945 20893 16957 20896
rect 16991 20893 17003 20927
rect 16945 20887 17003 20893
rect 17218 20884 17224 20936
rect 17276 20884 17282 20936
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20893 17831 20927
rect 17773 20887 17831 20893
rect 6362 20856 6368 20868
rect 6012 20828 6368 20856
rect 6362 20816 6368 20828
rect 6420 20816 6426 20868
rect 6641 20859 6699 20865
rect 6641 20825 6653 20859
rect 6687 20856 6699 20859
rect 6914 20856 6920 20868
rect 6687 20828 6920 20856
rect 6687 20825 6699 20828
rect 6641 20819 6699 20825
rect 6914 20816 6920 20828
rect 6972 20816 6978 20868
rect 9766 20865 9772 20868
rect 7024 20828 7130 20856
rect 7024 20800 7052 20828
rect 9760 20819 9772 20865
rect 9766 20816 9772 20819
rect 9824 20816 9830 20868
rect 14366 20865 14372 20868
rect 14360 20856 14372 20865
rect 14327 20828 14372 20856
rect 14360 20819 14372 20828
rect 14366 20816 14372 20819
rect 14424 20816 14430 20868
rect 14458 20816 14464 20868
rect 14516 20816 14522 20868
rect 15933 20859 15991 20865
rect 15933 20825 15945 20859
rect 15979 20856 15991 20859
rect 16393 20859 16451 20865
rect 16393 20856 16405 20859
rect 15979 20828 16405 20856
rect 15979 20825 15991 20828
rect 15933 20819 15991 20825
rect 16393 20825 16405 20828
rect 16439 20825 16451 20859
rect 16393 20819 16451 20825
rect 3326 20748 3332 20800
rect 3384 20748 3390 20800
rect 3418 20748 3424 20800
rect 3476 20788 3482 20800
rect 3789 20791 3847 20797
rect 3789 20788 3801 20791
rect 3476 20760 3801 20788
rect 3476 20748 3482 20760
rect 3789 20757 3801 20760
rect 3835 20757 3847 20791
rect 3789 20751 3847 20757
rect 4706 20748 4712 20800
rect 4764 20748 4770 20800
rect 7006 20748 7012 20800
rect 7064 20748 7070 20800
rect 10962 20748 10968 20800
rect 11020 20748 11026 20800
rect 12250 20748 12256 20800
rect 12308 20748 12314 20800
rect 15562 20748 15568 20800
rect 15620 20748 15626 20800
rect 17788 20788 17816 20887
rect 17954 20884 17960 20936
rect 18012 20884 18018 20936
rect 18138 20884 18144 20936
rect 18196 20884 18202 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19392 20896 19809 20924
rect 19392 20884 19398 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 20070 20884 20076 20936
rect 20128 20924 20134 20936
rect 20533 20927 20591 20933
rect 20533 20924 20545 20927
rect 20128 20896 20545 20924
rect 20128 20884 20134 20896
rect 20533 20893 20545 20896
rect 20579 20893 20591 20927
rect 20533 20887 20591 20893
rect 20901 20927 20959 20933
rect 20901 20893 20913 20927
rect 20947 20924 20959 20927
rect 21450 20924 21456 20936
rect 20947 20896 21456 20924
rect 20947 20893 20959 20896
rect 20901 20887 20959 20893
rect 21450 20884 21456 20896
rect 21508 20924 21514 20936
rect 22462 20924 22468 20936
rect 21508 20896 22468 20924
rect 21508 20884 21514 20896
rect 22462 20884 22468 20896
rect 22520 20884 22526 20936
rect 25774 20884 25780 20936
rect 25832 20884 25838 20936
rect 26237 20927 26295 20933
rect 26237 20893 26249 20927
rect 26283 20924 26295 20927
rect 26970 20924 26976 20936
rect 26283 20896 26976 20924
rect 26283 20893 26295 20896
rect 26237 20887 26295 20893
rect 26970 20884 26976 20896
rect 27028 20884 27034 20936
rect 28445 20927 28503 20933
rect 28445 20893 28457 20927
rect 28491 20924 28503 20927
rect 28534 20924 28540 20936
rect 28491 20896 28540 20924
rect 28491 20893 28503 20896
rect 28445 20887 28503 20893
rect 28534 20884 28540 20896
rect 28592 20884 28598 20936
rect 28718 20884 28724 20936
rect 28776 20884 28782 20936
rect 28810 20884 28816 20936
rect 28868 20884 28874 20936
rect 29914 20884 29920 20936
rect 29972 20884 29978 20936
rect 18049 20859 18107 20865
rect 18049 20825 18061 20859
rect 18095 20856 18107 20859
rect 18230 20856 18236 20868
rect 18095 20828 18236 20856
rect 18095 20825 18107 20828
rect 18049 20819 18107 20825
rect 18230 20816 18236 20828
rect 18288 20816 18294 20868
rect 19981 20859 20039 20865
rect 19981 20856 19993 20859
rect 18340 20828 19993 20856
rect 18340 20788 18368 20828
rect 19981 20825 19993 20828
rect 20027 20825 20039 20859
rect 19981 20819 20039 20825
rect 21168 20859 21226 20865
rect 21168 20825 21180 20859
rect 21214 20856 21226 20859
rect 21818 20856 21824 20868
rect 21214 20828 21824 20856
rect 21214 20825 21226 20828
rect 21168 20819 21226 20825
rect 21818 20816 21824 20828
rect 21876 20816 21882 20868
rect 24765 20859 24823 20865
rect 24765 20825 24777 20859
rect 24811 20856 24823 20859
rect 25225 20859 25283 20865
rect 25225 20856 25237 20859
rect 24811 20828 25237 20856
rect 24811 20825 24823 20828
rect 24765 20819 24823 20825
rect 25225 20825 25237 20828
rect 25271 20825 25283 20859
rect 25225 20819 25283 20825
rect 26326 20816 26332 20868
rect 26384 20856 26390 20868
rect 26482 20859 26540 20865
rect 26482 20856 26494 20859
rect 26384 20828 26494 20856
rect 26384 20816 26390 20828
rect 26482 20825 26494 20828
rect 26528 20825 26540 20859
rect 28629 20859 28687 20865
rect 28629 20856 28641 20859
rect 26482 20819 26540 20825
rect 26620 20828 28641 20856
rect 17788 20760 18368 20788
rect 19058 20748 19064 20800
rect 19116 20748 19122 20800
rect 23474 20748 23480 20800
rect 23532 20788 23538 20800
rect 24397 20791 24455 20797
rect 24397 20788 24409 20791
rect 23532 20760 24409 20788
rect 23532 20748 23538 20760
rect 24397 20757 24409 20760
rect 24443 20757 24455 20791
rect 24397 20751 24455 20757
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 25866 20788 25872 20800
rect 25372 20760 25872 20788
rect 25372 20748 25378 20760
rect 25866 20748 25872 20760
rect 25924 20788 25930 20800
rect 26620 20788 26648 20828
rect 28629 20825 28641 20828
rect 28675 20856 28687 20859
rect 30208 20856 30236 20955
rect 39206 20952 39212 21004
rect 39264 20952 39270 21004
rect 39390 20952 39396 21004
rect 39448 20952 39454 21004
rect 40034 20952 40040 21004
rect 40092 20992 40098 21004
rect 40402 20992 40408 21004
rect 40092 20964 40408 20992
rect 40092 20952 40098 20964
rect 40402 20952 40408 20964
rect 40460 20952 40466 21004
rect 30736 20927 30794 20933
rect 30736 20893 30748 20927
rect 30782 20924 30794 20927
rect 31110 20924 31116 20936
rect 30782 20896 31116 20924
rect 30782 20893 30794 20896
rect 30736 20887 30794 20893
rect 31110 20884 31116 20896
rect 31168 20884 31174 20936
rect 31754 20884 31760 20936
rect 31812 20924 31818 20936
rect 32122 20924 32128 20936
rect 31812 20896 32128 20924
rect 31812 20884 31818 20896
rect 32122 20884 32128 20896
rect 32180 20924 32186 20936
rect 32217 20927 32275 20933
rect 32217 20924 32229 20927
rect 32180 20896 32229 20924
rect 32180 20884 32186 20896
rect 32217 20893 32229 20896
rect 32263 20893 32275 20927
rect 32217 20887 32275 20893
rect 32484 20927 32542 20933
rect 32484 20893 32496 20927
rect 32530 20924 32542 20927
rect 33870 20924 33876 20936
rect 32530 20896 33876 20924
rect 32530 20893 32542 20896
rect 32484 20887 32542 20893
rect 33870 20884 33876 20896
rect 33928 20884 33934 20936
rect 35986 20884 35992 20936
rect 36044 20924 36050 20936
rect 36274 20927 36332 20933
rect 36274 20924 36286 20927
rect 36044 20896 36286 20924
rect 36044 20884 36050 20896
rect 36274 20893 36286 20896
rect 36320 20893 36332 20927
rect 36274 20887 36332 20893
rect 36538 20884 36544 20936
rect 36596 20924 36602 20936
rect 37182 20924 37188 20936
rect 36596 20896 37188 20924
rect 36596 20884 36602 20896
rect 37182 20884 37188 20896
rect 37240 20924 37246 20936
rect 37550 20933 37556 20936
rect 37277 20927 37335 20933
rect 37277 20924 37289 20927
rect 37240 20896 37289 20924
rect 37240 20884 37246 20896
rect 37277 20893 37289 20896
rect 37323 20893 37335 20927
rect 37277 20887 37335 20893
rect 37544 20887 37556 20933
rect 37550 20884 37556 20887
rect 37608 20884 37614 20936
rect 39408 20924 39436 20952
rect 39408 20896 40448 20924
rect 40420 20868 40448 20896
rect 34330 20856 34336 20868
rect 28675 20828 29684 20856
rect 30208 20828 34336 20856
rect 28675 20825 28687 20828
rect 28629 20819 28687 20825
rect 25924 20760 26648 20788
rect 25924 20748 25930 20760
rect 27614 20748 27620 20800
rect 27672 20788 27678 20800
rect 27709 20791 27767 20797
rect 27709 20788 27721 20791
rect 27672 20760 27721 20788
rect 27672 20748 27678 20760
rect 27709 20757 27721 20760
rect 27755 20757 27767 20791
rect 27709 20751 27767 20757
rect 29086 20748 29092 20800
rect 29144 20788 29150 20800
rect 29549 20791 29607 20797
rect 29549 20788 29561 20791
rect 29144 20760 29561 20788
rect 29144 20748 29150 20760
rect 29549 20757 29561 20760
rect 29595 20757 29607 20791
rect 29656 20788 29684 20828
rect 34330 20816 34336 20828
rect 34388 20816 34394 20868
rect 40402 20816 40408 20868
rect 40460 20816 40466 20868
rect 40678 20816 40684 20868
rect 40736 20816 40742 20868
rect 41230 20816 41236 20868
rect 41288 20816 41294 20868
rect 31478 20788 31484 20800
rect 29656 20760 31484 20788
rect 29549 20751 29607 20757
rect 31478 20748 31484 20760
rect 31536 20748 31542 20800
rect 31846 20748 31852 20800
rect 31904 20788 31910 20800
rect 32306 20788 32312 20800
rect 31904 20760 32312 20788
rect 31904 20748 31910 20760
rect 32306 20748 32312 20760
rect 32364 20748 32370 20800
rect 32490 20748 32496 20800
rect 32548 20788 32554 20800
rect 32766 20788 32772 20800
rect 32548 20760 32772 20788
rect 32548 20748 32554 20760
rect 32766 20748 32772 20760
rect 32824 20748 32830 20800
rect 33597 20791 33655 20797
rect 33597 20757 33609 20791
rect 33643 20788 33655 20791
rect 33686 20788 33692 20800
rect 33643 20760 33692 20788
rect 33643 20757 33655 20760
rect 33597 20751 33655 20757
rect 33686 20748 33692 20760
rect 33744 20748 33750 20800
rect 34606 20748 34612 20800
rect 34664 20788 34670 20800
rect 35161 20791 35219 20797
rect 35161 20788 35173 20791
rect 34664 20760 35173 20788
rect 34664 20748 34670 20760
rect 35161 20757 35173 20760
rect 35207 20788 35219 20791
rect 35618 20788 35624 20800
rect 35207 20760 35624 20788
rect 35207 20757 35219 20760
rect 35161 20751 35219 20757
rect 35618 20748 35624 20760
rect 35676 20748 35682 20800
rect 38746 20748 38752 20800
rect 38804 20748 38810 20800
rect 39117 20791 39175 20797
rect 39117 20757 39129 20791
rect 39163 20788 39175 20791
rect 39574 20788 39580 20800
rect 39163 20760 39580 20788
rect 39163 20757 39175 20760
rect 39117 20751 39175 20757
rect 39574 20748 39580 20760
rect 39632 20748 39638 20800
rect 42150 20748 42156 20800
rect 42208 20748 42214 20800
rect 1104 20698 42504 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 42504 20698
rect 1104 20624 42504 20646
rect 3053 20587 3111 20593
rect 3053 20553 3065 20587
rect 3099 20584 3111 20587
rect 3142 20584 3148 20596
rect 3099 20556 3148 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 4522 20544 4528 20596
rect 4580 20544 4586 20596
rect 6270 20544 6276 20596
rect 6328 20584 6334 20596
rect 6365 20587 6423 20593
rect 6365 20584 6377 20587
rect 6328 20556 6377 20584
rect 6328 20544 6334 20556
rect 6365 20553 6377 20556
rect 6411 20553 6423 20587
rect 6365 20547 6423 20553
rect 9766 20544 9772 20596
rect 9824 20544 9830 20596
rect 13170 20544 13176 20596
rect 13228 20584 13234 20596
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 13228 20556 13277 20584
rect 13228 20544 13234 20556
rect 13265 20553 13277 20556
rect 13311 20553 13323 20587
rect 13265 20547 13323 20553
rect 18417 20587 18475 20593
rect 18417 20553 18429 20587
rect 18463 20584 18475 20587
rect 18598 20584 18604 20596
rect 18463 20556 18604 20584
rect 18463 20553 18475 20556
rect 18417 20547 18475 20553
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 22278 20544 22284 20596
rect 22336 20544 22342 20596
rect 24857 20587 24915 20593
rect 24857 20553 24869 20587
rect 24903 20584 24915 20587
rect 25774 20584 25780 20596
rect 24903 20556 25780 20584
rect 24903 20553 24915 20556
rect 24857 20547 24915 20553
rect 25774 20544 25780 20556
rect 25832 20544 25838 20596
rect 26145 20587 26203 20593
rect 26145 20553 26157 20587
rect 26191 20584 26203 20587
rect 26326 20584 26332 20596
rect 26191 20556 26332 20584
rect 26191 20553 26203 20556
rect 26145 20547 26203 20553
rect 26326 20544 26332 20556
rect 26384 20544 26390 20596
rect 27706 20544 27712 20596
rect 27764 20584 27770 20596
rect 27801 20587 27859 20593
rect 27801 20584 27813 20587
rect 27764 20556 27813 20584
rect 27764 20544 27770 20556
rect 27801 20553 27813 20556
rect 27847 20553 27859 20587
rect 27801 20547 27859 20553
rect 28994 20544 29000 20596
rect 29052 20584 29058 20596
rect 32398 20584 32404 20596
rect 29052 20556 32404 20584
rect 29052 20544 29058 20556
rect 32398 20544 32404 20556
rect 32456 20544 32462 20596
rect 32692 20556 34836 20584
rect 8386 20476 8392 20528
rect 8444 20476 8450 20528
rect 12152 20519 12210 20525
rect 12152 20485 12164 20519
rect 12198 20516 12210 20519
rect 12250 20516 12256 20528
rect 12198 20488 12256 20516
rect 12198 20485 12210 20488
rect 12152 20479 12210 20485
rect 12250 20476 12256 20488
rect 12308 20476 12314 20528
rect 14728 20519 14786 20525
rect 14728 20485 14740 20519
rect 14774 20516 14786 20519
rect 15562 20516 15568 20528
rect 14774 20488 15568 20516
rect 14774 20485 14786 20488
rect 14728 20479 14786 20485
rect 15562 20476 15568 20488
rect 15620 20476 15626 20528
rect 18960 20519 19018 20525
rect 18960 20485 18972 20519
rect 19006 20516 19018 20519
rect 19058 20516 19064 20528
rect 19006 20488 19064 20516
rect 19006 20485 19018 20488
rect 18960 20479 19018 20485
rect 19058 20476 19064 20488
rect 19116 20476 19122 20528
rect 23385 20519 23443 20525
rect 23385 20485 23397 20519
rect 23431 20516 23443 20519
rect 23474 20516 23480 20528
rect 23431 20488 23480 20516
rect 23431 20485 23443 20488
rect 23385 20479 23443 20485
rect 23474 20476 23480 20488
rect 23532 20476 23538 20528
rect 25498 20516 25504 20528
rect 24610 20488 25504 20516
rect 25498 20476 25504 20488
rect 25556 20476 25562 20528
rect 25869 20519 25927 20525
rect 25869 20485 25881 20519
rect 25915 20516 25927 20519
rect 26050 20516 26056 20528
rect 25915 20488 26056 20516
rect 25915 20485 25927 20488
rect 25869 20479 25927 20485
rect 26050 20476 26056 20488
rect 26108 20476 26114 20528
rect 29178 20476 29184 20528
rect 29236 20476 29242 20528
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20448 1639 20451
rect 1670 20448 1676 20460
rect 1627 20420 1676 20448
rect 1627 20417 1639 20420
rect 1581 20411 1639 20417
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 1854 20457 1860 20460
rect 1848 20411 1860 20457
rect 1854 20408 1860 20411
rect 1912 20408 1918 20460
rect 3418 20408 3424 20460
rect 3476 20408 3482 20460
rect 4614 20408 4620 20460
rect 4672 20408 4678 20460
rect 5258 20408 5264 20460
rect 5316 20448 5322 20460
rect 6546 20448 6552 20460
rect 5316 20420 6552 20448
rect 5316 20408 5322 20420
rect 6546 20408 6552 20420
rect 6604 20448 6610 20460
rect 6733 20451 6791 20457
rect 6733 20448 6745 20451
rect 6604 20420 6745 20448
rect 6604 20408 6610 20420
rect 6733 20417 6745 20420
rect 6779 20448 6791 20451
rect 8938 20448 8944 20460
rect 6779 20420 8944 20448
rect 6779 20417 6791 20420
rect 6733 20411 6791 20417
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 9122 20408 9128 20460
rect 9180 20408 9186 20460
rect 9401 20451 9459 20457
rect 9401 20417 9413 20451
rect 9447 20448 9459 20451
rect 10962 20448 10968 20460
rect 9447 20420 10968 20448
rect 9447 20417 9459 20420
rect 9401 20411 9459 20417
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 11606 20408 11612 20460
rect 11664 20448 11670 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11664 20420 11897 20448
rect 11664 20408 11670 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 16666 20408 16672 20460
rect 16724 20408 16730 20460
rect 20714 20448 20720 20460
rect 18078 20420 20720 20448
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 21637 20451 21695 20457
rect 21637 20417 21649 20451
rect 21683 20448 21695 20451
rect 22189 20451 22247 20457
rect 22189 20448 22201 20451
rect 21683 20420 22201 20448
rect 21683 20417 21695 20420
rect 21637 20411 21695 20417
rect 22189 20417 22201 20420
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 25593 20451 25651 20457
rect 25593 20417 25605 20451
rect 25639 20417 25651 20451
rect 25593 20411 25651 20417
rect 25777 20451 25835 20457
rect 25777 20417 25789 20451
rect 25823 20417 25835 20451
rect 25777 20411 25835 20417
rect 3326 20340 3332 20392
rect 3384 20340 3390 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 6270 20340 6276 20392
rect 6328 20380 6334 20392
rect 6641 20383 6699 20389
rect 6641 20380 6653 20383
rect 6328 20352 6653 20380
rect 6328 20340 6334 20352
rect 6641 20349 6653 20352
rect 6687 20349 6699 20383
rect 6641 20343 6699 20349
rect 8478 20340 8484 20392
rect 8536 20380 8542 20392
rect 9309 20383 9367 20389
rect 9309 20380 9321 20383
rect 8536 20352 9321 20380
rect 8536 20340 8542 20352
rect 9309 20349 9321 20352
rect 9355 20349 9367 20383
rect 9309 20343 9367 20349
rect 14458 20340 14464 20392
rect 14516 20340 14522 20392
rect 16209 20383 16267 20389
rect 16209 20380 16221 20383
rect 15856 20352 16221 20380
rect 15856 20321 15884 20352
rect 16209 20349 16221 20352
rect 16255 20380 16267 20383
rect 16574 20380 16580 20392
rect 16255 20352 16580 20380
rect 16255 20349 16267 20352
rect 16209 20343 16267 20349
rect 16574 20340 16580 20352
rect 16632 20340 16638 20392
rect 16945 20383 17003 20389
rect 16945 20349 16957 20383
rect 16991 20380 17003 20383
rect 17310 20380 17316 20392
rect 16991 20352 17316 20380
rect 16991 20349 17003 20352
rect 16945 20343 17003 20349
rect 17310 20340 17316 20352
rect 17368 20340 17374 20392
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18693 20383 18751 20389
rect 18693 20380 18705 20383
rect 18012 20352 18705 20380
rect 18012 20340 18018 20352
rect 18693 20349 18705 20352
rect 18739 20349 18751 20383
rect 18693 20343 18751 20349
rect 21082 20340 21088 20392
rect 21140 20340 21146 20392
rect 22370 20340 22376 20392
rect 22428 20340 22434 20392
rect 22462 20340 22468 20392
rect 22520 20380 22526 20392
rect 23109 20383 23167 20389
rect 23109 20380 23121 20383
rect 22520 20352 23121 20380
rect 22520 20340 22526 20352
rect 23109 20349 23121 20352
rect 23155 20349 23167 20383
rect 23109 20343 23167 20349
rect 15841 20315 15899 20321
rect 15841 20281 15853 20315
rect 15887 20281 15899 20315
rect 25608 20312 25636 20411
rect 25792 20380 25820 20411
rect 25958 20408 25964 20460
rect 26016 20408 26022 20460
rect 28350 20408 28356 20460
rect 28408 20408 28414 20460
rect 32692 20457 32720 20556
rect 34808 20528 34836 20556
rect 40218 20544 40224 20596
rect 40276 20544 40282 20596
rect 40678 20544 40684 20596
rect 40736 20584 40742 20596
rect 41141 20587 41199 20593
rect 41141 20584 41153 20587
rect 40736 20556 41153 20584
rect 40736 20544 40742 20556
rect 41141 20553 41153 20556
rect 41187 20553 41199 20587
rect 41141 20547 41199 20553
rect 41601 20587 41659 20593
rect 41601 20553 41613 20587
rect 41647 20584 41659 20587
rect 41966 20584 41972 20596
rect 41647 20556 41972 20584
rect 41647 20553 41659 20556
rect 41601 20547 41659 20553
rect 41966 20544 41972 20556
rect 42024 20544 42030 20596
rect 32766 20476 32772 20528
rect 32824 20516 32830 20528
rect 32861 20519 32919 20525
rect 32861 20516 32873 20519
rect 32824 20488 32873 20516
rect 32824 20476 32830 20488
rect 32861 20485 32873 20488
rect 32907 20485 32919 20519
rect 32861 20479 32919 20485
rect 32953 20519 33011 20525
rect 32953 20485 32965 20519
rect 32999 20516 33011 20519
rect 33318 20516 33324 20528
rect 32999 20488 33324 20516
rect 32999 20485 33011 20488
rect 32953 20479 33011 20485
rect 33318 20476 33324 20488
rect 33376 20476 33382 20528
rect 34790 20476 34796 20528
rect 34848 20516 34854 20528
rect 36265 20519 36323 20525
rect 36265 20516 36277 20519
rect 34848 20488 36277 20516
rect 34848 20476 34854 20488
rect 36265 20485 36277 20488
rect 36311 20485 36323 20519
rect 36265 20479 36323 20485
rect 37182 20476 37188 20528
rect 37240 20516 37246 20528
rect 39942 20516 39948 20528
rect 37240 20488 39948 20516
rect 37240 20476 37246 20488
rect 32677 20451 32735 20457
rect 32677 20417 32689 20451
rect 32723 20417 32735 20451
rect 32677 20411 32735 20417
rect 33045 20451 33103 20457
rect 33045 20417 33057 20451
rect 33091 20448 33103 20451
rect 33134 20448 33140 20460
rect 33091 20420 33140 20448
rect 33091 20417 33103 20420
rect 33045 20411 33103 20417
rect 33134 20408 33140 20420
rect 33192 20448 33198 20460
rect 34422 20448 34428 20460
rect 33192 20420 34428 20448
rect 33192 20408 33198 20420
rect 34422 20408 34428 20420
rect 34480 20408 34486 20460
rect 35181 20451 35239 20457
rect 35181 20417 35193 20451
rect 35227 20448 35239 20451
rect 35342 20448 35348 20460
rect 35227 20420 35348 20448
rect 35227 20417 35239 20420
rect 35181 20411 35239 20417
rect 35342 20408 35348 20420
rect 35400 20408 35406 20460
rect 37292 20457 37320 20488
rect 38856 20460 38884 20488
rect 39942 20476 39948 20488
rect 40000 20476 40006 20528
rect 40494 20476 40500 20528
rect 40552 20516 40558 20528
rect 40773 20519 40831 20525
rect 40773 20516 40785 20519
rect 40552 20488 40785 20516
rect 40552 20476 40558 20488
rect 40773 20485 40785 20488
rect 40819 20485 40831 20519
rect 40773 20479 40831 20485
rect 35437 20451 35495 20457
rect 35437 20417 35449 20451
rect 35483 20448 35495 20451
rect 37277 20451 37335 20457
rect 37277 20448 37289 20451
rect 35483 20420 37289 20448
rect 35483 20417 35495 20420
rect 35437 20411 35495 20417
rect 37277 20417 37289 20420
rect 37323 20417 37335 20451
rect 37277 20411 37335 20417
rect 37544 20451 37602 20457
rect 37544 20417 37556 20451
rect 37590 20448 37602 20451
rect 38746 20448 38752 20460
rect 37590 20420 38752 20448
rect 37590 20417 37602 20420
rect 37544 20411 37602 20417
rect 38746 20408 38752 20420
rect 38804 20408 38810 20460
rect 38838 20408 38844 20460
rect 38896 20408 38902 20460
rect 39108 20451 39166 20457
rect 39108 20417 39120 20451
rect 39154 20448 39166 20451
rect 40681 20451 40739 20457
rect 39154 20420 40356 20448
rect 39154 20417 39166 20420
rect 39108 20411 39166 20417
rect 25866 20380 25872 20392
rect 25792 20352 25872 20380
rect 25866 20340 25872 20352
rect 25924 20340 25930 20392
rect 27893 20383 27951 20389
rect 27893 20349 27905 20383
rect 27939 20349 27951 20383
rect 27893 20343 27951 20349
rect 26970 20312 26976 20324
rect 25608 20284 26976 20312
rect 15841 20275 15899 20281
rect 26970 20272 26976 20284
rect 27028 20312 27034 20324
rect 27614 20312 27620 20324
rect 27028 20284 27620 20312
rect 27028 20272 27034 20284
rect 27614 20272 27620 20284
rect 27672 20272 27678 20324
rect 2961 20247 3019 20253
rect 2961 20213 2973 20247
rect 3007 20244 3019 20247
rect 3050 20244 3056 20256
rect 3007 20216 3056 20244
rect 3007 20213 3019 20216
rect 2961 20207 3019 20213
rect 3050 20204 3056 20216
rect 3108 20244 3114 20256
rect 3694 20244 3700 20256
rect 3108 20216 3700 20244
rect 3108 20204 3114 20216
rect 3694 20204 3700 20216
rect 3752 20204 3758 20256
rect 5258 20204 5264 20256
rect 5316 20204 5322 20256
rect 6733 20247 6791 20253
rect 6733 20213 6745 20247
rect 6779 20244 6791 20247
rect 6822 20244 6828 20256
rect 6779 20216 6828 20244
rect 6779 20213 6791 20216
rect 6733 20207 6791 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 16485 20247 16543 20253
rect 16485 20213 16497 20247
rect 16531 20244 16543 20247
rect 17126 20244 17132 20256
rect 16531 20216 17132 20244
rect 16531 20213 16543 20216
rect 16485 20207 16543 20213
rect 17126 20204 17132 20216
rect 17184 20204 17190 20256
rect 20070 20204 20076 20256
rect 20128 20204 20134 20256
rect 21821 20247 21879 20253
rect 21821 20213 21833 20247
rect 21867 20244 21879 20247
rect 22002 20244 22008 20256
rect 21867 20216 22008 20244
rect 21867 20213 21879 20216
rect 21821 20207 21879 20213
rect 22002 20204 22008 20216
rect 22060 20204 22066 20256
rect 26878 20204 26884 20256
rect 26936 20244 26942 20256
rect 27433 20247 27491 20253
rect 27433 20244 27445 20247
rect 26936 20216 27445 20244
rect 26936 20204 26942 20216
rect 27433 20213 27445 20216
rect 27479 20213 27491 20247
rect 27908 20244 27936 20343
rect 28074 20340 28080 20392
rect 28132 20340 28138 20392
rect 28629 20383 28687 20389
rect 28629 20349 28641 20383
rect 28675 20380 28687 20383
rect 29086 20380 29092 20392
rect 28675 20352 29092 20380
rect 28675 20349 28687 20352
rect 28629 20343 28687 20349
rect 29086 20340 29092 20352
rect 29144 20340 29150 20392
rect 30098 20340 30104 20392
rect 30156 20340 30162 20392
rect 32122 20340 32128 20392
rect 32180 20380 32186 20392
rect 33321 20383 33379 20389
rect 33321 20380 33333 20383
rect 32180 20352 33333 20380
rect 32180 20340 32186 20352
rect 33321 20349 33333 20352
rect 33367 20380 33379 20383
rect 33502 20380 33508 20392
rect 33367 20352 33508 20380
rect 33367 20349 33379 20352
rect 33321 20343 33379 20349
rect 33502 20340 33508 20352
rect 33560 20340 33566 20392
rect 35529 20383 35587 20389
rect 35529 20349 35541 20383
rect 35575 20349 35587 20383
rect 35529 20343 35587 20349
rect 29270 20244 29276 20256
rect 27908 20216 29276 20244
rect 27433 20207 27491 20213
rect 29270 20204 29276 20216
rect 29328 20204 29334 20256
rect 33229 20247 33287 20253
rect 33229 20213 33241 20247
rect 33275 20244 33287 20247
rect 33870 20244 33876 20256
rect 33275 20216 33876 20244
rect 33275 20213 33287 20216
rect 33229 20207 33287 20213
rect 33870 20204 33876 20216
rect 33928 20204 33934 20256
rect 33962 20204 33968 20256
rect 34020 20204 34026 20256
rect 34057 20247 34115 20253
rect 34057 20213 34069 20247
rect 34103 20244 34115 20247
rect 34146 20244 34152 20256
rect 34103 20216 34152 20244
rect 34103 20213 34115 20216
rect 34057 20207 34115 20213
rect 34146 20204 34152 20216
rect 34204 20244 34210 20256
rect 35544 20244 35572 20343
rect 36906 20340 36912 20392
rect 36964 20340 36970 20392
rect 40328 20321 40356 20420
rect 40681 20417 40693 20451
rect 40727 20448 40739 20451
rect 40954 20448 40960 20460
rect 40727 20420 40960 20448
rect 40727 20417 40739 20420
rect 40681 20411 40739 20417
rect 40954 20408 40960 20420
rect 41012 20408 41018 20460
rect 41506 20408 41512 20460
rect 41564 20408 41570 20460
rect 40402 20340 40408 20392
rect 40460 20380 40466 20392
rect 40865 20383 40923 20389
rect 40865 20380 40877 20383
rect 40460 20352 40877 20380
rect 40460 20340 40466 20352
rect 40865 20349 40877 20352
rect 40911 20349 40923 20383
rect 40865 20343 40923 20349
rect 41690 20340 41696 20392
rect 41748 20340 41754 20392
rect 40313 20315 40371 20321
rect 40313 20281 40325 20315
rect 40359 20281 40371 20315
rect 40313 20275 40371 20281
rect 34204 20216 35572 20244
rect 34204 20204 34210 20216
rect 36170 20204 36176 20256
rect 36228 20204 36234 20256
rect 38657 20247 38715 20253
rect 38657 20213 38669 20247
rect 38703 20244 38715 20247
rect 39022 20244 39028 20256
rect 38703 20216 39028 20244
rect 38703 20213 38715 20216
rect 38657 20207 38715 20213
rect 39022 20204 39028 20216
rect 39080 20204 39086 20256
rect 1104 20154 42504 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 42504 20154
rect 1104 20080 42504 20102
rect 3605 20043 3663 20049
rect 3605 20009 3617 20043
rect 3651 20040 3663 20043
rect 3878 20040 3884 20052
rect 3651 20012 3884 20040
rect 3651 20009 3663 20012
rect 3605 20003 3663 20009
rect 3878 20000 3884 20012
rect 3936 20000 3942 20052
rect 4249 20043 4307 20049
rect 4249 20009 4261 20043
rect 4295 20040 4307 20043
rect 4706 20040 4712 20052
rect 4295 20012 4712 20040
rect 4295 20009 4307 20012
rect 4249 20003 4307 20009
rect 4706 20000 4712 20012
rect 4764 20000 4770 20052
rect 5813 20043 5871 20049
rect 5813 20009 5825 20043
rect 5859 20040 5871 20043
rect 6454 20040 6460 20052
rect 5859 20012 6460 20040
rect 5859 20009 5871 20012
rect 5813 20003 5871 20009
rect 6454 20000 6460 20012
rect 6512 20040 6518 20052
rect 10042 20040 10048 20052
rect 6512 20012 10048 20040
rect 6512 20000 6518 20012
rect 10042 20000 10048 20012
rect 10100 20000 10106 20052
rect 11425 20043 11483 20049
rect 11425 20009 11437 20043
rect 11471 20040 11483 20043
rect 11790 20040 11796 20052
rect 11471 20012 11796 20040
rect 11471 20009 11483 20012
rect 11425 20003 11483 20009
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 17310 20000 17316 20052
rect 17368 20000 17374 20052
rect 19245 20043 19303 20049
rect 19245 20009 19257 20043
rect 19291 20040 19303 20043
rect 19334 20040 19340 20052
rect 19291 20012 19340 20040
rect 19291 20009 19303 20012
rect 19245 20003 19303 20009
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 19705 20043 19763 20049
rect 19705 20009 19717 20043
rect 19751 20040 19763 20043
rect 20530 20040 20536 20052
rect 19751 20012 20536 20040
rect 19751 20009 19763 20012
rect 19705 20003 19763 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 28994 20040 29000 20052
rect 23308 20012 29000 20040
rect 6638 19972 6644 19984
rect 5644 19944 6644 19972
rect 5644 19913 5672 19944
rect 6638 19932 6644 19944
rect 6696 19972 6702 19984
rect 8386 19972 8392 19984
rect 6696 19944 8392 19972
rect 6696 19932 6702 19944
rect 8386 19932 8392 19944
rect 8444 19972 8450 19984
rect 8444 19944 8984 19972
rect 8444 19932 8450 19944
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19873 5687 19907
rect 6086 19904 6092 19916
rect 5629 19867 5687 19873
rect 5920 19876 6092 19904
rect 1670 19796 1676 19848
rect 1728 19836 1734 19848
rect 2225 19839 2283 19845
rect 2225 19836 2237 19839
rect 1728 19808 2237 19836
rect 1728 19796 1734 19808
rect 2225 19805 2237 19808
rect 2271 19836 2283 19839
rect 3234 19836 3240 19848
rect 2271 19808 3240 19836
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 3694 19796 3700 19848
rect 3752 19836 3758 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3752 19808 3985 19836
rect 3752 19796 3758 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 4154 19796 4160 19848
rect 4212 19796 4218 19848
rect 5920 19845 5948 19876
rect 6086 19864 6092 19876
rect 6144 19904 6150 19916
rect 6822 19904 6828 19916
rect 6144 19876 6828 19904
rect 6144 19864 6150 19876
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 8956 19913 8984 19944
rect 10502 19932 10508 19984
rect 10560 19932 10566 19984
rect 11606 19932 11612 19984
rect 11664 19932 11670 19984
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19904 8263 19907
rect 8941 19907 8999 19913
rect 8251 19876 8524 19904
rect 8251 19873 8263 19876
rect 8205 19867 8263 19873
rect 8496 19848 8524 19876
rect 8941 19873 8953 19907
rect 8987 19873 8999 19907
rect 11624 19904 11652 19932
rect 11977 19907 12035 19913
rect 11977 19904 11989 19907
rect 11624 19876 11989 19904
rect 8941 19867 8999 19873
rect 11977 19873 11989 19876
rect 12023 19873 12035 19907
rect 11977 19867 12035 19873
rect 17865 19907 17923 19913
rect 17865 19873 17877 19907
rect 17911 19904 17923 19907
rect 18046 19904 18052 19916
rect 17911 19876 18052 19904
rect 17911 19873 17923 19876
rect 17865 19867 17923 19873
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19805 5779 19839
rect 5721 19799 5779 19805
rect 5905 19839 5963 19845
rect 5905 19805 5917 19839
rect 5951 19805 5963 19839
rect 6733 19839 6791 19845
rect 6733 19836 6745 19839
rect 5905 19799 5963 19805
rect 6104 19808 6745 19836
rect 2492 19771 2550 19777
rect 2492 19737 2504 19771
rect 2538 19768 2550 19771
rect 2538 19740 2774 19768
rect 2538 19737 2550 19740
rect 2492 19731 2550 19737
rect 2746 19700 2774 19740
rect 3050 19728 3056 19780
rect 3108 19768 3114 19780
rect 3789 19771 3847 19777
rect 3789 19768 3801 19771
rect 3108 19740 3801 19768
rect 3108 19728 3114 19740
rect 3789 19737 3801 19740
rect 3835 19737 3847 19771
rect 3789 19731 3847 19737
rect 4338 19728 4344 19780
rect 4396 19768 4402 19780
rect 5362 19771 5420 19777
rect 5362 19768 5374 19771
rect 4396 19740 5374 19768
rect 4396 19728 4402 19740
rect 5362 19737 5374 19740
rect 5408 19737 5420 19771
rect 5736 19768 5764 19799
rect 6104 19768 6132 19808
rect 6733 19805 6745 19808
rect 6779 19805 6791 19839
rect 8110 19836 8116 19848
rect 6733 19799 6791 19805
rect 7024 19808 8116 19836
rect 5736 19740 6132 19768
rect 5362 19731 5420 19737
rect 5920 19712 5948 19740
rect 6362 19728 6368 19780
rect 6420 19728 6426 19780
rect 6641 19771 6699 19777
rect 6641 19737 6653 19771
rect 6687 19768 6699 19771
rect 6822 19768 6828 19780
rect 6687 19740 6828 19768
rect 6687 19737 6699 19740
rect 6641 19731 6699 19737
rect 6822 19728 6828 19740
rect 6880 19728 6886 19780
rect 7024 19712 7052 19808
rect 8110 19796 8116 19808
rect 8168 19796 8174 19848
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 8297 19799 8355 19805
rect 7098 19728 7104 19780
rect 7156 19728 7162 19780
rect 4614 19700 4620 19712
rect 2746 19672 4620 19700
rect 4614 19660 4620 19672
rect 4672 19660 4678 19712
rect 5902 19660 5908 19712
rect 5960 19660 5966 19712
rect 6454 19660 6460 19712
rect 6512 19700 6518 19712
rect 6549 19703 6607 19709
rect 6549 19700 6561 19703
rect 6512 19672 6561 19700
rect 6512 19660 6518 19672
rect 6549 19669 6561 19672
rect 6595 19669 6607 19703
rect 6549 19663 6607 19669
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7006 19700 7012 19712
rect 6963 19672 7012 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7006 19660 7012 19672
rect 7064 19660 7070 19712
rect 7190 19660 7196 19712
rect 7248 19660 7254 19712
rect 8312 19700 8340 19799
rect 8478 19796 8484 19848
rect 8536 19796 8542 19848
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 8662 19836 8668 19848
rect 8619 19808 8668 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 8662 19796 8668 19808
rect 8720 19796 8726 19848
rect 8956 19836 8984 19867
rect 9766 19836 9772 19848
rect 8956 19808 9772 19836
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 10134 19796 10140 19848
rect 10192 19836 10198 19848
rect 10873 19839 10931 19845
rect 10873 19836 10885 19839
rect 10192 19808 10885 19836
rect 10192 19796 10198 19808
rect 10873 19805 10885 19808
rect 10919 19836 10931 19839
rect 10962 19836 10968 19848
rect 10919 19808 10968 19836
rect 10919 19805 10931 19808
rect 10873 19799 10931 19805
rect 10962 19796 10968 19808
rect 11020 19836 11026 19848
rect 11333 19839 11391 19845
rect 11333 19836 11345 19839
rect 11020 19808 11345 19836
rect 11020 19796 11026 19808
rect 11333 19805 11345 19808
rect 11379 19805 11391 19839
rect 11333 19799 11391 19805
rect 11514 19796 11520 19848
rect 11572 19796 11578 19848
rect 11606 19796 11612 19848
rect 11664 19796 11670 19848
rect 11992 19836 12020 19867
rect 18046 19864 18052 19876
rect 18104 19864 18110 19916
rect 18598 19864 18604 19916
rect 18656 19904 18662 19916
rect 18693 19907 18751 19913
rect 18693 19904 18705 19907
rect 18656 19876 18705 19904
rect 18656 19864 18662 19876
rect 18693 19873 18705 19876
rect 18739 19873 18751 19907
rect 20622 19904 20628 19916
rect 18693 19867 18751 19873
rect 19444 19876 20628 19904
rect 13814 19836 13820 19848
rect 11992 19808 13820 19836
rect 13814 19796 13820 19808
rect 13872 19836 13878 19848
rect 14458 19836 14464 19848
rect 13872 19808 14464 19836
rect 13872 19796 13878 19808
rect 14458 19796 14464 19808
rect 14516 19836 14522 19848
rect 14829 19839 14887 19845
rect 14829 19836 14841 19839
rect 14516 19808 14841 19836
rect 14516 19796 14522 19808
rect 14829 19805 14841 19808
rect 14875 19836 14887 19839
rect 15473 19839 15531 19845
rect 15473 19836 15485 19839
rect 14875 19808 15485 19836
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 15473 19805 15485 19808
rect 15519 19805 15531 19839
rect 18414 19836 18420 19848
rect 15473 19799 15531 19805
rect 17144 19808 18420 19836
rect 8757 19771 8815 19777
rect 8757 19737 8769 19771
rect 8803 19768 8815 19771
rect 9186 19771 9244 19777
rect 9186 19768 9198 19771
rect 8803 19740 9198 19768
rect 8803 19737 8815 19740
rect 8757 19731 8815 19737
rect 9186 19737 9198 19740
rect 9232 19737 9244 19771
rect 9186 19731 9244 19737
rect 9306 19728 9312 19780
rect 9364 19768 9370 19780
rect 12250 19777 12256 19780
rect 9364 19740 12204 19768
rect 9364 19728 9370 19740
rect 8846 19700 8852 19712
rect 8312 19672 8852 19700
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 10321 19703 10379 19709
rect 10321 19700 10333 19703
rect 9732 19672 10333 19700
rect 9732 19660 9738 19672
rect 10321 19669 10333 19672
rect 10367 19669 10379 19703
rect 10321 19663 10379 19669
rect 10410 19660 10416 19712
rect 10468 19660 10474 19712
rect 11793 19703 11851 19709
rect 11793 19669 11805 19703
rect 11839 19700 11851 19703
rect 12066 19700 12072 19712
rect 11839 19672 12072 19700
rect 11839 19669 11851 19672
rect 11793 19663 11851 19669
rect 12066 19660 12072 19672
rect 12124 19660 12130 19712
rect 12176 19700 12204 19740
rect 12244 19731 12256 19777
rect 12250 19728 12256 19731
rect 12308 19728 12314 19780
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 12406 19740 14105 19768
rect 12406 19700 12434 19740
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14093 19731 14151 19737
rect 15746 19728 15752 19780
rect 15804 19728 15810 19780
rect 16206 19768 16212 19780
rect 16132 19740 16212 19768
rect 12176 19672 12434 19700
rect 13170 19660 13176 19712
rect 13228 19700 13234 19712
rect 13357 19703 13415 19709
rect 13357 19700 13369 19703
rect 13228 19672 13369 19700
rect 13228 19660 13234 19672
rect 13357 19669 13369 19672
rect 13403 19669 13415 19703
rect 16132 19700 16160 19740
rect 16206 19728 16212 19740
rect 16264 19728 16270 19780
rect 17144 19700 17172 19808
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 19444 19845 19472 19876
rect 20622 19864 20628 19876
rect 20680 19864 20686 19916
rect 22002 19864 22008 19916
rect 22060 19864 22066 19916
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 17681 19771 17739 19777
rect 17681 19737 17693 19771
rect 17727 19768 17739 19771
rect 18141 19771 18199 19777
rect 18141 19768 18153 19771
rect 17727 19740 18153 19768
rect 17727 19737 17739 19740
rect 17681 19731 17739 19737
rect 18141 19737 18153 19740
rect 18187 19737 18199 19771
rect 18141 19731 18199 19737
rect 18598 19728 18604 19780
rect 18656 19768 18662 19780
rect 19536 19768 19564 19799
rect 19794 19796 19800 19848
rect 19852 19796 19858 19848
rect 23308 19845 23336 20012
rect 28994 20000 29000 20012
rect 29052 20000 29058 20052
rect 31938 20000 31944 20052
rect 31996 20040 32002 20052
rect 33042 20040 33048 20052
rect 31996 20012 33048 20040
rect 31996 20000 32002 20012
rect 33042 20000 33048 20012
rect 33100 20000 33106 20052
rect 35342 20000 35348 20052
rect 35400 20040 35406 20052
rect 36173 20043 36231 20049
rect 36173 20040 36185 20043
rect 35400 20012 36185 20040
rect 35400 20000 35406 20012
rect 36173 20009 36185 20012
rect 36219 20009 36231 20043
rect 36173 20003 36231 20009
rect 37918 20000 37924 20052
rect 37976 20040 37982 20052
rect 41690 20040 41696 20052
rect 37976 20012 41696 20040
rect 37976 20000 37982 20012
rect 41690 20000 41696 20012
rect 41748 20000 41754 20052
rect 32401 19975 32459 19981
rect 32401 19941 32413 19975
rect 32447 19972 32459 19975
rect 32447 19944 33364 19972
rect 32447 19941 32459 19944
rect 32401 19935 32459 19941
rect 26605 19907 26663 19913
rect 26605 19873 26617 19907
rect 26651 19904 26663 19907
rect 28350 19904 28356 19916
rect 26651 19876 28356 19904
rect 26651 19873 26663 19876
rect 26605 19867 26663 19873
rect 28350 19864 28356 19876
rect 28408 19864 28414 19916
rect 32858 19864 32864 19916
rect 32916 19904 32922 19916
rect 32953 19907 33011 19913
rect 32953 19904 32965 19907
rect 32916 19876 32965 19904
rect 32916 19864 32922 19876
rect 32953 19873 32965 19876
rect 32999 19873 33011 19907
rect 32953 19867 33011 19873
rect 33042 19864 33048 19916
rect 33100 19864 33106 19916
rect 33336 19913 33364 19944
rect 33321 19907 33379 19913
rect 33321 19873 33333 19907
rect 33367 19873 33379 19907
rect 33321 19867 33379 19873
rect 33870 19864 33876 19916
rect 33928 19904 33934 19916
rect 33928 19876 34836 19904
rect 33928 19864 33934 19876
rect 22281 19839 22339 19845
rect 22281 19805 22293 19839
rect 22327 19805 22339 19839
rect 22281 19799 22339 19805
rect 23293 19839 23351 19845
rect 23293 19805 23305 19839
rect 23339 19805 23351 19839
rect 23293 19799 23351 19805
rect 20438 19768 20444 19780
rect 18656 19740 20444 19768
rect 18656 19728 18662 19740
rect 20438 19728 20444 19740
rect 20496 19728 20502 19780
rect 20714 19728 20720 19780
rect 20772 19768 20778 19780
rect 22296 19768 22324 19799
rect 23750 19796 23756 19848
rect 23808 19836 23814 19848
rect 24029 19839 24087 19845
rect 24029 19836 24041 19839
rect 23808 19808 24041 19836
rect 23808 19796 23814 19808
rect 24029 19805 24041 19808
rect 24075 19805 24087 19839
rect 24029 19799 24087 19805
rect 31021 19839 31079 19845
rect 31021 19805 31033 19839
rect 31067 19805 31079 19839
rect 31021 19799 31079 19805
rect 22462 19768 22468 19780
rect 20772 19740 20838 19768
rect 22296 19740 22468 19768
rect 20772 19728 20778 19740
rect 22462 19728 22468 19740
rect 22520 19728 22526 19780
rect 26878 19728 26884 19780
rect 26936 19728 26942 19780
rect 28994 19768 29000 19780
rect 28106 19740 29000 19768
rect 28994 19728 29000 19740
rect 29052 19768 29058 19780
rect 29178 19768 29184 19780
rect 29052 19740 29184 19768
rect 29052 19728 29058 19740
rect 29178 19728 29184 19740
rect 29236 19728 29242 19780
rect 16132 19672 17172 19700
rect 13357 19663 13415 19669
rect 17218 19660 17224 19712
rect 17276 19660 17282 19712
rect 17770 19660 17776 19712
rect 17828 19660 17834 19712
rect 20533 19703 20591 19709
rect 20533 19669 20545 19703
rect 20579 19700 20591 19703
rect 21082 19700 21088 19712
rect 20579 19672 21088 19700
rect 20579 19669 20591 19672
rect 20533 19663 20591 19669
rect 21082 19660 21088 19672
rect 21140 19700 21146 19712
rect 21818 19700 21824 19712
rect 21140 19672 21824 19700
rect 21140 19660 21146 19672
rect 21818 19660 21824 19672
rect 21876 19660 21882 19712
rect 23474 19660 23480 19712
rect 23532 19660 23538 19712
rect 23566 19660 23572 19712
rect 23624 19700 23630 19712
rect 25038 19700 25044 19712
rect 23624 19672 25044 19700
rect 23624 19660 23630 19672
rect 25038 19660 25044 19672
rect 25096 19700 25102 19712
rect 25498 19700 25504 19712
rect 25096 19672 25504 19700
rect 25096 19660 25102 19672
rect 25498 19660 25504 19672
rect 25556 19660 25562 19712
rect 27706 19660 27712 19712
rect 27764 19700 27770 19712
rect 28353 19703 28411 19709
rect 28353 19700 28365 19703
rect 27764 19672 28365 19700
rect 27764 19660 27770 19672
rect 28353 19669 28365 19672
rect 28399 19669 28411 19703
rect 28353 19663 28411 19669
rect 29822 19660 29828 19712
rect 29880 19700 29886 19712
rect 31036 19700 31064 19799
rect 34422 19796 34428 19848
rect 34480 19796 34486 19848
rect 34698 19796 34704 19848
rect 34756 19796 34762 19848
rect 34808 19836 34836 19876
rect 36170 19864 36176 19916
rect 36228 19904 36234 19916
rect 36228 19876 36768 19904
rect 36228 19864 36234 19876
rect 34957 19839 35015 19845
rect 34957 19836 34969 19839
rect 34808 19808 34969 19836
rect 34957 19805 34969 19808
rect 35003 19805 35015 19839
rect 34957 19799 35015 19805
rect 36357 19839 36415 19845
rect 36357 19805 36369 19839
rect 36403 19805 36415 19839
rect 36357 19799 36415 19805
rect 36449 19839 36507 19845
rect 36449 19805 36461 19839
rect 36495 19836 36507 19839
rect 36630 19836 36636 19848
rect 36495 19808 36636 19836
rect 36495 19805 36507 19808
rect 36449 19799 36507 19805
rect 31288 19771 31346 19777
rect 31288 19737 31300 19771
rect 31334 19768 31346 19771
rect 34440 19768 34468 19796
rect 36372 19768 36400 19799
rect 36630 19796 36636 19808
rect 36688 19796 36694 19848
rect 36740 19845 36768 19876
rect 38838 19864 38844 19916
rect 38896 19904 38902 19916
rect 39945 19907 40003 19913
rect 39945 19904 39957 19907
rect 38896 19876 39957 19904
rect 38896 19864 38902 19876
rect 39945 19873 39957 19876
rect 39991 19873 40003 19907
rect 39945 19867 40003 19873
rect 36725 19839 36783 19845
rect 36725 19805 36737 19839
rect 36771 19805 36783 19839
rect 36725 19799 36783 19805
rect 39022 19796 39028 19848
rect 39080 19796 39086 19848
rect 31334 19740 32536 19768
rect 34440 19740 36400 19768
rect 31334 19737 31346 19740
rect 31288 19731 31346 19737
rect 31754 19700 31760 19712
rect 29880 19672 31760 19700
rect 29880 19660 29886 19672
rect 31754 19660 31760 19672
rect 31812 19660 31818 19712
rect 32508 19709 32536 19740
rect 36538 19728 36544 19780
rect 36596 19728 36602 19780
rect 38134 19740 38424 19768
rect 32493 19703 32551 19709
rect 32493 19669 32505 19703
rect 32539 19669 32551 19703
rect 32493 19663 32551 19669
rect 32861 19703 32919 19709
rect 32861 19669 32873 19703
rect 32907 19700 32919 19703
rect 33965 19703 34023 19709
rect 33965 19700 33977 19703
rect 32907 19672 33977 19700
rect 32907 19669 32919 19672
rect 32861 19663 32919 19669
rect 33965 19669 33977 19672
rect 34011 19700 34023 19703
rect 34422 19700 34428 19712
rect 34011 19672 34428 19700
rect 34011 19669 34023 19672
rect 33965 19663 34023 19669
rect 34422 19660 34428 19672
rect 34480 19660 34486 19712
rect 36081 19703 36139 19709
rect 36081 19669 36093 19703
rect 36127 19700 36139 19703
rect 36906 19700 36912 19712
rect 36127 19672 36912 19700
rect 36127 19669 36139 19672
rect 36081 19663 36139 19669
rect 36906 19660 36912 19672
rect 36964 19660 36970 19712
rect 37093 19703 37151 19709
rect 37093 19669 37105 19703
rect 37139 19700 37151 19703
rect 37182 19700 37188 19712
rect 37139 19672 37188 19700
rect 37139 19669 37151 19672
rect 37093 19663 37151 19669
rect 37182 19660 37188 19672
rect 37240 19660 37246 19712
rect 38396 19700 38424 19740
rect 38470 19728 38476 19780
rect 38528 19768 38534 19780
rect 38565 19771 38623 19777
rect 38565 19768 38577 19771
rect 38528 19740 38577 19768
rect 38528 19728 38534 19740
rect 38565 19737 38577 19740
rect 38611 19737 38623 19771
rect 38565 19731 38623 19737
rect 40218 19728 40224 19780
rect 40276 19728 40282 19780
rect 41230 19728 41236 19780
rect 41288 19728 41294 19780
rect 38654 19700 38660 19712
rect 38396 19672 38660 19700
rect 38654 19660 38660 19672
rect 38712 19660 38718 19712
rect 39574 19660 39580 19712
rect 39632 19660 39638 19712
rect 40862 19660 40868 19712
rect 40920 19700 40926 19712
rect 41693 19703 41751 19709
rect 41693 19700 41705 19703
rect 40920 19672 41705 19700
rect 40920 19660 40926 19672
rect 41693 19669 41705 19672
rect 41739 19669 41751 19703
rect 41693 19663 41751 19669
rect 1104 19610 42504 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 42504 19610
rect 1104 19536 42504 19558
rect 1765 19499 1823 19505
rect 1765 19465 1777 19499
rect 1811 19496 1823 19499
rect 1854 19496 1860 19508
rect 1811 19468 1860 19496
rect 1811 19465 1823 19468
rect 1765 19459 1823 19465
rect 1854 19456 1860 19468
rect 1912 19456 1918 19508
rect 3050 19496 3056 19508
rect 1964 19468 3056 19496
rect 1964 19369 1992 19468
rect 3050 19456 3056 19468
rect 3108 19456 3114 19508
rect 8294 19496 8300 19508
rect 3160 19468 8300 19496
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 3160 19428 3188 19468
rect 8294 19456 8300 19468
rect 8352 19496 8358 19508
rect 9122 19496 9128 19508
rect 8352 19468 9128 19496
rect 8352 19456 8358 19468
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 9677 19499 9735 19505
rect 9677 19465 9689 19499
rect 9723 19496 9735 19499
rect 10502 19496 10508 19508
rect 9723 19468 10508 19496
rect 9723 19465 9735 19468
rect 9677 19459 9735 19465
rect 10502 19456 10508 19468
rect 10560 19456 10566 19508
rect 10870 19456 10876 19508
rect 10928 19496 10934 19508
rect 11149 19499 11207 19505
rect 11149 19496 11161 19499
rect 10928 19468 11161 19496
rect 10928 19456 10934 19468
rect 11149 19465 11161 19468
rect 11195 19465 11207 19499
rect 11149 19459 11207 19465
rect 12250 19456 12256 19508
rect 12308 19496 12314 19508
rect 12437 19499 12495 19505
rect 12437 19496 12449 19499
rect 12308 19468 12449 19496
rect 12308 19456 12314 19468
rect 12437 19465 12449 19468
rect 12483 19465 12495 19499
rect 12437 19459 12495 19465
rect 15746 19456 15752 19508
rect 15804 19496 15810 19508
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 15804 19468 16681 19496
rect 15804 19456 15810 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 16669 19459 16727 19465
rect 17126 19456 17132 19508
rect 17184 19456 17190 19508
rect 17770 19496 17776 19508
rect 17604 19468 17776 19496
rect 2547 19400 3188 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 3234 19388 3240 19440
rect 3292 19388 3298 19440
rect 4154 19388 4160 19440
rect 4212 19428 4218 19440
rect 4890 19428 4896 19440
rect 4212 19400 4896 19428
rect 4212 19388 4218 19400
rect 4890 19388 4896 19400
rect 4948 19428 4954 19440
rect 4948 19400 5028 19428
rect 4948 19388 4954 19400
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19329 2007 19363
rect 1949 19323 2007 19329
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19360 3847 19363
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 3835 19332 4261 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5000 19369 5028 19400
rect 5902 19388 5908 19440
rect 5960 19428 5966 19440
rect 7190 19428 7196 19440
rect 5960 19400 6040 19428
rect 5960 19388 5966 19400
rect 4801 19363 4859 19369
rect 4801 19360 4813 19363
rect 4764 19332 4813 19360
rect 4764 19320 4770 19332
rect 4801 19329 4813 19332
rect 4847 19329 4859 19363
rect 4801 19323 4859 19329
rect 4985 19363 5043 19369
rect 4985 19329 4997 19363
rect 5031 19329 5043 19363
rect 4985 19323 5043 19329
rect 5169 19363 5227 19369
rect 5169 19329 5181 19363
rect 5215 19360 5227 19363
rect 5258 19360 5264 19372
rect 5215 19332 5264 19360
rect 5215 19329 5227 19332
rect 5169 19323 5227 19329
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 6012 19369 6040 19400
rect 6748 19400 7196 19428
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19329 6055 19363
rect 5997 19323 6055 19329
rect 6638 19320 6644 19372
rect 6696 19320 6702 19372
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19292 2191 19295
rect 3326 19292 3332 19304
rect 2179 19264 3332 19292
rect 2179 19261 2191 19264
rect 2133 19255 2191 19261
rect 3326 19252 3332 19264
rect 3384 19252 3390 19304
rect 3881 19295 3939 19301
rect 3881 19261 3893 19295
rect 3927 19261 3939 19295
rect 3881 19255 3939 19261
rect 4157 19295 4215 19301
rect 4157 19261 4169 19295
rect 4203 19292 4215 19295
rect 4338 19292 4344 19304
rect 4203 19264 4344 19292
rect 4203 19261 4215 19264
rect 4157 19255 4215 19261
rect 3896 19224 3924 19255
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 4614 19252 4620 19304
rect 4672 19292 4678 19304
rect 5077 19295 5135 19301
rect 5077 19292 5089 19295
rect 4672 19264 5089 19292
rect 4672 19252 4678 19264
rect 5077 19261 5089 19264
rect 5123 19261 5135 19295
rect 5077 19255 5135 19261
rect 5718 19252 5724 19304
rect 5776 19252 5782 19304
rect 5813 19295 5871 19301
rect 5813 19261 5825 19295
rect 5859 19261 5871 19295
rect 5813 19255 5871 19261
rect 5905 19295 5963 19301
rect 5905 19261 5917 19295
rect 5951 19292 5963 19295
rect 6086 19292 6092 19304
rect 5951 19264 6092 19292
rect 5951 19261 5963 19264
rect 5905 19255 5963 19261
rect 4798 19224 4804 19236
rect 3896 19196 4804 19224
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 5828 19224 5856 19255
rect 6086 19252 6092 19264
rect 6144 19252 6150 19304
rect 6748 19292 6776 19400
rect 7190 19388 7196 19400
rect 7248 19388 7254 19440
rect 8662 19388 8668 19440
rect 8720 19388 8726 19440
rect 8846 19388 8852 19440
rect 8904 19428 8910 19440
rect 10036 19431 10094 19437
rect 8904 19400 9352 19428
rect 8904 19388 8910 19400
rect 6914 19369 6920 19372
rect 6908 19323 6920 19369
rect 6914 19320 6920 19323
rect 6972 19320 6978 19372
rect 8110 19320 8116 19372
rect 8168 19360 8174 19372
rect 9324 19369 9352 19400
rect 10036 19397 10048 19431
rect 10082 19428 10094 19431
rect 10410 19428 10416 19440
rect 10082 19400 10416 19428
rect 10082 19397 10094 19400
rect 10036 19391 10094 19397
rect 10410 19388 10416 19400
rect 10468 19388 10474 19440
rect 10962 19388 10968 19440
rect 11020 19428 11026 19440
rect 17037 19431 17095 19437
rect 11020 19400 11928 19428
rect 11020 19388 11026 19400
rect 9033 19363 9091 19369
rect 9033 19360 9045 19363
rect 8168 19332 9045 19360
rect 8168 19320 8174 19332
rect 9033 19329 9045 19332
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 9309 19363 9367 19369
rect 9309 19329 9321 19363
rect 9355 19360 9367 19363
rect 9674 19360 9680 19372
rect 9355 19332 9680 19360
rect 9355 19329 9367 19332
rect 9309 19323 9367 19329
rect 6656 19264 6776 19292
rect 6656 19224 6684 19264
rect 5828 19196 6684 19224
rect 6181 19159 6239 19165
rect 6181 19125 6193 19159
rect 6227 19156 6239 19159
rect 6822 19156 6828 19168
rect 6227 19128 6828 19156
rect 6227 19125 6239 19128
rect 6181 19119 6239 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 8021 19159 8079 19165
rect 8021 19125 8033 19159
rect 8067 19156 8079 19159
rect 8110 19156 8116 19168
rect 8067 19128 8116 19156
rect 8067 19125 8079 19128
rect 8021 19119 8079 19125
rect 8110 19116 8116 19128
rect 8168 19116 8174 19168
rect 9048 19156 9076 19323
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 9766 19320 9772 19372
rect 9824 19320 9830 19372
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 11790 19360 11796 19372
rect 11747 19332 11796 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 11790 19320 11796 19332
rect 11848 19320 11854 19372
rect 11900 19369 11928 19400
rect 17037 19397 17049 19431
rect 17083 19428 17095 19431
rect 17604 19428 17632 19468
rect 17770 19456 17776 19468
rect 17828 19456 17834 19508
rect 22462 19496 22468 19508
rect 17972 19468 22468 19496
rect 17972 19440 18000 19468
rect 17954 19428 17960 19440
rect 17083 19400 17632 19428
rect 17696 19400 17960 19428
rect 17083 19397 17095 19400
rect 17037 19391 17095 19397
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19360 11943 19363
rect 11931 19332 12204 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 9214 19252 9220 19304
rect 9272 19252 9278 19304
rect 9398 19252 9404 19304
rect 9456 19252 9462 19304
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19261 9551 19295
rect 9493 19255 9551 19261
rect 9508 19156 9536 19255
rect 11330 19252 11336 19304
rect 11388 19292 11394 19304
rect 11514 19292 11520 19304
rect 11388 19264 11520 19292
rect 11388 19252 11394 19264
rect 11514 19252 11520 19264
rect 11572 19292 11578 19304
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11572 19264 11989 19292
rect 11572 19252 11578 19264
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 11977 19255 12035 19261
rect 11992 19224 12020 19255
rect 12066 19252 12072 19304
rect 12124 19252 12130 19304
rect 12176 19292 12204 19332
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 13725 19363 13783 19369
rect 12308 19332 12664 19360
rect 12308 19320 12314 19332
rect 12526 19292 12532 19304
rect 12176 19264 12532 19292
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 12636 19292 12664 19332
rect 13725 19329 13737 19363
rect 13771 19360 13783 19363
rect 13814 19360 13820 19372
rect 13771 19332 13820 19360
rect 13771 19329 13783 19332
rect 13725 19323 13783 19329
rect 13814 19320 13820 19332
rect 13872 19360 13878 19372
rect 14366 19360 14372 19372
rect 13872 19332 14372 19360
rect 13872 19320 13878 19332
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 17696 19369 17724 19400
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 18414 19388 18420 19440
rect 18472 19388 18478 19440
rect 19904 19369 19932 19468
rect 20714 19388 20720 19440
rect 20772 19388 20778 19440
rect 22066 19428 22094 19468
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 25406 19456 25412 19508
rect 25464 19496 25470 19508
rect 25593 19499 25651 19505
rect 25593 19496 25605 19499
rect 25464 19468 25605 19496
rect 25464 19456 25470 19468
rect 25593 19465 25605 19468
rect 25639 19465 25651 19499
rect 25593 19459 25651 19465
rect 26421 19499 26479 19505
rect 26421 19465 26433 19499
rect 26467 19496 26479 19499
rect 26786 19496 26792 19508
rect 26467 19468 26792 19496
rect 26467 19465 26479 19468
rect 26421 19459 26479 19465
rect 26786 19456 26792 19468
rect 26844 19456 26850 19508
rect 28626 19496 28632 19508
rect 28000 19468 28632 19496
rect 23566 19428 23572 19440
rect 22020 19400 22094 19428
rect 23506 19400 23572 19428
rect 22020 19369 22048 19400
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 25498 19428 25504 19440
rect 25346 19400 25504 19428
rect 25498 19388 25504 19400
rect 25556 19388 25562 19440
rect 17681 19363 17739 19369
rect 17681 19329 17693 19363
rect 17727 19329 17739 19363
rect 17681 19323 17739 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 13446 19292 13452 19304
rect 12636 19264 13452 19292
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19292 17371 19295
rect 17957 19295 18015 19301
rect 17359 19264 17816 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 13170 19224 13176 19236
rect 11992 19196 13176 19224
rect 13170 19184 13176 19196
rect 13228 19184 13234 19236
rect 9950 19156 9956 19168
rect 9048 19128 9956 19156
rect 9950 19116 9956 19128
rect 10008 19116 10014 19168
rect 17678 19116 17684 19168
rect 17736 19156 17742 19168
rect 17788 19156 17816 19264
rect 17957 19261 17969 19295
rect 18003 19292 18015 19295
rect 18322 19292 18328 19304
rect 18003 19264 18328 19292
rect 18003 19261 18015 19264
rect 17957 19255 18015 19261
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19300 19264 19441 19292
rect 19300 19252 19306 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 20165 19295 20223 19301
rect 20165 19261 20177 19295
rect 20211 19292 20223 19295
rect 20714 19292 20720 19304
rect 20211 19264 20720 19292
rect 20211 19261 20223 19264
rect 20165 19255 20223 19261
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 21637 19295 21695 19301
rect 21637 19292 21649 19295
rect 20956 19264 21649 19292
rect 20956 19252 20962 19264
rect 21637 19261 21649 19264
rect 21683 19261 21695 19295
rect 21637 19255 21695 19261
rect 22281 19295 22339 19301
rect 22281 19261 22293 19295
rect 22327 19292 22339 19295
rect 22738 19292 22744 19304
rect 22327 19264 22744 19292
rect 22327 19261 22339 19264
rect 22281 19255 22339 19261
rect 22738 19252 22744 19264
rect 22796 19252 22802 19304
rect 23860 19292 23888 19323
rect 26326 19320 26332 19372
rect 26384 19360 26390 19372
rect 28000 19369 28028 19468
rect 28626 19456 28632 19468
rect 28684 19496 28690 19508
rect 29822 19496 29828 19508
rect 28684 19468 29828 19496
rect 28684 19456 28690 19468
rect 29822 19456 29828 19468
rect 29880 19456 29886 19508
rect 31570 19456 31576 19508
rect 31628 19456 31634 19508
rect 32122 19456 32128 19508
rect 32180 19456 32186 19508
rect 32582 19456 32588 19508
rect 32640 19496 32646 19508
rect 34698 19496 34704 19508
rect 32640 19468 34704 19496
rect 32640 19456 32646 19468
rect 28994 19388 29000 19440
rect 29052 19388 29058 19440
rect 29564 19400 30590 19428
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26384 19332 26985 19360
rect 26384 19320 26390 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 27985 19363 28043 19369
rect 27985 19329 27997 19363
rect 28031 19329 28043 19363
rect 27985 19323 28043 19329
rect 23860 19264 23980 19292
rect 23750 19184 23756 19236
rect 23808 19184 23814 19236
rect 22370 19156 22376 19168
rect 17736 19128 22376 19156
rect 17736 19116 17742 19128
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 23952 19156 23980 19264
rect 24118 19252 24124 19304
rect 24176 19252 24182 19304
rect 26510 19252 26516 19304
rect 26568 19252 26574 19304
rect 26694 19252 26700 19304
rect 26752 19292 26758 19304
rect 27525 19295 27583 19301
rect 27525 19292 27537 19295
rect 26752 19264 27537 19292
rect 26752 19252 26758 19264
rect 27525 19261 27537 19264
rect 27571 19261 27583 19295
rect 27525 19255 27583 19261
rect 28258 19252 28264 19304
rect 28316 19252 28322 19304
rect 28994 19252 29000 19304
rect 29052 19292 29058 19304
rect 29564 19292 29592 19400
rect 33134 19388 33140 19440
rect 33192 19388 33198 19440
rect 29822 19320 29828 19372
rect 29880 19320 29886 19372
rect 33888 19369 33916 19468
rect 34698 19456 34704 19468
rect 34756 19456 34762 19508
rect 36354 19456 36360 19508
rect 36412 19496 36418 19508
rect 36817 19499 36875 19505
rect 36817 19496 36829 19499
rect 36412 19468 36829 19496
rect 36412 19456 36418 19468
rect 36817 19465 36829 19468
rect 36863 19465 36875 19499
rect 36817 19459 36875 19465
rect 38470 19456 38476 19508
rect 38528 19456 38534 19508
rect 40218 19456 40224 19508
rect 40276 19456 40282 19508
rect 40681 19499 40739 19505
rect 40681 19465 40693 19499
rect 40727 19496 40739 19499
rect 40954 19496 40960 19508
rect 40727 19468 40960 19496
rect 40727 19465 40739 19468
rect 40681 19459 40739 19465
rect 40954 19456 40960 19468
rect 41012 19456 41018 19508
rect 41506 19456 41512 19508
rect 41564 19456 41570 19508
rect 33962 19388 33968 19440
rect 34020 19428 34026 19440
rect 34333 19431 34391 19437
rect 34333 19428 34345 19431
rect 34020 19400 34345 19428
rect 34020 19388 34026 19400
rect 34333 19397 34345 19400
rect 34379 19397 34391 19431
rect 34333 19391 34391 19397
rect 34422 19388 34428 19440
rect 34480 19388 34486 19440
rect 38013 19431 38071 19437
rect 38013 19397 38025 19431
rect 38059 19428 38071 19431
rect 39574 19428 39580 19440
rect 38059 19400 39580 19428
rect 38059 19397 38071 19400
rect 38013 19391 38071 19397
rect 39574 19388 39580 19400
rect 39632 19388 39638 19440
rect 33873 19363 33931 19369
rect 33873 19329 33885 19363
rect 33919 19329 33931 19363
rect 33873 19323 33931 19329
rect 29052 19264 29592 19292
rect 29052 19252 29058 19264
rect 29638 19252 29644 19304
rect 29696 19292 29702 19304
rect 29733 19295 29791 19301
rect 29733 19292 29745 19295
rect 29696 19264 29745 19292
rect 29696 19252 29702 19264
rect 29733 19261 29745 19264
rect 29779 19261 29791 19295
rect 29733 19255 29791 19261
rect 30101 19295 30159 19301
rect 30101 19261 30113 19295
rect 30147 19292 30159 19295
rect 30466 19292 30472 19304
rect 30147 19264 30472 19292
rect 30147 19261 30159 19264
rect 30101 19255 30159 19261
rect 30466 19252 30472 19264
rect 30524 19252 30530 19304
rect 33597 19295 33655 19301
rect 33597 19261 33609 19295
rect 33643 19292 33655 19295
rect 33643 19264 34008 19292
rect 33643 19261 33655 19264
rect 33597 19255 33655 19261
rect 33980 19233 34008 19264
rect 34330 19252 34336 19304
rect 34388 19292 34394 19304
rect 34609 19295 34667 19301
rect 34609 19292 34621 19295
rect 34388 19264 34621 19292
rect 34388 19252 34394 19264
rect 34609 19261 34621 19264
rect 34655 19261 34667 19295
rect 34609 19255 34667 19261
rect 33965 19227 34023 19233
rect 33965 19193 33977 19227
rect 34011 19193 34023 19227
rect 33965 19187 34023 19193
rect 25222 19156 25228 19168
rect 23952 19128 25228 19156
rect 25222 19116 25228 19128
rect 25280 19116 25286 19168
rect 25958 19116 25964 19168
rect 26016 19116 26022 19168
rect 33226 19116 33232 19168
rect 33284 19156 33290 19168
rect 34624 19156 34652 19255
rect 34698 19252 34704 19304
rect 34756 19292 34762 19304
rect 35069 19295 35127 19301
rect 35069 19292 35081 19295
rect 34756 19264 35081 19292
rect 34756 19252 34762 19264
rect 35069 19261 35081 19264
rect 35115 19261 35127 19295
rect 35069 19255 35127 19261
rect 35342 19252 35348 19304
rect 35400 19252 35406 19304
rect 36464 19292 36492 19346
rect 38102 19320 38108 19372
rect 38160 19320 38166 19372
rect 40586 19320 40592 19372
rect 40644 19320 40650 19372
rect 40862 19320 40868 19372
rect 40920 19360 40926 19372
rect 41049 19363 41107 19369
rect 41049 19360 41061 19363
rect 40920 19332 41061 19360
rect 40920 19320 40926 19332
rect 41049 19329 41061 19332
rect 41095 19329 41107 19363
rect 41049 19323 41107 19329
rect 41233 19363 41291 19369
rect 41233 19329 41245 19363
rect 41279 19329 41291 19363
rect 41233 19323 41291 19329
rect 36538 19292 36544 19304
rect 36464 19264 36544 19292
rect 36538 19252 36544 19264
rect 36596 19252 36602 19304
rect 37918 19252 37924 19304
rect 37976 19252 37982 19304
rect 40773 19295 40831 19301
rect 40773 19261 40785 19295
rect 40819 19261 40831 19295
rect 40773 19255 40831 19261
rect 40788 19156 40816 19255
rect 41046 19184 41052 19236
rect 41104 19224 41110 19236
rect 41248 19224 41276 19323
rect 42150 19252 42156 19304
rect 42208 19252 42214 19304
rect 41104 19196 41276 19224
rect 41104 19184 41110 19196
rect 33284 19128 40816 19156
rect 41141 19159 41199 19165
rect 33284 19116 33290 19128
rect 41141 19125 41153 19159
rect 41187 19156 41199 19159
rect 41322 19156 41328 19168
rect 41187 19128 41328 19156
rect 41187 19125 41199 19128
rect 41141 19119 41199 19125
rect 41322 19116 41328 19128
rect 41380 19116 41386 19168
rect 1104 19066 42504 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 42504 19066
rect 1104 18992 42504 19014
rect 4065 18955 4123 18961
rect 4065 18921 4077 18955
rect 4111 18952 4123 18955
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 4111 18924 4537 18952
rect 4111 18921 4123 18924
rect 4065 18915 4123 18921
rect 4525 18921 4537 18924
rect 4571 18952 4583 18955
rect 4706 18952 4712 18964
rect 4571 18924 4712 18952
rect 4571 18921 4583 18924
rect 4525 18915 4583 18921
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 5718 18912 5724 18964
rect 5776 18952 5782 18964
rect 6362 18952 6368 18964
rect 5776 18924 6368 18952
rect 5776 18912 5782 18924
rect 6362 18912 6368 18924
rect 6420 18912 6426 18964
rect 6822 18912 6828 18964
rect 6880 18912 6886 18964
rect 7576 18924 10088 18952
rect 3970 18884 3976 18896
rect 3896 18856 3976 18884
rect 3896 18825 3924 18856
rect 3970 18844 3976 18856
rect 4028 18844 4034 18896
rect 6641 18887 6699 18893
rect 6641 18853 6653 18887
rect 6687 18884 6699 18887
rect 6914 18884 6920 18896
rect 6687 18856 6920 18884
rect 6687 18853 6699 18856
rect 6641 18847 6699 18853
rect 6914 18844 6920 18856
rect 6972 18844 6978 18896
rect 7006 18844 7012 18896
rect 7064 18884 7070 18896
rect 7193 18887 7251 18893
rect 7193 18884 7205 18887
rect 7064 18856 7205 18884
rect 7064 18844 7070 18856
rect 7193 18853 7205 18856
rect 7239 18853 7251 18887
rect 7193 18847 7251 18853
rect 3881 18819 3939 18825
rect 3881 18785 3893 18819
rect 3927 18785 3939 18819
rect 3881 18779 3939 18785
rect 3694 18708 3700 18760
rect 3752 18748 3758 18760
rect 3789 18751 3847 18757
rect 3789 18748 3801 18751
rect 3752 18720 3801 18748
rect 3752 18708 3758 18720
rect 3789 18717 3801 18720
rect 3835 18717 3847 18751
rect 3789 18711 3847 18717
rect 3970 18708 3976 18760
rect 4028 18748 4034 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 4028 18720 4077 18748
rect 4028 18708 4034 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4798 18748 4804 18760
rect 4065 18711 4123 18717
rect 4540 18720 4804 18748
rect 4080 18680 4108 18711
rect 4540 18689 4568 18720
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 7576 18757 7604 18924
rect 9585 18887 9643 18893
rect 7668 18856 9536 18884
rect 7561 18751 7619 18757
rect 7561 18717 7573 18751
rect 7607 18717 7619 18751
rect 7561 18711 7619 18717
rect 4341 18683 4399 18689
rect 4341 18680 4353 18683
rect 4080 18652 4353 18680
rect 4341 18649 4353 18652
rect 4387 18649 4399 18683
rect 4540 18683 4599 18689
rect 4540 18652 4553 18683
rect 4341 18643 4399 18649
rect 4541 18649 4553 18652
rect 4587 18649 4599 18683
rect 7668 18680 7696 18856
rect 8113 18819 8171 18825
rect 8113 18785 8125 18819
rect 8159 18785 8171 18819
rect 8113 18779 8171 18785
rect 8297 18819 8355 18825
rect 8297 18785 8309 18819
rect 8343 18816 8355 18819
rect 8478 18816 8484 18828
rect 8343 18788 8484 18816
rect 8343 18785 8355 18788
rect 8297 18779 8355 18785
rect 4541 18643 4599 18649
rect 4632 18652 7696 18680
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 4632 18612 4660 18652
rect 7742 18640 7748 18692
rect 7800 18640 7806 18692
rect 8128 18680 8156 18779
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 9508 18816 9536 18856
rect 9585 18853 9597 18887
rect 9631 18884 9643 18887
rect 9674 18884 9680 18896
rect 9631 18856 9680 18884
rect 9631 18853 9643 18856
rect 9585 18847 9643 18853
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 10060 18884 10088 18924
rect 10134 18912 10140 18964
rect 10192 18912 10198 18964
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 10873 18955 10931 18961
rect 10873 18952 10885 18955
rect 10836 18924 10885 18952
rect 10836 18912 10842 18924
rect 10873 18921 10885 18924
rect 10919 18921 10931 18955
rect 12250 18952 12256 18964
rect 10873 18915 10931 18921
rect 12084 18924 12256 18952
rect 12084 18884 12112 18924
rect 12250 18912 12256 18924
rect 12308 18912 12314 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 17865 18955 17923 18961
rect 17865 18952 17877 18955
rect 17828 18924 17877 18952
rect 17828 18912 17834 18924
rect 17865 18921 17877 18924
rect 17911 18921 17923 18955
rect 17865 18915 17923 18921
rect 18322 18912 18328 18964
rect 18380 18912 18386 18964
rect 18414 18912 18420 18964
rect 18472 18952 18478 18964
rect 19429 18955 19487 18961
rect 19429 18952 19441 18955
rect 18472 18924 19441 18952
rect 18472 18912 18478 18924
rect 19429 18921 19441 18924
rect 19475 18921 19487 18955
rect 19429 18915 19487 18921
rect 20714 18912 20720 18964
rect 20772 18912 20778 18964
rect 22738 18912 22744 18964
rect 22796 18912 22802 18964
rect 24118 18912 24124 18964
rect 24176 18952 24182 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 24176 18924 24409 18952
rect 24176 18912 24182 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24397 18915 24455 18921
rect 24946 18912 24952 18964
rect 25004 18912 25010 18964
rect 26694 18912 26700 18964
rect 26752 18912 26758 18964
rect 28258 18912 28264 18964
rect 28316 18952 28322 18964
rect 28445 18955 28503 18961
rect 28445 18952 28457 18955
rect 28316 18924 28457 18952
rect 28316 18912 28322 18924
rect 28445 18921 28457 18924
rect 28491 18921 28503 18955
rect 28445 18915 28503 18921
rect 30466 18912 30472 18964
rect 30524 18912 30530 18964
rect 33594 18912 33600 18964
rect 33652 18952 33658 18964
rect 34333 18955 34391 18961
rect 34333 18952 34345 18955
rect 33652 18924 34345 18952
rect 33652 18912 33658 18924
rect 34333 18921 34345 18924
rect 34379 18921 34391 18955
rect 36538 18952 36544 18964
rect 34333 18915 34391 18921
rect 34440 18924 36544 18952
rect 10060 18856 12112 18884
rect 12161 18887 12219 18893
rect 12161 18853 12173 18887
rect 12207 18884 12219 18887
rect 24964 18884 24992 18912
rect 12207 18856 13860 18884
rect 12207 18853 12219 18856
rect 12161 18847 12219 18853
rect 10502 18816 10508 18828
rect 9508 18788 10508 18816
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 8386 18708 8392 18760
rect 8444 18708 8450 18760
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9272 18720 9781 18748
rect 9272 18708 9278 18720
rect 9769 18717 9781 18720
rect 9815 18748 9827 18751
rect 10042 18748 10048 18760
rect 9815 18720 10048 18748
rect 9815 18717 9827 18720
rect 9769 18711 9827 18717
rect 10042 18708 10048 18720
rect 10100 18748 10106 18760
rect 10870 18748 10876 18760
rect 10100 18720 10876 18748
rect 10100 18708 10106 18720
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11103 18720 11744 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 8662 18680 8668 18692
rect 7852 18652 8668 18680
rect 4295 18584 4660 18612
rect 4709 18615 4767 18621
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 4709 18581 4721 18615
rect 4755 18612 4767 18615
rect 4890 18612 4896 18624
rect 4755 18584 4896 18612
rect 4755 18581 4767 18584
rect 4709 18575 4767 18581
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 6825 18615 6883 18621
rect 6825 18581 6837 18615
rect 6871 18612 6883 18615
rect 7377 18615 7435 18621
rect 7377 18612 7389 18615
rect 6871 18584 7389 18612
rect 6871 18581 6883 18584
rect 6825 18575 6883 18581
rect 7377 18581 7389 18584
rect 7423 18612 7435 18615
rect 7852 18612 7880 18652
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 9950 18640 9956 18692
rect 10008 18640 10014 18692
rect 10778 18680 10784 18692
rect 10152 18652 10784 18680
rect 7423 18584 7880 18612
rect 7423 18581 7435 18584
rect 7377 18575 7435 18581
rect 7926 18572 7932 18624
rect 7984 18612 7990 18624
rect 8113 18615 8171 18621
rect 8113 18612 8125 18615
rect 7984 18584 8125 18612
rect 7984 18572 7990 18584
rect 8113 18581 8125 18584
rect 8159 18581 8171 18615
rect 8113 18575 8171 18581
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 9858 18612 9864 18624
rect 9456 18584 9864 18612
rect 9456 18572 9462 18584
rect 9858 18572 9864 18584
rect 9916 18612 9922 18624
rect 10152 18612 10180 18652
rect 10778 18640 10784 18652
rect 10836 18640 10842 18692
rect 11330 18640 11336 18692
rect 11388 18640 11394 18692
rect 11716 18680 11744 18720
rect 12066 18708 12072 18760
rect 12124 18708 12130 18760
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18748 12311 18751
rect 12360 18748 12388 18779
rect 12526 18776 12532 18828
rect 12584 18816 12590 18828
rect 12584 18788 13400 18816
rect 12584 18776 12590 18788
rect 12299 18720 12388 18748
rect 12621 18751 12679 18757
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 12621 18717 12633 18751
rect 12667 18717 12679 18751
rect 12621 18711 12679 18717
rect 12526 18680 12532 18692
rect 11716 18652 12532 18680
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 9916 18584 10180 18612
rect 9916 18572 9922 18584
rect 10226 18572 10232 18624
rect 10284 18612 10290 18624
rect 10689 18615 10747 18621
rect 10689 18612 10701 18615
rect 10284 18584 10701 18612
rect 10284 18572 10290 18584
rect 10689 18581 10701 18584
rect 10735 18581 10747 18615
rect 12636 18612 12664 18711
rect 12710 18708 12716 18760
rect 12768 18708 12774 18760
rect 12802 18708 12808 18760
rect 12860 18748 12866 18760
rect 13372 18757 13400 18788
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 12860 18720 13277 18748
rect 12860 18708 12866 18720
rect 13265 18717 13277 18720
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 13630 18748 13636 18760
rect 13587 18720 13636 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 13630 18708 13636 18720
rect 13688 18708 13694 18760
rect 13832 18757 13860 18856
rect 23308 18856 24992 18884
rect 17218 18776 17224 18828
rect 17276 18776 17282 18828
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18969 18819 19027 18825
rect 18969 18816 18981 18819
rect 18104 18788 18981 18816
rect 18104 18776 18110 18788
rect 18969 18785 18981 18788
rect 19015 18816 19027 18819
rect 21269 18819 21327 18825
rect 19015 18788 19840 18816
rect 19015 18785 19027 18788
rect 18969 18779 19027 18785
rect 13817 18751 13875 18757
rect 13817 18717 13829 18751
rect 13863 18717 13875 18751
rect 13817 18711 13875 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18748 18751 18751
rect 19242 18748 19248 18760
rect 18739 18720 19248 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 19242 18708 19248 18720
rect 19300 18708 19306 18760
rect 12728 18680 12756 18708
rect 19812 18692 19840 18788
rect 21269 18785 21281 18819
rect 21315 18785 21327 18819
rect 21269 18779 21327 18785
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20956 18720 21097 18748
rect 20956 18708 20962 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 12989 18683 13047 18689
rect 12989 18680 13001 18683
rect 12728 18652 13001 18680
rect 12989 18649 13001 18652
rect 13035 18680 13047 18683
rect 13078 18680 13084 18692
rect 13035 18652 13084 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 13078 18640 13084 18652
rect 13136 18640 13142 18692
rect 13170 18640 13176 18692
rect 13228 18640 13234 18692
rect 19702 18640 19708 18692
rect 19760 18640 19766 18692
rect 19794 18640 19800 18692
rect 19852 18680 19858 18692
rect 21284 18680 21312 18779
rect 23198 18776 23204 18828
rect 23256 18776 23262 18828
rect 23308 18825 23336 18856
rect 23293 18819 23351 18825
rect 23293 18785 23305 18819
rect 23339 18785 23351 18819
rect 24949 18819 25007 18825
rect 24949 18816 24961 18819
rect 23293 18779 23351 18785
rect 23492 18788 24961 18816
rect 23109 18751 23167 18757
rect 23109 18717 23121 18751
rect 23155 18748 23167 18751
rect 23382 18748 23388 18760
rect 23155 18720 23388 18748
rect 23155 18717 23167 18720
rect 23109 18711 23167 18717
rect 23382 18708 23388 18720
rect 23440 18708 23446 18760
rect 23492 18680 23520 18788
rect 24949 18785 24961 18788
rect 24995 18785 25007 18819
rect 24949 18779 25007 18785
rect 28074 18776 28080 18828
rect 28132 18816 28138 18828
rect 28997 18819 29055 18825
rect 28997 18816 29009 18819
rect 28132 18788 29009 18816
rect 28132 18776 28138 18788
rect 28997 18785 29009 18788
rect 29043 18816 29055 18819
rect 31018 18816 31024 18828
rect 29043 18788 31024 18816
rect 29043 18785 29055 18788
rect 28997 18779 29055 18785
rect 31018 18776 31024 18788
rect 31076 18776 31082 18828
rect 33318 18776 33324 18828
rect 33376 18816 33382 18828
rect 33376 18788 34008 18816
rect 33376 18776 33382 18788
rect 25222 18708 25228 18760
rect 25280 18748 25286 18760
rect 25317 18751 25375 18757
rect 25317 18748 25329 18751
rect 25280 18720 25329 18748
rect 25280 18708 25286 18720
rect 25317 18717 25329 18720
rect 25363 18717 25375 18751
rect 25317 18711 25375 18717
rect 25584 18751 25642 18757
rect 25584 18717 25596 18751
rect 25630 18748 25642 18751
rect 25958 18748 25964 18760
rect 25630 18720 25964 18748
rect 25630 18717 25642 18720
rect 25584 18711 25642 18717
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 28813 18751 28871 18757
rect 28813 18717 28825 18751
rect 28859 18748 28871 18751
rect 29638 18748 29644 18760
rect 28859 18720 29644 18748
rect 28859 18717 28871 18720
rect 28813 18711 28871 18717
rect 29638 18708 29644 18720
rect 29696 18708 29702 18760
rect 30837 18751 30895 18757
rect 30837 18717 30849 18751
rect 30883 18748 30895 18751
rect 31570 18748 31576 18760
rect 30883 18720 31576 18748
rect 30883 18717 30895 18720
rect 30837 18711 30895 18717
rect 31570 18708 31576 18720
rect 31628 18708 31634 18760
rect 31754 18708 31760 18760
rect 31812 18748 31818 18760
rect 32125 18751 32183 18757
rect 32125 18748 32137 18751
rect 31812 18720 32137 18748
rect 31812 18708 31818 18720
rect 32125 18717 32137 18720
rect 32171 18748 32183 18751
rect 32582 18748 32588 18760
rect 32171 18720 32588 18748
rect 32171 18717 32183 18720
rect 32125 18711 32183 18717
rect 32582 18708 32588 18720
rect 32640 18708 32646 18760
rect 33980 18748 34008 18788
rect 34440 18748 34468 18924
rect 36538 18912 36544 18924
rect 36596 18912 36602 18964
rect 38102 18912 38108 18964
rect 38160 18952 38166 18964
rect 38289 18955 38347 18961
rect 38289 18952 38301 18955
rect 38160 18924 38301 18952
rect 38160 18912 38166 18924
rect 38289 18921 38301 18924
rect 38335 18921 38347 18955
rect 38289 18915 38347 18921
rect 40586 18912 40592 18964
rect 40644 18952 40650 18964
rect 41233 18955 41291 18961
rect 41233 18952 41245 18955
rect 40644 18924 41245 18952
rect 40644 18912 40650 18924
rect 41233 18921 41245 18924
rect 41279 18921 41291 18955
rect 41233 18915 41291 18921
rect 40221 18887 40279 18893
rect 40221 18853 40233 18887
rect 40267 18884 40279 18887
rect 42058 18884 42064 18896
rect 40267 18856 42064 18884
rect 40267 18853 40279 18856
rect 40221 18847 40279 18853
rect 42058 18844 42064 18856
rect 42116 18844 42122 18896
rect 34698 18776 34704 18828
rect 34756 18816 34762 18828
rect 34977 18819 35035 18825
rect 34977 18816 34989 18819
rect 34756 18788 34989 18816
rect 34756 18776 34762 18788
rect 34977 18785 34989 18788
rect 35023 18785 35035 18819
rect 34977 18779 35035 18785
rect 37182 18776 37188 18828
rect 37240 18816 37246 18828
rect 37645 18819 37703 18825
rect 37645 18816 37657 18819
rect 37240 18788 37657 18816
rect 37240 18776 37246 18788
rect 37645 18785 37657 18788
rect 37691 18785 37703 18819
rect 41785 18819 41843 18825
rect 41785 18816 41797 18819
rect 37645 18779 37703 18785
rect 40880 18788 41797 18816
rect 40880 18760 40908 18788
rect 41785 18785 41797 18788
rect 41831 18785 41843 18819
rect 41785 18779 41843 18785
rect 33980 18734 34468 18748
rect 33994 18720 34468 18734
rect 39298 18708 39304 18760
rect 39356 18708 39362 18760
rect 40037 18751 40095 18757
rect 40037 18717 40049 18751
rect 40083 18717 40095 18751
rect 40037 18711 40095 18717
rect 40221 18751 40279 18757
rect 40221 18717 40233 18751
rect 40267 18748 40279 18751
rect 40862 18748 40868 18760
rect 40267 18720 40868 18748
rect 40267 18717 40279 18720
rect 40221 18711 40279 18717
rect 19852 18652 23520 18680
rect 19852 18640 19858 18652
rect 24394 18640 24400 18692
rect 24452 18680 24458 18692
rect 24857 18683 24915 18689
rect 24857 18680 24869 18683
rect 24452 18652 24869 18680
rect 24452 18640 24458 18652
rect 24857 18649 24869 18652
rect 24903 18649 24915 18683
rect 24857 18643 24915 18649
rect 32861 18683 32919 18689
rect 32861 18649 32873 18683
rect 32907 18680 32919 18683
rect 33134 18680 33140 18692
rect 32907 18652 33140 18680
rect 32907 18649 32919 18652
rect 32861 18643 32919 18649
rect 33134 18640 33140 18652
rect 33192 18640 33198 18692
rect 35253 18683 35311 18689
rect 35253 18649 35265 18683
rect 35299 18649 35311 18683
rect 36538 18680 36544 18692
rect 36478 18652 36544 18680
rect 35253 18643 35311 18649
rect 13188 18612 13216 18640
rect 12636 18584 13216 18612
rect 13725 18615 13783 18621
rect 10689 18575 10747 18581
rect 13725 18581 13737 18615
rect 13771 18612 13783 18615
rect 14182 18612 14188 18624
rect 13771 18584 14188 18612
rect 13771 18581 13783 18584
rect 13725 18575 13783 18581
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 18785 18615 18843 18621
rect 18785 18581 18797 18615
rect 18831 18612 18843 18615
rect 19334 18612 19340 18624
rect 18831 18584 19340 18612
rect 18831 18581 18843 18584
rect 18785 18575 18843 18581
rect 19334 18572 19340 18584
rect 19392 18572 19398 18624
rect 21177 18615 21235 18621
rect 21177 18581 21189 18615
rect 21223 18612 21235 18615
rect 21450 18612 21456 18624
rect 21223 18584 21456 18612
rect 21223 18581 21235 18584
rect 21177 18575 21235 18581
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18612 24823 18615
rect 25406 18612 25412 18624
rect 24811 18584 25412 18612
rect 24811 18581 24823 18584
rect 24765 18575 24823 18581
rect 25406 18572 25412 18584
rect 25464 18572 25470 18624
rect 28902 18572 28908 18624
rect 28960 18572 28966 18624
rect 30926 18572 30932 18624
rect 30984 18572 30990 18624
rect 35268 18612 35296 18643
rect 36538 18640 36544 18652
rect 36596 18640 36602 18692
rect 40052 18680 40080 18711
rect 40862 18708 40868 18720
rect 40920 18708 40926 18760
rect 40957 18751 41015 18757
rect 40957 18717 40969 18751
rect 41003 18748 41015 18751
rect 41598 18748 41604 18760
rect 41003 18720 41604 18748
rect 41003 18717 41015 18720
rect 40957 18711 41015 18717
rect 41598 18708 41604 18720
rect 41656 18708 41662 18760
rect 41046 18680 41052 18692
rect 40052 18652 41052 18680
rect 41046 18640 41052 18652
rect 41104 18640 41110 18692
rect 35434 18612 35440 18624
rect 35268 18584 35440 18612
rect 35434 18572 35440 18584
rect 35492 18572 35498 18624
rect 36078 18572 36084 18624
rect 36136 18612 36142 18624
rect 36725 18615 36783 18621
rect 36725 18612 36737 18615
rect 36136 18584 36737 18612
rect 36136 18572 36142 18584
rect 36725 18581 36737 18584
rect 36771 18581 36783 18615
rect 36725 18575 36783 18581
rect 37918 18572 37924 18624
rect 37976 18612 37982 18624
rect 38657 18615 38715 18621
rect 38657 18612 38669 18615
rect 37976 18584 38669 18612
rect 37976 18572 37982 18584
rect 38657 18581 38669 18584
rect 38703 18581 38715 18615
rect 38657 18575 38715 18581
rect 40218 18572 40224 18624
rect 40276 18612 40282 18624
rect 40313 18615 40371 18621
rect 40313 18612 40325 18615
rect 40276 18584 40325 18612
rect 40276 18572 40282 18584
rect 40313 18581 40325 18584
rect 40359 18581 40371 18615
rect 40313 18575 40371 18581
rect 1104 18522 42504 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 42504 18522
rect 1104 18448 42504 18470
rect 8297 18411 8355 18417
rect 8297 18377 8309 18411
rect 8343 18408 8355 18411
rect 8386 18408 8392 18420
rect 8343 18380 8392 18408
rect 8343 18377 8355 18380
rect 8297 18371 8355 18377
rect 8386 18368 8392 18380
rect 8444 18368 8450 18420
rect 10134 18368 10140 18420
rect 10192 18368 10198 18420
rect 11057 18411 11115 18417
rect 11057 18377 11069 18411
rect 11103 18408 11115 18411
rect 11606 18408 11612 18420
rect 11103 18380 11612 18408
rect 11103 18377 11115 18380
rect 11057 18371 11115 18377
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 17129 18411 17187 18417
rect 17129 18377 17141 18411
rect 17175 18408 17187 18411
rect 19889 18411 19947 18417
rect 17175 18380 19748 18408
rect 17175 18377 17187 18380
rect 17129 18371 17187 18377
rect 9858 18300 9864 18352
rect 9916 18300 9922 18352
rect 10152 18340 10180 18368
rect 12526 18340 12532 18352
rect 10152 18312 10916 18340
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18272 7895 18275
rect 8478 18272 8484 18284
rect 7883 18244 8484 18272
rect 7883 18241 7895 18244
rect 7837 18235 7895 18241
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 9214 18232 9220 18284
rect 9272 18232 9278 18284
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9674 18272 9680 18284
rect 9631 18244 9680 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 10042 18232 10048 18284
rect 10100 18232 10106 18284
rect 10137 18275 10195 18281
rect 10137 18241 10149 18275
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 8021 18207 8079 18213
rect 8021 18173 8033 18207
rect 8067 18204 8079 18207
rect 8846 18204 8852 18216
rect 8067 18176 8852 18204
rect 8067 18173 8079 18176
rect 8021 18167 8079 18173
rect 8846 18164 8852 18176
rect 8904 18204 8910 18216
rect 9125 18207 9183 18213
rect 9125 18204 9137 18207
rect 8904 18176 9137 18204
rect 8904 18164 8910 18176
rect 9125 18173 9137 18176
rect 9171 18173 9183 18207
rect 9692 18204 9720 18232
rect 10152 18204 10180 18235
rect 10594 18232 10600 18284
rect 10652 18232 10658 18284
rect 10888 18281 10916 18312
rect 12084 18312 12532 18340
rect 12084 18281 12112 18312
rect 12526 18300 12532 18312
rect 12584 18300 12590 18352
rect 14182 18300 14188 18352
rect 14240 18349 14246 18352
rect 14240 18340 14252 18349
rect 14240 18312 14285 18340
rect 14240 18303 14252 18312
rect 14240 18300 14246 18303
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 19720 18340 19748 18380
rect 19889 18377 19901 18411
rect 19935 18408 19947 18411
rect 19978 18408 19984 18420
rect 19935 18380 19984 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20806 18368 20812 18420
rect 20864 18408 20870 18420
rect 21453 18411 21511 18417
rect 21453 18408 21465 18411
rect 20864 18380 21465 18408
rect 20864 18368 20870 18380
rect 21453 18377 21465 18380
rect 21499 18377 21511 18411
rect 21453 18371 21511 18377
rect 26326 18368 26332 18420
rect 26384 18368 26390 18420
rect 31938 18408 31944 18420
rect 28092 18380 31944 18408
rect 20346 18340 20352 18352
rect 18472 18312 18906 18340
rect 19720 18312 20352 18340
rect 18472 18300 18478 18312
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 25038 18300 25044 18352
rect 25096 18340 25102 18352
rect 28092 18349 28120 18380
rect 31938 18368 31944 18380
rect 31996 18368 32002 18420
rect 33134 18368 33140 18420
rect 33192 18408 33198 18420
rect 33413 18411 33471 18417
rect 33413 18408 33425 18411
rect 33192 18380 33425 18408
rect 33192 18368 33198 18380
rect 33413 18377 33425 18380
rect 33459 18377 33471 18411
rect 33413 18371 33471 18377
rect 33594 18368 33600 18420
rect 33652 18408 33658 18420
rect 33781 18411 33839 18417
rect 33781 18408 33793 18411
rect 33652 18380 33793 18408
rect 33652 18368 33658 18380
rect 33781 18377 33793 18380
rect 33827 18377 33839 18411
rect 33781 18371 33839 18377
rect 35342 18368 35348 18420
rect 35400 18408 35406 18420
rect 35805 18411 35863 18417
rect 35805 18408 35817 18411
rect 35400 18380 35817 18408
rect 35400 18368 35406 18380
rect 35805 18377 35817 18380
rect 35851 18377 35863 18411
rect 35805 18371 35863 18377
rect 36173 18411 36231 18417
rect 36173 18377 36185 18411
rect 36219 18408 36231 18411
rect 36354 18408 36360 18420
rect 36219 18380 36360 18408
rect 36219 18377 36231 18380
rect 36173 18371 36231 18377
rect 36354 18368 36360 18380
rect 36412 18368 36418 18420
rect 38654 18368 38660 18420
rect 38712 18408 38718 18420
rect 38712 18380 40356 18408
rect 38712 18368 38718 18380
rect 27709 18343 27767 18349
rect 27709 18340 27721 18343
rect 25096 18312 27721 18340
rect 25096 18300 25102 18312
rect 27709 18309 27721 18312
rect 27755 18309 27767 18343
rect 27709 18303 27767 18309
rect 28077 18343 28135 18349
rect 28077 18309 28089 18343
rect 28123 18309 28135 18343
rect 28077 18303 28135 18309
rect 29086 18300 29092 18352
rect 29144 18340 29150 18352
rect 29144 18312 29486 18340
rect 29144 18300 29150 18312
rect 32582 18300 32588 18352
rect 32640 18340 32646 18352
rect 32861 18343 32919 18349
rect 32861 18340 32873 18343
rect 32640 18312 32873 18340
rect 32640 18300 32646 18312
rect 32861 18309 32873 18312
rect 32907 18309 32919 18343
rect 32861 18303 32919 18309
rect 36265 18343 36323 18349
rect 36265 18309 36277 18343
rect 36311 18340 36323 18343
rect 37918 18340 37924 18352
rect 36311 18312 37924 18340
rect 36311 18309 36323 18312
rect 36265 18303 36323 18309
rect 37918 18300 37924 18312
rect 37976 18300 37982 18352
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18241 12127 18275
rect 12069 18235 12127 18241
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18272 12495 18275
rect 13170 18272 13176 18284
rect 12483 18244 13176 18272
rect 12483 18241 12495 18244
rect 12437 18235 12495 18241
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 14366 18232 14372 18284
rect 14424 18272 14430 18284
rect 14461 18275 14519 18281
rect 14461 18272 14473 18275
rect 14424 18244 14473 18272
rect 14424 18232 14430 18244
rect 14461 18241 14473 18244
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 17034 18232 17040 18284
rect 17092 18232 17098 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18141 18275 18199 18281
rect 18141 18272 18153 18275
rect 18012 18244 18153 18272
rect 18012 18232 18018 18244
rect 18141 18241 18153 18244
rect 18187 18241 18199 18275
rect 18141 18235 18199 18241
rect 19702 18232 19708 18284
rect 19760 18272 19766 18284
rect 21361 18275 21419 18281
rect 21361 18272 21373 18275
rect 19760 18244 21373 18272
rect 19760 18232 19766 18244
rect 21361 18241 21373 18244
rect 21407 18241 21419 18275
rect 21361 18235 21419 18241
rect 26237 18275 26295 18281
rect 26237 18241 26249 18275
rect 26283 18272 26295 18275
rect 26973 18275 27031 18281
rect 26973 18272 26985 18275
rect 26283 18244 26985 18272
rect 26283 18241 26295 18244
rect 26237 18235 26295 18241
rect 26973 18241 26985 18244
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 28626 18232 28632 18284
rect 28684 18272 28690 18284
rect 28721 18275 28779 18281
rect 28721 18272 28733 18275
rect 28684 18244 28733 18272
rect 28684 18232 28690 18244
rect 28721 18241 28733 18244
rect 28767 18241 28779 18275
rect 28721 18235 28779 18241
rect 31570 18232 31576 18284
rect 31628 18272 31634 18284
rect 31665 18275 31723 18281
rect 31665 18272 31677 18275
rect 31628 18244 31677 18272
rect 31628 18232 31634 18244
rect 31665 18241 31677 18244
rect 31711 18241 31723 18275
rect 31665 18235 31723 18241
rect 32125 18275 32183 18281
rect 32125 18241 32137 18275
rect 32171 18272 32183 18275
rect 32398 18272 32404 18284
rect 32171 18244 32404 18272
rect 32171 18241 32183 18244
rect 32125 18235 32183 18241
rect 32398 18232 32404 18244
rect 32456 18232 32462 18284
rect 33873 18275 33931 18281
rect 33873 18241 33885 18275
rect 33919 18272 33931 18275
rect 34514 18272 34520 18284
rect 33919 18244 34520 18272
rect 33919 18241 33931 18244
rect 33873 18235 33931 18241
rect 34514 18232 34520 18244
rect 34572 18232 34578 18284
rect 38948 18258 38976 18380
rect 40129 18343 40187 18349
rect 40129 18309 40141 18343
rect 40175 18340 40187 18343
rect 40218 18340 40224 18352
rect 40175 18312 40224 18340
rect 40175 18309 40187 18312
rect 40129 18303 40187 18309
rect 40218 18300 40224 18312
rect 40276 18300 40282 18352
rect 40328 18340 40356 18380
rect 41046 18368 41052 18420
rect 41104 18408 41110 18420
rect 41601 18411 41659 18417
rect 41601 18408 41613 18411
rect 41104 18380 41613 18408
rect 41104 18368 41110 18380
rect 41601 18377 41613 18380
rect 41647 18377 41659 18411
rect 41601 18371 41659 18377
rect 40328 18312 40618 18340
rect 42058 18300 42064 18352
rect 42116 18340 42122 18352
rect 42153 18343 42211 18349
rect 42153 18340 42165 18343
rect 42116 18312 42165 18340
rect 42116 18300 42122 18312
rect 42153 18309 42165 18312
rect 42199 18340 42211 18343
rect 42242 18340 42248 18352
rect 42199 18312 42248 18340
rect 42199 18309 42211 18312
rect 42153 18303 42211 18309
rect 42242 18300 42248 18312
rect 42300 18300 42306 18352
rect 9692 18176 10180 18204
rect 10689 18207 10747 18213
rect 9125 18167 9183 18173
rect 10689 18173 10701 18207
rect 10735 18173 10747 18207
rect 10689 18167 10747 18173
rect 6362 18096 6368 18148
rect 6420 18136 6426 18148
rect 8110 18136 8116 18148
rect 6420 18108 8116 18136
rect 6420 18096 6426 18108
rect 8110 18096 8116 18108
rect 8168 18136 8174 18148
rect 10321 18139 10379 18145
rect 8168 18108 9904 18136
rect 8168 18096 8174 18108
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 7374 18068 7380 18080
rect 4856 18040 7380 18068
rect 4856 18028 4862 18040
rect 7374 18028 7380 18040
rect 7432 18068 7438 18080
rect 9600 18077 9628 18108
rect 7653 18071 7711 18077
rect 7653 18068 7665 18071
rect 7432 18040 7665 18068
rect 7432 18028 7438 18040
rect 7653 18037 7665 18040
rect 7699 18037 7711 18071
rect 7653 18031 7711 18037
rect 9585 18071 9643 18077
rect 9585 18037 9597 18071
rect 9631 18037 9643 18071
rect 9585 18031 9643 18037
rect 9766 18028 9772 18080
rect 9824 18028 9830 18080
rect 9876 18077 9904 18108
rect 10321 18105 10333 18139
rect 10367 18136 10379 18139
rect 10704 18136 10732 18167
rect 12526 18164 12532 18216
rect 12584 18204 12590 18216
rect 12802 18204 12808 18216
rect 12584 18176 12808 18204
rect 12584 18164 12590 18176
rect 12802 18164 12808 18176
rect 12860 18204 12866 18216
rect 17313 18207 17371 18213
rect 12860 18176 13124 18204
rect 12860 18164 12866 18176
rect 13096 18145 13124 18176
rect 17313 18173 17325 18207
rect 17359 18204 17371 18207
rect 17402 18204 17408 18216
rect 17359 18176 17408 18204
rect 17359 18173 17371 18176
rect 17313 18167 17371 18173
rect 17402 18164 17408 18176
rect 17460 18164 17466 18216
rect 18414 18164 18420 18216
rect 18472 18164 18478 18216
rect 22186 18164 22192 18216
rect 22244 18204 22250 18216
rect 22373 18207 22431 18213
rect 22373 18204 22385 18207
rect 22244 18176 22385 18204
rect 22244 18164 22250 18176
rect 22373 18173 22385 18176
rect 22419 18173 22431 18207
rect 22373 18167 22431 18173
rect 24302 18164 24308 18216
rect 24360 18204 24366 18216
rect 24946 18204 24952 18216
rect 24360 18176 24952 18204
rect 24360 18164 24366 18176
rect 24946 18164 24952 18176
rect 25004 18204 25010 18216
rect 26421 18207 26479 18213
rect 26421 18204 26433 18207
rect 25004 18176 26433 18204
rect 25004 18164 25010 18176
rect 26421 18173 26433 18176
rect 26467 18173 26479 18207
rect 26421 18167 26479 18173
rect 27522 18164 27528 18216
rect 27580 18164 27586 18216
rect 28994 18164 29000 18216
rect 29052 18164 29058 18216
rect 31018 18164 31024 18216
rect 31076 18204 31082 18216
rect 34057 18207 34115 18213
rect 34057 18204 34069 18207
rect 31076 18176 34069 18204
rect 31076 18164 31082 18176
rect 34057 18173 34069 18176
rect 34103 18204 34115 18207
rect 36446 18204 36452 18216
rect 34103 18176 36452 18204
rect 34103 18173 34115 18176
rect 34057 18167 34115 18173
rect 36446 18164 36452 18176
rect 36504 18164 36510 18216
rect 37458 18164 37464 18216
rect 37516 18204 37522 18216
rect 37553 18207 37611 18213
rect 37553 18204 37565 18207
rect 37516 18176 37565 18204
rect 37516 18164 37522 18176
rect 37553 18173 37565 18176
rect 37599 18173 37611 18207
rect 37553 18167 37611 18173
rect 11885 18139 11943 18145
rect 11885 18136 11897 18139
rect 10367 18108 10732 18136
rect 10888 18108 11897 18136
rect 10367 18105 10379 18108
rect 10321 18099 10379 18105
rect 10888 18077 10916 18108
rect 11885 18105 11897 18108
rect 11931 18105 11943 18139
rect 11885 18099 11943 18105
rect 13081 18139 13139 18145
rect 13081 18105 13093 18139
rect 13127 18105 13139 18139
rect 13081 18099 13139 18105
rect 20898 18096 20904 18148
rect 20956 18136 20962 18148
rect 21821 18139 21879 18145
rect 21821 18136 21833 18139
rect 20956 18108 21833 18136
rect 20956 18096 20962 18108
rect 21821 18105 21833 18108
rect 21867 18105 21879 18139
rect 21821 18099 21879 18105
rect 34790 18096 34796 18148
rect 34848 18136 34854 18148
rect 35986 18136 35992 18148
rect 34848 18108 35992 18136
rect 34848 18096 34854 18108
rect 35986 18096 35992 18108
rect 36044 18096 36050 18148
rect 9861 18071 9919 18077
rect 9861 18037 9873 18071
rect 9907 18037 9919 18071
rect 9861 18031 9919 18037
rect 10873 18071 10931 18077
rect 10873 18037 10885 18071
rect 10919 18037 10931 18071
rect 10873 18031 10931 18037
rect 12161 18071 12219 18077
rect 12161 18037 12173 18071
rect 12207 18068 12219 18071
rect 12802 18068 12808 18080
rect 12207 18040 12808 18068
rect 12207 18037 12219 18040
rect 12161 18031 12219 18037
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 16666 18028 16672 18080
rect 16724 18028 16730 18080
rect 25498 18028 25504 18080
rect 25556 18068 25562 18080
rect 25869 18071 25927 18077
rect 25869 18068 25881 18071
rect 25556 18040 25881 18068
rect 25556 18028 25562 18040
rect 25869 18037 25881 18040
rect 25915 18037 25927 18071
rect 25869 18031 25927 18037
rect 30466 18028 30472 18080
rect 30524 18028 30530 18080
rect 30742 18028 30748 18080
rect 30800 18068 30806 18080
rect 31389 18071 31447 18077
rect 31389 18068 31401 18071
rect 30800 18040 31401 18068
rect 30800 18028 30806 18040
rect 31389 18037 31401 18040
rect 31435 18037 31447 18071
rect 31389 18031 31447 18037
rect 35526 18028 35532 18080
rect 35584 18068 35590 18080
rect 36354 18068 36360 18080
rect 35584 18040 36360 18068
rect 35584 18028 35590 18040
rect 36354 18028 36360 18040
rect 36412 18068 36418 18080
rect 37182 18068 37188 18080
rect 36412 18040 37188 18068
rect 36412 18028 36418 18040
rect 37182 18028 37188 18040
rect 37240 18028 37246 18080
rect 37568 18068 37596 18167
rect 37826 18164 37832 18216
rect 37884 18164 37890 18216
rect 39853 18207 39911 18213
rect 39853 18204 39865 18207
rect 38856 18176 39865 18204
rect 38856 18068 38884 18176
rect 39853 18173 39865 18176
rect 39899 18173 39911 18207
rect 39853 18167 39911 18173
rect 41322 18164 41328 18216
rect 41380 18204 41386 18216
rect 41380 18176 41828 18204
rect 41380 18164 41386 18176
rect 41800 18145 41828 18176
rect 41785 18139 41843 18145
rect 41785 18105 41797 18139
rect 41831 18105 41843 18139
rect 41785 18099 41843 18105
rect 37568 18040 38884 18068
rect 39298 18028 39304 18080
rect 39356 18068 39362 18080
rect 41414 18068 41420 18080
rect 39356 18040 41420 18068
rect 39356 18028 39362 18040
rect 41414 18028 41420 18040
rect 41472 18028 41478 18080
rect 41690 18028 41696 18080
rect 41748 18028 41754 18080
rect 1104 17978 42504 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 42504 17978
rect 1104 17904 42504 17926
rect 5721 17867 5779 17873
rect 5721 17833 5733 17867
rect 5767 17864 5779 17867
rect 5810 17864 5816 17876
rect 5767 17836 5816 17864
rect 5767 17833 5779 17836
rect 5721 17827 5779 17833
rect 5810 17824 5816 17836
rect 5868 17824 5874 17876
rect 10321 17867 10379 17873
rect 10321 17833 10333 17867
rect 10367 17864 10379 17867
rect 10413 17867 10471 17873
rect 10413 17864 10425 17867
rect 10367 17836 10425 17864
rect 10367 17833 10379 17836
rect 10321 17827 10379 17833
rect 10413 17833 10425 17836
rect 10459 17833 10471 17867
rect 10413 17827 10471 17833
rect 10870 17824 10876 17876
rect 10928 17824 10934 17876
rect 18414 17824 18420 17876
rect 18472 17864 18478 17876
rect 19245 17867 19303 17873
rect 19245 17864 19257 17867
rect 18472 17836 19257 17864
rect 18472 17824 18478 17836
rect 19245 17833 19257 17836
rect 19291 17833 19303 17867
rect 19245 17827 19303 17833
rect 23750 17824 23756 17876
rect 23808 17864 23814 17876
rect 24394 17864 24400 17876
rect 23808 17836 24400 17864
rect 23808 17824 23814 17836
rect 24394 17824 24400 17836
rect 24452 17824 24458 17876
rect 26510 17824 26516 17876
rect 26568 17864 26574 17876
rect 26973 17867 27031 17873
rect 26973 17864 26985 17867
rect 26568 17836 26985 17864
rect 26568 17824 26574 17836
rect 26973 17833 26985 17836
rect 27019 17864 27031 17867
rect 27522 17864 27528 17876
rect 27019 17836 27528 17864
rect 27019 17833 27031 17836
rect 26973 17827 27031 17833
rect 27522 17824 27528 17836
rect 27580 17824 27586 17876
rect 35434 17824 35440 17876
rect 35492 17864 35498 17876
rect 35713 17867 35771 17873
rect 35713 17864 35725 17867
rect 35492 17836 35725 17864
rect 35492 17824 35498 17836
rect 35713 17833 35725 17836
rect 35759 17833 35771 17867
rect 35713 17827 35771 17833
rect 41598 17824 41604 17876
rect 41656 17824 41662 17876
rect 4614 17756 4620 17808
rect 4672 17796 4678 17808
rect 5166 17796 5172 17808
rect 4672 17768 5172 17796
rect 4672 17756 4678 17768
rect 5166 17756 5172 17768
rect 5224 17796 5230 17808
rect 5902 17796 5908 17808
rect 5224 17768 5908 17796
rect 5224 17756 5230 17768
rect 5902 17756 5908 17768
rect 5960 17756 5966 17808
rect 5994 17756 6000 17808
rect 6052 17796 6058 17808
rect 14093 17799 14151 17805
rect 14093 17796 14105 17799
rect 6052 17768 6408 17796
rect 6052 17756 6058 17768
rect 1578 17688 1584 17740
rect 1636 17728 1642 17740
rect 1765 17731 1823 17737
rect 1765 17728 1777 17731
rect 1636 17700 1777 17728
rect 1636 17688 1642 17700
rect 1765 17697 1777 17700
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17728 4951 17731
rect 5442 17728 5448 17740
rect 4939 17700 5448 17728
rect 4939 17697 4951 17700
rect 4893 17691 4951 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 6089 17731 6147 17737
rect 6089 17728 6101 17731
rect 5592 17700 6101 17728
rect 5592 17688 5598 17700
rect 6089 17697 6101 17700
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17660 1455 17663
rect 1670 17660 1676 17672
rect 1443 17632 1676 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 3191 17663 3249 17669
rect 3191 17629 3203 17663
rect 3237 17660 3249 17663
rect 4341 17663 4399 17669
rect 4341 17660 4353 17663
rect 3237 17632 4353 17660
rect 3237 17629 3249 17632
rect 3191 17623 3249 17629
rect 4341 17629 4353 17632
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 4706 17620 4712 17672
rect 4764 17660 4770 17672
rect 5077 17663 5135 17669
rect 5077 17660 5089 17663
rect 4764 17632 5089 17660
rect 4764 17620 4770 17632
rect 5077 17629 5089 17632
rect 5123 17629 5135 17663
rect 5077 17623 5135 17629
rect 5166 17620 5172 17672
rect 5224 17620 5230 17672
rect 5905 17663 5963 17669
rect 5905 17660 5917 17663
rect 5276 17632 5917 17660
rect 2774 17552 2780 17604
rect 2832 17552 2838 17604
rect 4798 17552 4804 17604
rect 4856 17592 4862 17604
rect 5276 17601 5304 17632
rect 5905 17629 5917 17632
rect 5951 17629 5963 17663
rect 5905 17623 5963 17629
rect 5261 17595 5319 17601
rect 5261 17592 5273 17595
rect 4856 17564 5273 17592
rect 4856 17552 4862 17564
rect 5261 17561 5273 17564
rect 5307 17561 5319 17595
rect 5261 17555 5319 17561
rect 5629 17595 5687 17601
rect 5629 17561 5641 17595
rect 5675 17561 5687 17595
rect 5920 17592 5948 17623
rect 5994 17620 6000 17672
rect 6052 17620 6058 17672
rect 6178 17620 6184 17672
rect 6236 17620 6242 17672
rect 6380 17669 6408 17768
rect 13924 17768 14105 17796
rect 10226 17688 10232 17740
rect 10284 17688 10290 17740
rect 12526 17688 12532 17740
rect 12584 17688 12590 17740
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 13924 17737 13952 17768
rect 14093 17765 14105 17768
rect 14139 17765 14151 17799
rect 14093 17759 14151 17765
rect 16945 17799 17003 17805
rect 16945 17765 16957 17799
rect 16991 17796 17003 17799
rect 16991 17768 18460 17796
rect 16991 17765 17003 17768
rect 16945 17759 17003 17765
rect 13909 17731 13967 17737
rect 13909 17728 13921 17731
rect 12860 17700 13921 17728
rect 12860 17688 12866 17700
rect 13909 17697 13921 17700
rect 13955 17697 13967 17731
rect 13909 17691 13967 17697
rect 17034 17688 17040 17740
rect 17092 17728 17098 17740
rect 17497 17731 17555 17737
rect 17497 17728 17509 17731
rect 17092 17700 17509 17728
rect 17092 17688 17098 17700
rect 17497 17697 17509 17700
rect 17543 17697 17555 17731
rect 17497 17691 17555 17697
rect 6365 17663 6423 17669
rect 6365 17629 6377 17663
rect 6411 17629 6423 17663
rect 6365 17623 6423 17629
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17660 7159 17663
rect 7650 17660 7656 17672
rect 7147 17632 7656 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10134 17660 10140 17672
rect 10091 17632 10140 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10502 17620 10508 17672
rect 10560 17660 10566 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 10560 17632 10609 17660
rect 10560 17620 10566 17632
rect 10597 17629 10609 17632
rect 10643 17629 10655 17663
rect 10597 17623 10655 17629
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17660 11023 17663
rect 11011 17632 12204 17660
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 6546 17592 6552 17604
rect 5920 17564 6552 17592
rect 5629 17555 5687 17561
rect 3050 17484 3056 17536
rect 3108 17524 3114 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 3108 17496 3801 17524
rect 3108 17484 3114 17496
rect 3789 17493 3801 17496
rect 3835 17493 3847 17527
rect 5644 17524 5672 17555
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 7368 17595 7426 17601
rect 7368 17561 7380 17595
rect 7414 17592 7426 17595
rect 7466 17592 7472 17604
rect 7414 17564 7472 17592
rect 7414 17561 7426 17564
rect 7368 17555 7426 17561
rect 7466 17552 7472 17564
rect 7524 17552 7530 17604
rect 9766 17552 9772 17604
rect 9824 17592 9830 17604
rect 10321 17595 10379 17601
rect 10321 17592 10333 17595
rect 9824 17564 10333 17592
rect 9824 17552 9830 17564
rect 10321 17561 10333 17564
rect 10367 17561 10379 17595
rect 10321 17555 10379 17561
rect 6086 17524 6092 17536
rect 5644 17496 6092 17524
rect 3789 17487 3847 17493
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 8481 17527 8539 17533
rect 8481 17493 8493 17527
rect 8527 17524 8539 17527
rect 8846 17524 8852 17536
rect 8527 17496 8852 17524
rect 8527 17493 8539 17496
rect 8481 17487 8539 17493
rect 8846 17484 8852 17496
rect 8904 17524 8910 17536
rect 9398 17524 9404 17536
rect 8904 17496 9404 17524
rect 8904 17484 8910 17496
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 9858 17484 9864 17536
rect 9916 17484 9922 17536
rect 12176 17533 12204 17632
rect 15470 17620 15476 17672
rect 15528 17660 15534 17672
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 15528 17632 15577 17660
rect 15528 17620 15534 17632
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 15832 17663 15890 17669
rect 15832 17629 15844 17663
rect 15878 17660 15890 17663
rect 16666 17660 16672 17672
rect 15878 17632 16672 17660
rect 15878 17629 15890 17632
rect 15832 17623 15890 17629
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 17512 17660 17540 17691
rect 17678 17688 17684 17740
rect 17736 17728 17742 17740
rect 18322 17728 18328 17740
rect 17736 17700 18328 17728
rect 17736 17688 17742 17700
rect 18322 17688 18328 17700
rect 18380 17688 18386 17740
rect 18432 17737 18460 17768
rect 22002 17756 22008 17808
rect 22060 17796 22066 17808
rect 22373 17799 22431 17805
rect 22373 17796 22385 17799
rect 22060 17768 22385 17796
rect 22060 17756 22066 17768
rect 22373 17765 22385 17768
rect 22419 17765 22431 17799
rect 33318 17796 33324 17808
rect 22373 17759 22431 17765
rect 32324 17768 33324 17796
rect 18417 17731 18475 17737
rect 18417 17697 18429 17731
rect 18463 17697 18475 17731
rect 18417 17691 18475 17697
rect 19702 17688 19708 17740
rect 19760 17728 19766 17740
rect 19797 17731 19855 17737
rect 19797 17728 19809 17731
rect 19760 17700 19809 17728
rect 19760 17688 19766 17700
rect 19797 17697 19809 17700
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 19886 17688 19892 17740
rect 19944 17728 19950 17740
rect 20625 17731 20683 17737
rect 20625 17728 20637 17731
rect 19944 17700 20637 17728
rect 19944 17688 19950 17700
rect 20625 17697 20637 17700
rect 20671 17728 20683 17731
rect 24213 17731 24271 17737
rect 20671 17700 22508 17728
rect 20671 17697 20683 17700
rect 20625 17691 20683 17697
rect 22480 17672 22508 17700
rect 24213 17697 24225 17731
rect 24259 17728 24271 17731
rect 24946 17728 24952 17740
rect 24259 17700 24952 17728
rect 24259 17697 24271 17700
rect 24213 17691 24271 17697
rect 24946 17688 24952 17700
rect 25004 17688 25010 17740
rect 25222 17688 25228 17740
rect 25280 17688 25286 17740
rect 25498 17688 25504 17740
rect 25556 17688 25562 17740
rect 30190 17728 30196 17740
rect 29380 17700 30196 17728
rect 17865 17663 17923 17669
rect 17865 17660 17877 17663
rect 17512 17632 17877 17660
rect 17865 17629 17877 17632
rect 17911 17629 17923 17663
rect 17865 17623 17923 17629
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19978 17660 19984 17672
rect 19659 17632 19984 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 22462 17620 22468 17672
rect 22520 17620 22526 17672
rect 29380 17669 29408 17700
rect 30190 17688 30196 17700
rect 30248 17728 30254 17740
rect 30837 17731 30895 17737
rect 30248 17700 30788 17728
rect 30248 17688 30254 17700
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 29181 17663 29239 17669
rect 29181 17629 29193 17663
rect 29227 17629 29239 17663
rect 29181 17623 29239 17629
rect 29365 17663 29423 17669
rect 29365 17629 29377 17663
rect 29411 17629 29423 17663
rect 29365 17623 29423 17629
rect 30285 17663 30343 17669
rect 30285 17629 30297 17663
rect 30331 17660 30343 17663
rect 30466 17660 30472 17672
rect 30331 17632 30472 17660
rect 30331 17629 30343 17632
rect 30285 17623 30343 17629
rect 12342 17601 12348 17604
rect 12320 17595 12348 17601
rect 12320 17561 12332 17595
rect 12320 17555 12348 17561
rect 12342 17552 12348 17555
rect 12400 17552 12406 17604
rect 13906 17552 13912 17604
rect 13964 17592 13970 17604
rect 15206 17595 15264 17601
rect 15206 17592 15218 17595
rect 13964 17564 15218 17592
rect 13964 17552 13970 17564
rect 15206 17561 15218 17564
rect 15252 17561 15264 17595
rect 15206 17555 15264 17561
rect 20898 17552 20904 17604
rect 20956 17552 20962 17604
rect 22126 17564 22692 17592
rect 12161 17527 12219 17533
rect 12161 17493 12173 17527
rect 12207 17493 12219 17527
rect 12161 17487 12219 17493
rect 12437 17527 12495 17533
rect 12437 17493 12449 17527
rect 12483 17524 12495 17527
rect 12710 17524 12716 17536
rect 12483 17496 12716 17524
rect 12483 17493 12495 17496
rect 12437 17487 12495 17493
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 13265 17527 13323 17533
rect 13265 17493 13277 17527
rect 13311 17524 13323 17527
rect 13538 17524 13544 17536
rect 13311 17496 13544 17524
rect 13311 17493 13323 17496
rect 13265 17487 13323 17493
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 17034 17484 17040 17536
rect 17092 17484 17098 17536
rect 17402 17484 17408 17536
rect 17460 17484 17466 17536
rect 19702 17484 19708 17536
rect 19760 17484 19766 17536
rect 22664 17524 22692 17564
rect 22738 17552 22744 17604
rect 22796 17552 22802 17604
rect 25038 17592 25044 17604
rect 23966 17564 25044 17592
rect 24044 17524 24072 17564
rect 25038 17552 25044 17564
rect 25096 17592 25102 17604
rect 27080 17592 27108 17623
rect 25096 17564 25990 17592
rect 27080 17564 27200 17592
rect 25096 17552 25102 17564
rect 22664 17496 24072 17524
rect 27172 17524 27200 17564
rect 27338 17552 27344 17604
rect 27396 17552 27402 17604
rect 29086 17592 29092 17604
rect 28566 17564 29092 17592
rect 29086 17552 29092 17564
rect 29144 17552 29150 17604
rect 29196 17592 29224 17623
rect 30300 17592 30328 17623
rect 30466 17620 30472 17632
rect 30524 17660 30530 17672
rect 30760 17669 30788 17700
rect 30837 17697 30849 17731
rect 30883 17728 30895 17731
rect 31754 17728 31760 17740
rect 30883 17700 31760 17728
rect 30883 17697 30895 17700
rect 30837 17691 30895 17697
rect 31754 17688 31760 17700
rect 31812 17688 31818 17740
rect 30561 17663 30619 17669
rect 30561 17660 30573 17663
rect 30524 17632 30573 17660
rect 30524 17620 30530 17632
rect 30561 17629 30573 17632
rect 30607 17629 30619 17663
rect 30561 17623 30619 17629
rect 30745 17663 30803 17669
rect 30745 17629 30757 17663
rect 30791 17629 30803 17663
rect 32324 17660 32352 17768
rect 33318 17756 33324 17768
rect 33376 17756 33382 17808
rect 35066 17756 35072 17808
rect 35124 17796 35130 17808
rect 35124 17768 36571 17796
rect 35124 17756 35130 17768
rect 32585 17731 32643 17737
rect 32585 17697 32597 17731
rect 32631 17728 32643 17731
rect 33229 17731 33287 17737
rect 33229 17728 33241 17731
rect 32631 17700 33241 17728
rect 32631 17697 32643 17700
rect 32585 17691 32643 17697
rect 33229 17697 33241 17700
rect 33275 17697 33287 17731
rect 33229 17691 33287 17697
rect 36357 17731 36415 17737
rect 36357 17697 36369 17731
rect 36403 17728 36415 17731
rect 36446 17728 36452 17740
rect 36403 17700 36452 17728
rect 36403 17697 36415 17700
rect 36357 17691 36415 17697
rect 32246 17632 32352 17660
rect 33244 17660 33272 17691
rect 36446 17688 36452 17700
rect 36504 17688 36510 17740
rect 36543 17728 36571 17768
rect 39574 17756 39580 17808
rect 39632 17796 39638 17808
rect 39632 17768 42196 17796
rect 39632 17756 39638 17768
rect 39393 17731 39451 17737
rect 36543 17700 39344 17728
rect 33413 17663 33471 17669
rect 33413 17660 33425 17663
rect 33244 17632 33425 17660
rect 30745 17623 30803 17629
rect 33413 17629 33425 17632
rect 33459 17629 33471 17663
rect 33413 17623 33471 17629
rect 29196 17564 30328 17592
rect 31110 17552 31116 17604
rect 31168 17552 31174 17604
rect 32677 17595 32735 17601
rect 32677 17592 32689 17595
rect 32416 17564 32689 17592
rect 27614 17524 27620 17536
rect 27172 17496 27620 17524
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 28718 17484 28724 17536
rect 28776 17524 28782 17536
rect 28813 17527 28871 17533
rect 28813 17524 28825 17527
rect 28776 17496 28825 17524
rect 28776 17484 28782 17496
rect 28813 17493 28825 17496
rect 28859 17493 28871 17527
rect 28813 17487 28871 17493
rect 29273 17527 29331 17533
rect 29273 17493 29285 17527
rect 29319 17524 29331 17527
rect 29454 17524 29460 17536
rect 29319 17496 29460 17524
rect 29319 17493 29331 17496
rect 29273 17487 29331 17493
rect 29454 17484 29460 17496
rect 29512 17484 29518 17536
rect 29641 17527 29699 17533
rect 29641 17493 29653 17527
rect 29687 17524 29699 17527
rect 29730 17524 29736 17536
rect 29687 17496 29736 17524
rect 29687 17493 29699 17496
rect 29641 17487 29699 17493
rect 29730 17484 29736 17496
rect 29788 17484 29794 17536
rect 30190 17484 30196 17536
rect 30248 17524 30254 17536
rect 30377 17527 30435 17533
rect 30377 17524 30389 17527
rect 30248 17496 30389 17524
rect 30248 17484 30254 17496
rect 30377 17493 30389 17496
rect 30423 17493 30435 17527
rect 30377 17487 30435 17493
rect 30650 17484 30656 17536
rect 30708 17524 30714 17536
rect 32416 17524 32444 17564
rect 32677 17561 32689 17564
rect 32723 17561 32735 17595
rect 33428 17592 33456 17623
rect 33502 17620 33508 17672
rect 33560 17660 33566 17672
rect 33597 17663 33655 17669
rect 33597 17660 33609 17663
rect 33560 17632 33609 17660
rect 33560 17620 33566 17632
rect 33597 17629 33609 17632
rect 33643 17629 33655 17663
rect 33597 17623 33655 17629
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 34790 17660 34796 17672
rect 34572 17632 34796 17660
rect 34572 17620 34578 17632
rect 34790 17620 34796 17632
rect 34848 17620 34854 17672
rect 34974 17620 34980 17672
rect 35032 17660 35038 17672
rect 36541 17663 36599 17669
rect 36541 17660 36553 17663
rect 35032 17632 36553 17660
rect 35032 17620 35038 17632
rect 36541 17629 36553 17632
rect 36587 17629 36599 17663
rect 36541 17623 36599 17629
rect 36998 17620 37004 17672
rect 37056 17660 37062 17672
rect 37093 17663 37151 17669
rect 37093 17660 37105 17663
rect 37056 17632 37105 17660
rect 37056 17620 37062 17632
rect 37093 17629 37105 17632
rect 37139 17629 37151 17663
rect 37093 17623 37151 17629
rect 37458 17620 37464 17672
rect 37516 17660 37522 17672
rect 37645 17663 37703 17669
rect 37645 17660 37657 17663
rect 37516 17632 37657 17660
rect 37516 17620 37522 17632
rect 37645 17629 37657 17632
rect 37691 17629 37703 17663
rect 39316 17660 39344 17700
rect 39393 17697 39405 17731
rect 39439 17728 39451 17731
rect 39942 17728 39948 17740
rect 39439 17700 39948 17728
rect 39439 17697 39451 17700
rect 39393 17691 39451 17697
rect 39942 17688 39948 17700
rect 40000 17728 40006 17740
rect 40405 17731 40463 17737
rect 40405 17728 40417 17731
rect 40000 17700 40417 17728
rect 40000 17688 40006 17700
rect 40405 17697 40417 17700
rect 40451 17697 40463 17731
rect 40405 17691 40463 17697
rect 40957 17731 41015 17737
rect 40957 17697 40969 17731
rect 41003 17728 41015 17731
rect 41046 17728 41052 17740
rect 41003 17700 41052 17728
rect 41003 17697 41015 17700
rect 40957 17691 41015 17697
rect 41046 17688 41052 17700
rect 41104 17688 41110 17740
rect 41509 17731 41567 17737
rect 41509 17697 41521 17731
rect 41555 17728 41567 17731
rect 41555 17700 42012 17728
rect 41555 17697 41567 17700
rect 41509 17691 41567 17697
rect 39850 17660 39856 17672
rect 39316 17632 39856 17660
rect 37645 17623 37703 17629
rect 39850 17620 39856 17632
rect 39908 17620 39914 17672
rect 41414 17620 41420 17672
rect 41472 17660 41478 17672
rect 41984 17669 42012 17700
rect 42168 17669 42196 17768
rect 41785 17663 41843 17669
rect 41785 17660 41797 17663
rect 41472 17632 41797 17660
rect 41472 17620 41478 17632
rect 41785 17629 41797 17632
rect 41831 17629 41843 17663
rect 41785 17623 41843 17629
rect 41969 17663 42027 17669
rect 41969 17629 41981 17663
rect 42015 17629 42027 17663
rect 41969 17623 42027 17629
rect 42153 17663 42211 17669
rect 42153 17629 42165 17663
rect 42199 17629 42211 17663
rect 42153 17623 42211 17629
rect 33778 17592 33784 17604
rect 33428 17564 33784 17592
rect 32677 17555 32735 17561
rect 33778 17552 33784 17564
rect 33836 17552 33842 17604
rect 34698 17552 34704 17604
rect 34756 17592 34762 17604
rect 35345 17595 35403 17601
rect 35345 17592 35357 17595
rect 34756 17564 35357 17592
rect 34756 17552 34762 17564
rect 35345 17561 35357 17564
rect 35391 17561 35403 17595
rect 35345 17555 35403 17561
rect 35526 17552 35532 17604
rect 35584 17552 35590 17604
rect 36078 17552 36084 17604
rect 36136 17552 36142 17604
rect 37921 17595 37979 17601
rect 37921 17561 37933 17595
rect 37967 17592 37979 17595
rect 38010 17592 38016 17604
rect 37967 17564 38016 17592
rect 37967 17561 37979 17564
rect 37921 17555 37979 17561
rect 38010 17552 38016 17564
rect 38068 17552 38074 17604
rect 38654 17552 38660 17604
rect 38712 17552 38718 17604
rect 39868 17592 39896 17620
rect 41877 17595 41935 17601
rect 41877 17592 41889 17595
rect 39868 17564 41889 17592
rect 41877 17561 41889 17564
rect 41923 17561 41935 17595
rect 41877 17555 41935 17561
rect 30708 17496 32444 17524
rect 30708 17484 30714 17496
rect 33502 17484 33508 17536
rect 33560 17484 33566 17536
rect 34514 17484 34520 17536
rect 34572 17524 34578 17536
rect 35161 17527 35219 17533
rect 35161 17524 35173 17527
rect 34572 17496 35173 17524
rect 34572 17484 34578 17496
rect 35161 17493 35173 17496
rect 35207 17524 35219 17527
rect 35434 17524 35440 17536
rect 35207 17496 35440 17524
rect 35207 17493 35219 17496
rect 35161 17487 35219 17493
rect 35434 17484 35440 17496
rect 35492 17484 35498 17536
rect 36173 17527 36231 17533
rect 36173 17493 36185 17527
rect 36219 17524 36231 17527
rect 38838 17524 38844 17536
rect 36219 17496 38844 17524
rect 36219 17493 36231 17496
rect 36173 17487 36231 17493
rect 38838 17484 38844 17496
rect 38896 17524 38902 17536
rect 39853 17527 39911 17533
rect 39853 17524 39865 17527
rect 38896 17496 39865 17524
rect 38896 17484 38902 17496
rect 39853 17493 39865 17496
rect 39899 17493 39911 17527
rect 39853 17487 39911 17493
rect 1104 17434 42504 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 42504 17434
rect 1104 17360 42504 17382
rect 4479 17323 4537 17329
rect 4479 17289 4491 17323
rect 4525 17320 4537 17323
rect 4798 17320 4804 17332
rect 4525 17292 4804 17320
rect 4525 17289 4537 17292
rect 4479 17283 4537 17289
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 5169 17323 5227 17329
rect 5169 17289 5181 17323
rect 5215 17320 5227 17323
rect 5258 17320 5264 17332
rect 5215 17292 5264 17320
rect 5215 17289 5227 17292
rect 5169 17283 5227 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5994 17320 6000 17332
rect 5368 17292 6000 17320
rect 4982 17252 4988 17264
rect 4094 17238 4988 17252
rect 4080 17224 4988 17238
rect 842 17144 848 17196
rect 900 17184 906 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 900 17156 1409 17184
rect 900 17144 906 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 3970 17144 3976 17196
rect 4028 17184 4034 17196
rect 4080 17184 4108 17224
rect 4982 17212 4988 17224
rect 5040 17212 5046 17264
rect 5368 17252 5396 17292
rect 5994 17280 6000 17292
rect 6052 17320 6058 17332
rect 6089 17323 6147 17329
rect 6089 17320 6101 17323
rect 6052 17292 6101 17320
rect 6052 17280 6058 17292
rect 6089 17289 6101 17292
rect 6135 17289 6147 17323
rect 6089 17283 6147 17289
rect 7466 17280 7472 17332
rect 7524 17280 7530 17332
rect 10505 17323 10563 17329
rect 10505 17289 10517 17323
rect 10551 17320 10563 17323
rect 10594 17320 10600 17332
rect 10551 17292 10600 17320
rect 10551 17289 10563 17292
rect 10505 17283 10563 17289
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 12492 17292 12541 17320
rect 12492 17280 12498 17292
rect 12529 17289 12541 17292
rect 12575 17320 12587 17323
rect 12802 17320 12808 17332
rect 12575 17292 12808 17320
rect 12575 17289 12587 17292
rect 12529 17283 12587 17289
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 12989 17323 13047 17329
rect 12989 17289 13001 17323
rect 13035 17289 13047 17323
rect 12989 17283 13047 17289
rect 6917 17255 6975 17261
rect 6917 17252 6929 17255
rect 5092 17224 5396 17252
rect 5444 17224 6929 17252
rect 4028 17156 4108 17184
rect 4028 17144 4034 17156
rect 4890 17144 4896 17196
rect 4948 17144 4954 17196
rect 5092 17193 5120 17224
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5444 17184 5472 17224
rect 6917 17221 6929 17224
rect 6963 17221 6975 17255
rect 6917 17215 6975 17221
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 13004 17252 13032 17283
rect 17402 17280 17408 17332
rect 17460 17320 17466 17332
rect 17497 17323 17555 17329
rect 17497 17320 17509 17323
rect 17460 17292 17509 17320
rect 17460 17280 17466 17292
rect 17497 17289 17509 17292
rect 17543 17289 17555 17323
rect 17497 17283 17555 17289
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 25222 17320 25228 17332
rect 22520 17292 25228 17320
rect 22520 17280 22526 17292
rect 12400 17224 13032 17252
rect 12400 17212 12406 17224
rect 5316 17156 5472 17184
rect 5537 17187 5595 17193
rect 5316 17144 5322 17156
rect 5537 17153 5549 17187
rect 5583 17153 5595 17187
rect 5537 17147 5595 17153
rect 1762 17076 1768 17128
rect 1820 17116 1826 17128
rect 2685 17119 2743 17125
rect 2685 17116 2697 17119
rect 1820 17088 2697 17116
rect 1820 17076 1826 17088
rect 2685 17085 2697 17088
rect 2731 17085 2743 17119
rect 2685 17079 2743 17085
rect 5166 17076 5172 17128
rect 5224 17116 5230 17128
rect 5552 17116 5580 17147
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6086 17144 6092 17196
rect 6144 17184 6150 17196
rect 6181 17187 6239 17193
rect 6181 17184 6193 17187
rect 6144 17156 6193 17184
rect 6144 17144 6150 17156
rect 6181 17153 6193 17156
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 6546 17144 6552 17196
rect 6604 17184 6610 17196
rect 6641 17187 6699 17193
rect 6641 17184 6653 17187
rect 6604 17156 6653 17184
rect 6604 17144 6610 17156
rect 6641 17153 6653 17156
rect 6687 17153 6699 17187
rect 6641 17147 6699 17153
rect 5224 17088 5580 17116
rect 5224 17076 5230 17088
rect 5626 17076 5632 17128
rect 5684 17076 5690 17128
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17085 5871 17119
rect 5813 17079 5871 17085
rect 5828 17048 5856 17079
rect 6362 17076 6368 17128
rect 6420 17076 6426 17128
rect 6656 17116 6684 17147
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6788 17156 7205 17184
rect 6788 17144 6794 17156
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7374 17144 7380 17196
rect 7432 17144 7438 17196
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 7926 17184 7932 17196
rect 7607 17156 7932 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8110 17193 8116 17196
rect 8104 17147 8116 17193
rect 8110 17144 8116 17147
rect 8168 17144 8174 17196
rect 9398 17144 9404 17196
rect 9456 17144 9462 17196
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17184 9919 17187
rect 9950 17184 9956 17196
rect 9907 17156 9956 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6656 17088 6929 17116
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 7650 17076 7656 17128
rect 7708 17116 7714 17128
rect 7837 17119 7895 17125
rect 7837 17116 7849 17119
rect 7708 17088 7849 17116
rect 7708 17076 7714 17088
rect 7837 17085 7849 17088
rect 7883 17085 7895 17119
rect 9508 17116 9536 17147
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 10689 17187 10747 17193
rect 10689 17153 10701 17187
rect 10735 17184 10747 17187
rect 10965 17187 11023 17193
rect 10735 17156 10916 17184
rect 10735 17153 10747 17156
rect 10689 17147 10747 17153
rect 7837 17079 7895 17085
rect 9416 17088 9536 17116
rect 10781 17119 10839 17125
rect 6825 17051 6883 17057
rect 6825 17048 6837 17051
rect 5828 17020 6837 17048
rect 6825 17017 6837 17020
rect 6871 17017 6883 17051
rect 6825 17011 6883 17017
rect 9416 16992 9444 17088
rect 10781 17085 10793 17119
rect 10827 17085 10839 17119
rect 10888 17116 10916 17156
rect 10965 17153 10977 17187
rect 11011 17184 11023 17187
rect 11422 17184 11428 17196
rect 11011 17156 11428 17184
rect 11011 17153 11023 17156
rect 10965 17147 11023 17153
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 12437 17187 12495 17193
rect 12437 17153 12449 17187
rect 12483 17184 12495 17187
rect 12618 17184 12624 17196
rect 12483 17156 12624 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 11054 17116 11060 17128
rect 10888 17088 11060 17116
rect 10781 17079 10839 17085
rect 10045 17051 10103 17057
rect 10045 17017 10057 17051
rect 10091 17048 10103 17051
rect 10796 17048 10824 17079
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 12176 17116 12204 17147
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 12728 17193 12756 17224
rect 20806 17212 20812 17264
rect 20864 17212 20870 17264
rect 23750 17212 23756 17264
rect 23808 17212 23814 17264
rect 12713 17187 12771 17193
rect 12713 17153 12725 17187
rect 12759 17153 12771 17187
rect 12713 17147 12771 17153
rect 13262 17144 13268 17196
rect 13320 17184 13326 17196
rect 14102 17187 14160 17193
rect 14102 17184 14114 17187
rect 13320 17156 14114 17184
rect 13320 17144 13326 17156
rect 14102 17153 14114 17156
rect 14148 17153 14160 17187
rect 14102 17147 14160 17153
rect 19886 17144 19892 17196
rect 19944 17144 19950 17196
rect 21818 17144 21824 17196
rect 21876 17144 21882 17196
rect 22002 17144 22008 17196
rect 22060 17184 22066 17196
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 22060 17156 22385 17184
rect 22060 17144 22066 17156
rect 22373 17153 22385 17156
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17153 23719 17187
rect 23661 17147 23719 17153
rect 12526 17116 12532 17128
rect 12176 17088 12532 17116
rect 12526 17076 12532 17088
rect 12584 17116 12590 17128
rect 12802 17116 12808 17128
rect 12584 17088 12808 17116
rect 12584 17076 12590 17088
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 14366 17076 14372 17128
rect 14424 17076 14430 17128
rect 18138 17076 18144 17128
rect 18196 17076 18202 17128
rect 20165 17119 20223 17125
rect 20165 17085 20177 17119
rect 20211 17116 20223 17119
rect 20806 17116 20812 17128
rect 20211 17088 20812 17116
rect 20211 17085 20223 17088
rect 20165 17079 20223 17085
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 10091 17020 10824 17048
rect 12253 17051 12311 17057
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 12986 17048 12992 17060
rect 12299 17020 12992 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12986 17008 12992 17020
rect 13044 17008 13050 17060
rect 21637 17051 21695 17057
rect 21637 17017 21649 17051
rect 21683 17048 21695 17051
rect 22094 17048 22100 17060
rect 21683 17020 22100 17048
rect 21683 17017 21695 17020
rect 21637 17011 21695 17017
rect 22094 17008 22100 17020
rect 22152 17008 22158 17060
rect 22738 17008 22744 17060
rect 22796 17048 22802 17060
rect 23477 17051 23535 17057
rect 23477 17048 23489 17051
rect 22796 17020 23489 17048
rect 22796 17008 22802 17020
rect 23477 17017 23489 17020
rect 23523 17017 23535 17051
rect 23477 17011 23535 17017
rect 1578 16940 1584 16992
rect 1636 16940 1642 16992
rect 4614 16940 4620 16992
rect 4672 16940 4678 16992
rect 4893 16983 4951 16989
rect 4893 16949 4905 16983
rect 4939 16980 4951 16983
rect 5442 16980 5448 16992
rect 4939 16952 5448 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 5902 16940 5908 16992
rect 5960 16980 5966 16992
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 5960 16952 6469 16980
rect 5960 16940 5966 16952
rect 6457 16949 6469 16952
rect 6503 16949 6515 16983
rect 6457 16943 6515 16949
rect 6546 16940 6552 16992
rect 6604 16980 6610 16992
rect 7101 16983 7159 16989
rect 7101 16980 7113 16983
rect 6604 16952 7113 16980
rect 6604 16940 6610 16952
rect 7101 16949 7113 16952
rect 7147 16949 7159 16983
rect 7101 16943 7159 16949
rect 9214 16940 9220 16992
rect 9272 16980 9278 16992
rect 9398 16980 9404 16992
rect 9272 16952 9404 16980
rect 9272 16940 9278 16952
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 9861 16983 9919 16989
rect 9861 16949 9873 16983
rect 9907 16980 9919 16983
rect 10318 16980 10324 16992
rect 9907 16952 10324 16980
rect 9907 16949 9919 16952
rect 9861 16943 9919 16949
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10560 16952 10701 16980
rect 10560 16940 10566 16952
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10689 16943 10747 16949
rect 12894 16940 12900 16992
rect 12952 16940 12958 16992
rect 21358 16940 21364 16992
rect 21416 16980 21422 16992
rect 21913 16983 21971 16989
rect 21913 16980 21925 16983
rect 21416 16952 21925 16980
rect 21416 16940 21422 16952
rect 21913 16949 21925 16952
rect 21959 16949 21971 16983
rect 21913 16943 21971 16949
rect 22554 16940 22560 16992
rect 22612 16980 22618 16992
rect 23017 16983 23075 16989
rect 23017 16980 23029 16983
rect 22612 16952 23029 16980
rect 22612 16940 22618 16952
rect 23017 16949 23029 16952
rect 23063 16949 23075 16983
rect 23676 16980 23704 17147
rect 23842 17144 23848 17196
rect 23900 17144 23906 17196
rect 24136 17193 24164 17292
rect 25222 17280 25228 17292
rect 25280 17280 25286 17332
rect 27338 17280 27344 17332
rect 27396 17320 27402 17332
rect 27893 17323 27951 17329
rect 27893 17320 27905 17323
rect 27396 17292 27905 17320
rect 27396 17280 27402 17292
rect 27893 17289 27905 17292
rect 27939 17289 27951 17323
rect 27893 17283 27951 17289
rect 28994 17280 29000 17332
rect 29052 17320 29058 17332
rect 29365 17323 29423 17329
rect 29365 17320 29377 17323
rect 29052 17292 29377 17320
rect 29052 17280 29058 17292
rect 29365 17289 29377 17292
rect 29411 17289 29423 17323
rect 29365 17283 29423 17289
rect 30285 17323 30343 17329
rect 30285 17289 30297 17323
rect 30331 17320 30343 17323
rect 30331 17292 31064 17320
rect 30331 17289 30343 17292
rect 30285 17283 30343 17289
rect 24394 17212 24400 17264
rect 24452 17212 24458 17264
rect 25038 17212 25044 17264
rect 25096 17212 25102 17264
rect 28261 17255 28319 17261
rect 28261 17252 28273 17255
rect 25700 17224 28273 17252
rect 24029 17187 24087 17193
rect 24029 17153 24041 17187
rect 24075 17153 24087 17187
rect 24029 17147 24087 17153
rect 24121 17187 24179 17193
rect 24121 17153 24133 17187
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 24044 17116 24072 17147
rect 24486 17116 24492 17128
rect 24044 17088 24492 17116
rect 24486 17076 24492 17088
rect 24544 17116 24550 17128
rect 25700 17116 25728 17224
rect 28261 17221 28273 17224
rect 28307 17221 28319 17255
rect 28261 17215 28319 17221
rect 28399 17255 28457 17261
rect 28399 17221 28411 17255
rect 28445 17252 28457 17255
rect 28902 17252 28908 17264
rect 28445 17224 28908 17252
rect 28445 17221 28457 17224
rect 28399 17215 28457 17221
rect 28902 17212 28908 17224
rect 28960 17252 28966 17264
rect 29273 17255 29331 17261
rect 29273 17252 29285 17255
rect 28960 17224 29285 17252
rect 28960 17212 28966 17224
rect 29273 17221 29285 17224
rect 29319 17252 29331 17255
rect 29319 17224 29592 17252
rect 29319 17221 29331 17224
rect 29273 17215 29331 17221
rect 27430 17144 27436 17196
rect 27488 17144 27494 17196
rect 27617 17187 27675 17193
rect 27617 17153 27629 17187
rect 27663 17184 27675 17187
rect 27706 17184 27712 17196
rect 27663 17156 27712 17184
rect 27663 17153 27675 17156
rect 27617 17147 27675 17153
rect 27706 17144 27712 17156
rect 27764 17144 27770 17196
rect 28074 17144 28080 17196
rect 28132 17144 28138 17196
rect 28166 17144 28172 17196
rect 28224 17144 28230 17196
rect 28718 17144 28724 17196
rect 28776 17144 28782 17196
rect 29564 17193 29592 17224
rect 29730 17212 29736 17264
rect 29788 17212 29794 17264
rect 30650 17212 30656 17264
rect 30708 17212 30714 17264
rect 31036 17252 31064 17292
rect 31110 17280 31116 17332
rect 31168 17280 31174 17332
rect 34609 17323 34667 17329
rect 32968 17292 34468 17320
rect 32030 17252 32036 17264
rect 31036 17224 32036 17252
rect 32030 17212 32036 17224
rect 32088 17252 32094 17264
rect 32088 17224 32720 17252
rect 32088 17212 32094 17224
rect 29549 17187 29607 17193
rect 29549 17153 29561 17187
rect 29595 17153 29607 17187
rect 29549 17147 29607 17153
rect 29638 17144 29644 17196
rect 29696 17144 29702 17196
rect 29917 17187 29975 17193
rect 29917 17153 29929 17187
rect 29963 17153 29975 17187
rect 29917 17147 29975 17153
rect 24544 17088 25728 17116
rect 25869 17119 25927 17125
rect 24544 17076 24550 17088
rect 25869 17085 25881 17119
rect 25915 17116 25927 17119
rect 26050 17116 26056 17128
rect 25915 17088 26056 17116
rect 25915 17085 25927 17088
rect 25869 17079 25927 17085
rect 26050 17076 26056 17088
rect 26108 17116 26114 17128
rect 26513 17119 26571 17125
rect 26513 17116 26525 17119
rect 26108 17088 26525 17116
rect 26108 17076 26114 17088
rect 26513 17085 26525 17088
rect 26559 17085 26571 17119
rect 26513 17079 26571 17085
rect 28537 17119 28595 17125
rect 28537 17085 28549 17119
rect 28583 17085 28595 17119
rect 28537 17079 28595 17085
rect 25498 17008 25504 17060
rect 25556 17048 25562 17060
rect 25961 17051 26019 17057
rect 25961 17048 25973 17051
rect 25556 17020 25973 17048
rect 25556 17008 25562 17020
rect 25961 17017 25973 17020
rect 26007 17017 26019 17051
rect 28552 17048 28580 17079
rect 28994 17076 29000 17128
rect 29052 17116 29058 17128
rect 29932 17116 29960 17147
rect 30190 17144 30196 17196
rect 30248 17144 30254 17196
rect 30469 17187 30527 17193
rect 30469 17153 30481 17187
rect 30515 17184 30527 17187
rect 30558 17184 30564 17196
rect 30515 17156 30564 17184
rect 30515 17153 30527 17156
rect 30469 17147 30527 17153
rect 30558 17144 30564 17156
rect 30616 17144 30622 17196
rect 30742 17144 30748 17196
rect 30800 17144 30806 17196
rect 30837 17187 30895 17193
rect 30837 17153 30849 17187
rect 30883 17153 30895 17187
rect 30837 17147 30895 17153
rect 29052 17088 29960 17116
rect 29052 17076 29058 17088
rect 30374 17076 30380 17128
rect 30432 17116 30438 17128
rect 30852 17116 30880 17147
rect 31938 17144 31944 17196
rect 31996 17184 32002 17196
rect 32692 17193 32720 17224
rect 32968 17193 32996 17292
rect 34440 17264 34468 17292
rect 34609 17289 34621 17323
rect 34655 17289 34667 17323
rect 34609 17283 34667 17289
rect 33689 17255 33747 17261
rect 33689 17252 33701 17255
rect 33060 17224 33701 17252
rect 32125 17187 32183 17193
rect 32125 17184 32137 17187
rect 31996 17156 32137 17184
rect 31996 17144 32002 17156
rect 32125 17153 32137 17156
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 32677 17187 32735 17193
rect 32677 17153 32689 17187
rect 32723 17153 32735 17187
rect 32677 17147 32735 17153
rect 32953 17187 33011 17193
rect 32953 17153 32965 17187
rect 32999 17153 33011 17187
rect 32953 17147 33011 17153
rect 30432 17088 30880 17116
rect 31665 17119 31723 17125
rect 30432 17076 30438 17088
rect 31665 17085 31677 17119
rect 31711 17085 31723 17119
rect 31665 17079 31723 17085
rect 32769 17119 32827 17125
rect 32769 17085 32781 17119
rect 32815 17116 32827 17119
rect 33060 17116 33088 17224
rect 33244 17196 33272 17224
rect 33689 17221 33701 17224
rect 33735 17221 33747 17255
rect 33689 17215 33747 17221
rect 34422 17212 34428 17264
rect 34480 17212 34486 17264
rect 34624 17252 34652 17283
rect 37826 17280 37832 17332
rect 37884 17320 37890 17332
rect 37921 17323 37979 17329
rect 37921 17320 37933 17323
rect 37884 17292 37933 17320
rect 37884 17280 37890 17292
rect 37921 17289 37933 17292
rect 37967 17289 37979 17323
rect 37921 17283 37979 17289
rect 38010 17280 38016 17332
rect 38068 17320 38074 17332
rect 38565 17323 38623 17329
rect 38565 17320 38577 17323
rect 38068 17292 38577 17320
rect 38068 17280 38074 17292
rect 38565 17289 38577 17292
rect 38611 17289 38623 17323
rect 40034 17320 40040 17332
rect 38565 17283 38623 17289
rect 38948 17292 40040 17320
rect 35529 17255 35587 17261
rect 35529 17252 35541 17255
rect 34624 17224 35541 17252
rect 35529 17221 35541 17224
rect 35575 17221 35587 17255
rect 35529 17215 35587 17221
rect 36538 17212 36544 17264
rect 36596 17212 36602 17264
rect 37476 17224 38424 17252
rect 33137 17187 33195 17193
rect 33137 17153 33149 17187
rect 33183 17153 33195 17187
rect 33137 17147 33195 17153
rect 32815 17088 33088 17116
rect 33152 17116 33180 17147
rect 33226 17144 33232 17196
rect 33284 17144 33290 17196
rect 33594 17144 33600 17196
rect 33652 17144 33658 17196
rect 33778 17144 33784 17196
rect 33836 17144 33842 17196
rect 34241 17187 34299 17193
rect 34241 17153 34253 17187
rect 34287 17153 34299 17187
rect 34241 17147 34299 17153
rect 33502 17116 33508 17128
rect 33152 17088 33508 17116
rect 32815 17085 32827 17088
rect 32769 17079 32827 17085
rect 25961 17011 26019 17017
rect 26068 17020 28580 17048
rect 31021 17051 31079 17057
rect 25406 16980 25412 16992
rect 23676 16952 25412 16980
rect 23017 16943 23075 16949
rect 25406 16940 25412 16952
rect 25464 16980 25470 16992
rect 26068 16980 26096 17020
rect 31021 17017 31033 17051
rect 31067 17048 31079 17051
rect 31680 17048 31708 17079
rect 33502 17076 33508 17088
rect 33560 17076 33566 17128
rect 34256 17116 34284 17147
rect 34514 17144 34520 17196
rect 34572 17144 34578 17196
rect 34790 17144 34796 17196
rect 34848 17144 34854 17196
rect 34885 17187 34943 17193
rect 34885 17153 34897 17187
rect 34931 17153 34943 17187
rect 34885 17147 34943 17153
rect 34900 17116 34928 17147
rect 34974 17144 34980 17196
rect 35032 17144 35038 17196
rect 37476 17193 37504 17224
rect 35161 17187 35219 17193
rect 35161 17153 35173 17187
rect 35207 17153 35219 17187
rect 35161 17147 35219 17153
rect 37461 17187 37519 17193
rect 37461 17153 37473 17187
rect 37507 17153 37519 17187
rect 37461 17147 37519 17153
rect 35066 17116 35072 17128
rect 34256 17088 34468 17116
rect 31067 17020 31708 17048
rect 31067 17017 31079 17020
rect 31021 17011 31079 17017
rect 31846 17008 31852 17060
rect 31904 17048 31910 17060
rect 32861 17051 32919 17057
rect 32861 17048 32873 17051
rect 31904 17020 32873 17048
rect 31904 17008 31910 17020
rect 32861 17017 32873 17020
rect 32907 17017 32919 17051
rect 32861 17011 32919 17017
rect 33413 17051 33471 17057
rect 33413 17017 33425 17051
rect 33459 17048 33471 17051
rect 34440 17048 34468 17088
rect 34900 17088 35072 17116
rect 33459 17020 34468 17048
rect 33459 17017 33471 17020
rect 33413 17011 33471 17017
rect 25464 16952 26096 16980
rect 25464 16940 25470 16952
rect 27798 16940 27804 16992
rect 27856 16940 27862 16992
rect 30282 16940 30288 16992
rect 30340 16980 30346 16992
rect 32309 16983 32367 16989
rect 32309 16980 32321 16983
rect 30340 16952 32321 16980
rect 30340 16940 30346 16952
rect 32309 16949 32321 16952
rect 32355 16949 32367 16983
rect 32309 16943 32367 16949
rect 32490 16940 32496 16992
rect 32548 16940 32554 16992
rect 33318 16940 33324 16992
rect 33376 16940 33382 16992
rect 34054 16940 34060 16992
rect 34112 16980 34118 16992
rect 34333 16983 34391 16989
rect 34333 16980 34345 16983
rect 34112 16952 34345 16980
rect 34112 16940 34118 16952
rect 34333 16949 34345 16952
rect 34379 16949 34391 16983
rect 34440 16980 34468 17020
rect 34514 17008 34520 17060
rect 34572 17048 34578 17060
rect 34900 17048 34928 17088
rect 35066 17076 35072 17088
rect 35124 17076 35130 17128
rect 34572 17020 34928 17048
rect 35176 17048 35204 17147
rect 38010 17144 38016 17196
rect 38068 17184 38074 17196
rect 38105 17187 38163 17193
rect 38105 17184 38117 17187
rect 38068 17156 38117 17184
rect 38068 17144 38074 17156
rect 38105 17153 38117 17156
rect 38151 17153 38163 17187
rect 38105 17147 38163 17153
rect 38197 17187 38255 17193
rect 38197 17153 38209 17187
rect 38243 17153 38255 17187
rect 38197 17147 38255 17153
rect 38289 17187 38347 17193
rect 38289 17153 38301 17187
rect 38335 17153 38347 17187
rect 38289 17147 38347 17153
rect 35250 17076 35256 17128
rect 35308 17076 35314 17128
rect 35360 17088 37504 17116
rect 35360 17048 35388 17088
rect 35176 17020 35388 17048
rect 34572 17008 34578 17020
rect 35710 16980 35716 16992
rect 34440 16952 35716 16980
rect 34333 16943 34391 16949
rect 35710 16940 35716 16952
rect 35768 16940 35774 16992
rect 36998 16940 37004 16992
rect 37056 16940 37062 16992
rect 37476 16980 37504 17088
rect 37550 17076 37556 17128
rect 37608 17076 37614 17128
rect 37918 17076 37924 17128
rect 37976 17116 37982 17128
rect 38212 17116 38240 17147
rect 37976 17088 38240 17116
rect 37976 17076 37982 17088
rect 37829 17051 37887 17057
rect 37829 17017 37841 17051
rect 37875 17048 37887 17051
rect 38304 17048 38332 17147
rect 38396 17116 38424 17224
rect 38838 17212 38844 17264
rect 38896 17212 38902 17264
rect 38948 17261 38976 17292
rect 40034 17280 40040 17292
rect 40092 17280 40098 17332
rect 40126 17280 40132 17332
rect 40184 17320 40190 17332
rect 41969 17323 42027 17329
rect 41969 17320 41981 17323
rect 40184 17292 41981 17320
rect 40184 17280 40190 17292
rect 41969 17289 41981 17292
rect 42015 17289 42027 17323
rect 41969 17283 42027 17289
rect 38933 17255 38991 17261
rect 38933 17221 38945 17255
rect 38979 17221 38991 17255
rect 39761 17255 39819 17261
rect 38933 17215 38991 17221
rect 39040 17224 39712 17252
rect 38470 17144 38476 17196
rect 38528 17144 38534 17196
rect 38562 17144 38568 17196
rect 38620 17184 38626 17196
rect 38749 17187 38807 17193
rect 38749 17184 38761 17187
rect 38620 17156 38761 17184
rect 38620 17144 38626 17156
rect 38749 17153 38761 17156
rect 38795 17153 38807 17187
rect 38749 17147 38807 17153
rect 39040 17116 39068 17224
rect 39117 17187 39175 17193
rect 39117 17153 39129 17187
rect 39163 17153 39175 17187
rect 39117 17147 39175 17153
rect 38396 17088 39068 17116
rect 37875 17020 38332 17048
rect 37875 17017 37887 17020
rect 37829 17011 37887 17017
rect 38470 17008 38476 17060
rect 38528 17048 38534 17060
rect 39132 17048 39160 17147
rect 39574 17144 39580 17196
rect 39632 17144 39638 17196
rect 39684 17116 39712 17224
rect 39761 17221 39773 17255
rect 39807 17252 39819 17255
rect 41141 17255 41199 17261
rect 41141 17252 41153 17255
rect 39807 17224 41153 17252
rect 39807 17221 39819 17224
rect 39761 17215 39819 17221
rect 41141 17221 41153 17224
rect 41187 17221 41199 17255
rect 41141 17215 41199 17221
rect 39850 17144 39856 17196
rect 39908 17144 39914 17196
rect 39942 17144 39948 17196
rect 40000 17144 40006 17196
rect 41785 17187 41843 17193
rect 40052 17156 41414 17184
rect 40052 17116 40080 17156
rect 39684 17088 40080 17116
rect 40405 17119 40463 17125
rect 40405 17085 40417 17119
rect 40451 17085 40463 17119
rect 40405 17079 40463 17085
rect 38528 17020 39160 17048
rect 40129 17051 40187 17057
rect 38528 17008 38534 17020
rect 40129 17017 40141 17051
rect 40175 17048 40187 17051
rect 40420 17048 40448 17079
rect 40175 17020 40448 17048
rect 41386 17048 41414 17156
rect 41785 17153 41797 17187
rect 41831 17184 41843 17187
rect 41877 17187 41935 17193
rect 41877 17184 41889 17187
rect 41831 17156 41889 17184
rect 41831 17153 41843 17156
rect 41785 17147 41843 17153
rect 41877 17153 41889 17156
rect 41923 17184 41935 17187
rect 41966 17184 41972 17196
rect 41923 17156 41972 17184
rect 41923 17153 41935 17156
rect 41877 17147 41935 17153
rect 41966 17144 41972 17156
rect 42024 17144 42030 17196
rect 42061 17187 42119 17193
rect 42061 17153 42073 17187
rect 42107 17184 42119 17187
rect 42150 17184 42156 17196
rect 42107 17156 42156 17184
rect 42107 17153 42119 17156
rect 42061 17147 42119 17153
rect 42150 17144 42156 17156
rect 42208 17144 42214 17196
rect 41690 17048 41696 17060
rect 41386 17020 41696 17048
rect 40175 17017 40187 17020
rect 40129 17011 40187 17017
rect 41690 17008 41696 17020
rect 41748 17008 41754 17060
rect 39574 16980 39580 16992
rect 37476 16952 39580 16980
rect 39574 16940 39580 16952
rect 39632 16980 39638 16992
rect 40402 16980 40408 16992
rect 39632 16952 40408 16980
rect 39632 16940 39638 16952
rect 40402 16940 40408 16952
rect 40460 16940 40466 16992
rect 40494 16940 40500 16992
rect 40552 16980 40558 16992
rect 41049 16983 41107 16989
rect 41049 16980 41061 16983
rect 40552 16952 41061 16980
rect 40552 16940 40558 16952
rect 41049 16949 41061 16952
rect 41095 16949 41107 16983
rect 41049 16943 41107 16949
rect 1104 16890 42504 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 42504 16890
rect 1104 16816 42504 16838
rect 5077 16779 5135 16785
rect 5077 16745 5089 16779
rect 5123 16776 5135 16779
rect 5626 16776 5632 16788
rect 5123 16748 5632 16776
rect 5123 16745 5135 16748
rect 5077 16739 5135 16745
rect 5626 16736 5632 16748
rect 5684 16736 5690 16788
rect 5994 16736 6000 16788
rect 6052 16776 6058 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 6052 16748 6285 16776
rect 6052 16736 6058 16748
rect 6273 16745 6285 16748
rect 6319 16776 6331 16779
rect 6546 16776 6552 16788
rect 6319 16748 6552 16776
rect 6319 16745 6331 16748
rect 6273 16739 6331 16745
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 8110 16776 8116 16788
rect 8067 16748 8116 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 8205 16779 8263 16785
rect 8205 16745 8217 16779
rect 8251 16776 8263 16779
rect 8941 16779 8999 16785
rect 8941 16776 8953 16779
rect 8251 16748 8953 16776
rect 8251 16745 8263 16748
rect 8205 16739 8263 16745
rect 8941 16745 8953 16748
rect 8987 16745 8999 16779
rect 8941 16739 8999 16745
rect 10781 16779 10839 16785
rect 10781 16745 10793 16779
rect 10827 16745 10839 16779
rect 10781 16739 10839 16745
rect 4890 16668 4896 16720
rect 4948 16708 4954 16720
rect 5813 16711 5871 16717
rect 5813 16708 5825 16711
rect 4948 16680 5396 16708
rect 4948 16668 4954 16680
rect 5368 16652 5396 16680
rect 5552 16680 5825 16708
rect 1578 16600 1584 16652
rect 1636 16640 1642 16652
rect 1765 16643 1823 16649
rect 1765 16640 1777 16643
rect 1636 16612 1777 16640
rect 1636 16600 1642 16612
rect 1765 16609 1777 16612
rect 1811 16609 1823 16643
rect 1765 16603 1823 16609
rect 3191 16643 3249 16649
rect 3191 16609 3203 16643
rect 3237 16640 3249 16643
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3237 16612 4353 16640
rect 3237 16609 3249 16612
rect 3191 16603 3249 16609
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 5258 16600 5264 16652
rect 5316 16600 5322 16652
rect 5350 16600 5356 16652
rect 5408 16600 5414 16652
rect 5442 16600 5448 16652
rect 5500 16600 5506 16652
rect 5552 16649 5580 16680
rect 5813 16677 5825 16680
rect 5859 16677 5871 16711
rect 5813 16671 5871 16677
rect 5902 16668 5908 16720
rect 5960 16708 5966 16720
rect 10796 16708 10824 16739
rect 10870 16736 10876 16788
rect 10928 16776 10934 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10928 16748 10977 16776
rect 10928 16736 10934 16748
rect 10965 16745 10977 16748
rect 11011 16745 11023 16779
rect 10965 16739 11023 16745
rect 11422 16736 11428 16788
rect 11480 16736 11486 16788
rect 12342 16776 12348 16788
rect 11624 16748 12348 16776
rect 11054 16708 11060 16720
rect 5960 16680 6408 16708
rect 10796 16680 11060 16708
rect 5960 16668 5966 16680
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16609 5595 16643
rect 5537 16603 5595 16609
rect 5721 16643 5779 16649
rect 5721 16609 5733 16643
rect 5767 16640 5779 16643
rect 6178 16640 6184 16652
rect 5767 16612 6184 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16572 1455 16575
rect 1670 16572 1676 16584
rect 1443 16544 1676 16572
rect 1443 16541 1455 16544
rect 1397 16535 1455 16541
rect 1670 16532 1676 16544
rect 1728 16532 1734 16584
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 6380 16581 6408 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 9309 16643 9367 16649
rect 9309 16609 9321 16643
rect 9355 16640 9367 16643
rect 9950 16640 9956 16652
rect 9355 16612 9956 16640
rect 9355 16609 9367 16612
rect 9309 16603 9367 16609
rect 9950 16600 9956 16612
rect 10008 16640 10014 16652
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 10008 16612 10609 16640
rect 10008 16600 10014 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 4856 16544 5304 16572
rect 4856 16532 4862 16544
rect 2774 16464 2780 16516
rect 2832 16504 2838 16516
rect 3970 16504 3976 16516
rect 2832 16476 3976 16504
rect 2832 16464 2838 16476
rect 3970 16464 3976 16476
rect 4028 16464 4034 16516
rect 4890 16464 4896 16516
rect 4948 16464 4954 16516
rect 5077 16507 5135 16513
rect 5077 16473 5089 16507
rect 5123 16504 5135 16507
rect 5166 16504 5172 16516
rect 5123 16476 5172 16504
rect 5123 16473 5135 16476
rect 5077 16467 5135 16473
rect 5166 16464 5172 16476
rect 5224 16464 5230 16516
rect 5276 16504 5304 16544
rect 5460 16544 6009 16572
rect 5460 16504 5488 16544
rect 5997 16541 6009 16544
rect 6043 16541 6055 16575
rect 5997 16535 6055 16541
rect 6365 16575 6423 16581
rect 6365 16541 6377 16575
rect 6411 16541 6423 16575
rect 6365 16535 6423 16541
rect 8478 16532 8484 16584
rect 8536 16532 8542 16584
rect 9122 16532 9128 16584
rect 9180 16532 9186 16584
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 5276 16476 5488 16504
rect 8389 16507 8447 16513
rect 8389 16473 8401 16507
rect 8435 16504 8447 16507
rect 8662 16504 8668 16516
rect 8435 16476 8668 16504
rect 8435 16473 8447 16476
rect 8389 16467 8447 16473
rect 8662 16464 8668 16476
rect 8720 16504 8726 16516
rect 8846 16504 8852 16516
rect 8720 16476 8852 16504
rect 8720 16464 8726 16476
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 9232 16504 9260 16535
rect 9398 16532 9404 16584
rect 9456 16532 9462 16584
rect 11624 16581 11652 16748
rect 12342 16736 12348 16748
rect 12400 16776 12406 16788
rect 12621 16779 12679 16785
rect 12621 16776 12633 16779
rect 12400 16748 12633 16776
rect 12400 16736 12406 16748
rect 12621 16745 12633 16748
rect 12667 16745 12679 16779
rect 12621 16739 12679 16745
rect 12802 16736 12808 16788
rect 12860 16736 12866 16788
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12952 16748 13093 16776
rect 12952 16736 12958 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13081 16739 13139 16745
rect 13262 16736 13268 16788
rect 13320 16736 13326 16788
rect 13906 16736 13912 16788
rect 13964 16736 13970 16788
rect 20806 16736 20812 16788
rect 20864 16736 20870 16788
rect 23753 16779 23811 16785
rect 23753 16745 23765 16779
rect 23799 16776 23811 16779
rect 23842 16776 23848 16788
rect 23799 16748 23848 16776
rect 23799 16745 23811 16748
rect 23753 16739 23811 16745
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 24394 16736 24400 16788
rect 24452 16736 24458 16788
rect 24762 16736 24768 16788
rect 24820 16776 24826 16788
rect 25777 16779 25835 16785
rect 25777 16776 25789 16779
rect 24820 16748 25789 16776
rect 24820 16736 24826 16748
rect 25777 16745 25789 16748
rect 25823 16745 25835 16779
rect 25777 16739 25835 16745
rect 28074 16736 28080 16788
rect 28132 16776 28138 16788
rect 28905 16779 28963 16785
rect 28905 16776 28917 16779
rect 28132 16748 28917 16776
rect 28132 16736 28138 16748
rect 28905 16745 28917 16748
rect 28951 16745 28963 16779
rect 28905 16739 28963 16745
rect 29086 16736 29092 16788
rect 29144 16776 29150 16788
rect 30282 16776 30288 16788
rect 29144 16748 30288 16776
rect 29144 16736 29150 16748
rect 30282 16736 30288 16748
rect 30340 16736 30346 16788
rect 32490 16736 32496 16788
rect 32548 16776 32554 16788
rect 32548 16748 34376 16776
rect 32548 16736 32554 16748
rect 17034 16668 17040 16720
rect 17092 16668 17098 16720
rect 25133 16711 25191 16717
rect 25133 16708 25145 16711
rect 25056 16680 25145 16708
rect 13630 16640 13636 16652
rect 11716 16612 11928 16640
rect 11716 16581 11744 16612
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16541 10839 16575
rect 10781 16535 10839 16541
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 11701 16575 11759 16581
rect 11701 16541 11713 16575
rect 11747 16541 11759 16575
rect 11701 16535 11759 16541
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16541 11851 16575
rect 11900 16572 11928 16612
rect 12820 16612 13636 16640
rect 11900 16544 12112 16572
rect 11793 16535 11851 16541
rect 9674 16504 9680 16516
rect 9232 16476 9680 16504
rect 9674 16464 9680 16476
rect 9732 16504 9738 16516
rect 10318 16504 10324 16516
rect 9732 16476 10324 16504
rect 9732 16464 9738 16476
rect 10318 16464 10324 16476
rect 10376 16504 10382 16516
rect 10505 16507 10563 16513
rect 10505 16504 10517 16507
rect 10376 16476 10517 16504
rect 10376 16464 10382 16476
rect 10505 16473 10517 16476
rect 10551 16473 10563 16507
rect 10796 16504 10824 16535
rect 11808 16504 11836 16535
rect 11974 16504 11980 16516
rect 10796 16476 11980 16504
rect 10505 16467 10563 16473
rect 11974 16464 11980 16476
rect 12032 16464 12038 16516
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3016 16408 3801 16436
rect 3016 16396 3022 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 5184 16436 5212 16464
rect 5626 16436 5632 16448
rect 5184 16408 5632 16436
rect 3789 16399 3847 16405
rect 5626 16396 5632 16408
rect 5684 16396 5690 16448
rect 8189 16439 8247 16445
rect 8189 16405 8201 16439
rect 8235 16436 8247 16439
rect 8573 16439 8631 16445
rect 8573 16436 8585 16439
rect 8235 16408 8585 16436
rect 8235 16405 8247 16408
rect 8189 16399 8247 16405
rect 8573 16405 8585 16408
rect 8619 16405 8631 16439
rect 8573 16399 8631 16405
rect 11882 16396 11888 16448
rect 11940 16436 11946 16448
rect 12084 16436 12112 16544
rect 12434 16464 12440 16516
rect 12492 16464 12498 16516
rect 12618 16464 12624 16516
rect 12676 16513 12682 16516
rect 12676 16507 12711 16513
rect 12699 16504 12711 16507
rect 12820 16504 12848 16612
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 17052 16640 17080 16668
rect 20625 16643 20683 16649
rect 20625 16640 20637 16643
rect 15979 16612 17080 16640
rect 19720 16612 20637 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 19720 16584 19748 16612
rect 20625 16609 20637 16612
rect 20671 16609 20683 16643
rect 20625 16603 20683 16609
rect 21376 16612 21588 16640
rect 13538 16532 13544 16584
rect 13596 16532 13602 16584
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 15470 16572 15476 16584
rect 15252 16544 15476 16572
rect 15252 16532 15258 16544
rect 15470 16532 15476 16544
rect 15528 16572 15534 16584
rect 15657 16575 15715 16581
rect 15657 16572 15669 16575
rect 15528 16544 15669 16572
rect 15528 16532 15534 16544
rect 15657 16541 15669 16544
rect 15703 16541 15715 16575
rect 15657 16535 15715 16541
rect 17494 16532 17500 16584
rect 17552 16532 17558 16584
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 18196 16544 18337 16572
rect 18196 16532 18202 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16572 18567 16575
rect 18690 16572 18696 16584
rect 18555 16544 18696 16572
rect 18555 16541 18567 16544
rect 18509 16535 18567 16541
rect 12699 16476 12848 16504
rect 12699 16473 12711 16476
rect 12676 16467 12711 16473
rect 12676 16464 12682 16467
rect 12894 16464 12900 16516
rect 12952 16464 12958 16516
rect 12986 16464 12992 16516
rect 13044 16504 13050 16516
rect 13097 16507 13155 16513
rect 13097 16504 13109 16507
rect 13044 16476 13109 16504
rect 13044 16464 13050 16476
rect 13097 16473 13109 16476
rect 13143 16473 13155 16507
rect 13097 16467 13155 16473
rect 15378 16464 15384 16516
rect 15436 16504 15442 16516
rect 16206 16504 16212 16516
rect 15436 16476 16212 16504
rect 15436 16464 15442 16476
rect 16206 16464 16212 16476
rect 16264 16504 16270 16516
rect 18340 16504 18368 16535
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 18785 16575 18843 16581
rect 18785 16541 18797 16575
rect 18831 16572 18843 16575
rect 18966 16572 18972 16584
rect 18831 16544 18972 16572
rect 18831 16541 18843 16544
rect 18785 16535 18843 16541
rect 18800 16504 18828 16535
rect 18966 16532 18972 16544
rect 19024 16532 19030 16584
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16572 19487 16575
rect 19702 16572 19708 16584
rect 19475 16544 19708 16572
rect 19475 16541 19487 16544
rect 19429 16535 19487 16541
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 20073 16575 20131 16581
rect 19852 16544 20024 16572
rect 19852 16532 19858 16544
rect 16264 16476 16422 16504
rect 17420 16476 18828 16504
rect 16264 16464 16270 16476
rect 12802 16436 12808 16448
rect 11940 16408 12808 16436
rect 11940 16396 11946 16408
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 17420 16445 17448 16476
rect 19518 16464 19524 16516
rect 19576 16464 19582 16516
rect 19613 16507 19671 16513
rect 19613 16473 19625 16507
rect 19659 16504 19671 16507
rect 19886 16504 19892 16516
rect 19659 16476 19892 16504
rect 19659 16473 19671 16476
rect 19613 16467 19671 16473
rect 19886 16464 19892 16476
rect 19944 16464 19950 16516
rect 19996 16504 20024 16544
rect 20073 16541 20085 16575
rect 20119 16572 20131 16575
rect 20254 16572 20260 16584
rect 20119 16544 20260 16572
rect 20119 16541 20131 16544
rect 20073 16535 20131 16541
rect 20254 16532 20260 16544
rect 20312 16532 20318 16584
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 21376 16581 21404 16612
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20772 16544 21005 16572
rect 20772 16532 20778 16544
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 21085 16575 21143 16581
rect 21085 16541 21097 16575
rect 21131 16572 21143 16575
rect 21361 16575 21419 16581
rect 21131 16544 21312 16572
rect 21131 16541 21143 16544
rect 21085 16535 21143 16541
rect 19996 16476 20760 16504
rect 17405 16439 17463 16445
rect 17405 16405 17417 16439
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 18138 16396 18144 16448
rect 18196 16396 18202 16448
rect 18414 16396 18420 16448
rect 18472 16396 18478 16448
rect 18782 16396 18788 16448
rect 18840 16436 18846 16448
rect 18969 16439 19027 16445
rect 18969 16436 18981 16439
rect 18840 16408 18981 16436
rect 18840 16396 18846 16408
rect 18969 16405 18981 16408
rect 19015 16405 19027 16439
rect 18969 16399 19027 16405
rect 19150 16396 19156 16448
rect 19208 16436 19214 16448
rect 19245 16439 19303 16445
rect 19245 16436 19257 16439
rect 19208 16408 19257 16436
rect 19208 16396 19214 16408
rect 19245 16405 19257 16408
rect 19291 16405 19303 16439
rect 19536 16436 19564 16464
rect 20622 16436 20628 16448
rect 19536 16408 20628 16436
rect 19245 16399 19303 16405
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 20732 16436 20760 16476
rect 21174 16464 21180 16516
rect 21232 16464 21238 16516
rect 21284 16504 21312 16544
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 21450 16532 21456 16584
rect 21508 16532 21514 16584
rect 21560 16572 21588 16612
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 22152 16612 22416 16640
rect 22152 16600 22158 16612
rect 21726 16572 21732 16584
rect 21560 16544 21732 16572
rect 21726 16532 21732 16544
rect 21784 16532 21790 16584
rect 22388 16581 22416 16612
rect 24118 16600 24124 16652
rect 24176 16600 24182 16652
rect 25056 16649 25084 16680
rect 25133 16677 25145 16680
rect 25179 16677 25191 16711
rect 25133 16671 25191 16677
rect 25866 16668 25872 16720
rect 25924 16708 25930 16720
rect 27982 16708 27988 16720
rect 25924 16680 26280 16708
rect 25924 16668 25930 16680
rect 25041 16643 25099 16649
rect 25041 16609 25053 16643
rect 25087 16609 25099 16643
rect 25884 16640 25912 16668
rect 25041 16603 25099 16609
rect 25792 16612 25912 16640
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16541 22431 16575
rect 22373 16535 22431 16541
rect 22554 16532 22560 16584
rect 22612 16532 22618 16584
rect 22741 16575 22799 16581
rect 22741 16541 22753 16575
rect 22787 16572 22799 16575
rect 22922 16572 22928 16584
rect 22787 16544 22928 16572
rect 22787 16541 22799 16544
rect 22741 16535 22799 16541
rect 22922 16532 22928 16544
rect 22980 16532 22986 16584
rect 24029 16575 24087 16581
rect 24029 16541 24041 16575
rect 24075 16572 24087 16575
rect 24210 16572 24216 16584
rect 24075 16544 24216 16572
rect 24075 16541 24087 16544
rect 24029 16535 24087 16541
rect 24210 16532 24216 16544
rect 24268 16532 24274 16584
rect 24946 16532 24952 16584
rect 25004 16572 25010 16584
rect 25317 16575 25375 16581
rect 25317 16572 25329 16575
rect 25004 16544 25329 16572
rect 25004 16532 25010 16544
rect 25317 16541 25329 16544
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 25498 16532 25504 16584
rect 25556 16532 25562 16584
rect 25590 16532 25596 16584
rect 25648 16572 25654 16584
rect 25792 16581 25820 16612
rect 25685 16575 25743 16581
rect 25685 16572 25697 16575
rect 25648 16544 25697 16572
rect 25648 16532 25654 16544
rect 25685 16541 25697 16544
rect 25731 16541 25743 16575
rect 25685 16535 25743 16541
rect 25777 16575 25835 16581
rect 25777 16541 25789 16575
rect 25823 16541 25835 16575
rect 25777 16535 25835 16541
rect 25955 16575 26013 16581
rect 25955 16541 25967 16575
rect 26001 16574 26013 16575
rect 26050 16574 26056 16584
rect 26001 16546 26056 16574
rect 26001 16541 26013 16546
rect 25955 16535 26013 16541
rect 26050 16532 26056 16546
rect 26108 16532 26114 16584
rect 26252 16581 26280 16680
rect 27632 16680 27988 16708
rect 26878 16600 26884 16652
rect 26936 16640 26942 16652
rect 27632 16649 27660 16680
rect 27982 16668 27988 16680
rect 28040 16668 28046 16720
rect 28166 16668 28172 16720
rect 28224 16708 28230 16720
rect 29641 16711 29699 16717
rect 29641 16708 29653 16711
rect 28224 16680 29653 16708
rect 28224 16668 28230 16680
rect 29641 16677 29653 16680
rect 29687 16677 29699 16711
rect 29641 16671 29699 16677
rect 27617 16643 27675 16649
rect 26936 16612 27568 16640
rect 26936 16600 26942 16612
rect 26237 16575 26295 16581
rect 26237 16541 26249 16575
rect 26283 16541 26295 16575
rect 27540 16572 27568 16612
rect 27617 16609 27629 16643
rect 27663 16609 27675 16643
rect 27617 16603 27675 16609
rect 27709 16643 27767 16649
rect 27709 16609 27721 16643
rect 27755 16609 27767 16643
rect 27709 16603 27767 16609
rect 29288 16612 29868 16640
rect 27724 16572 27752 16603
rect 27540 16544 27752 16572
rect 26237 16535 26295 16541
rect 28534 16532 28540 16584
rect 28592 16572 28598 16584
rect 29288 16581 29316 16612
rect 28721 16575 28779 16581
rect 28721 16572 28733 16575
rect 28592 16544 28733 16572
rect 28592 16532 28598 16544
rect 28721 16541 28733 16544
rect 28767 16541 28779 16575
rect 28721 16535 28779 16541
rect 29089 16575 29147 16581
rect 29089 16541 29101 16575
rect 29135 16541 29147 16575
rect 29089 16535 29147 16541
rect 29273 16575 29331 16581
rect 29273 16541 29285 16575
rect 29319 16541 29331 16575
rect 29273 16535 29331 16541
rect 29365 16575 29423 16581
rect 29365 16541 29377 16575
rect 29411 16572 29423 16575
rect 29454 16572 29460 16584
rect 29411 16544 29460 16572
rect 29411 16541 29423 16544
rect 29365 16535 29423 16541
rect 21468 16504 21496 16532
rect 21284 16476 21496 16504
rect 22465 16507 22523 16513
rect 22465 16473 22477 16507
rect 22511 16504 22523 16507
rect 22830 16504 22836 16516
rect 22511 16476 22836 16504
rect 22511 16473 22523 16476
rect 22465 16467 22523 16473
rect 22830 16464 22836 16476
rect 22888 16504 22894 16516
rect 25409 16507 25467 16513
rect 25409 16504 25421 16507
rect 22888 16476 25421 16504
rect 22888 16464 22894 16476
rect 25409 16473 25421 16476
rect 25455 16504 25467 16507
rect 26142 16504 26148 16516
rect 25455 16476 26148 16504
rect 25455 16473 25467 16476
rect 25409 16467 25467 16473
rect 26142 16464 26148 16476
rect 26200 16464 26206 16516
rect 27525 16507 27583 16513
rect 27525 16473 27537 16507
rect 27571 16504 27583 16507
rect 28169 16507 28227 16513
rect 28169 16504 28181 16507
rect 27571 16476 28181 16504
rect 27571 16473 27583 16476
rect 27525 16467 27583 16473
rect 28169 16473 28181 16476
rect 28215 16473 28227 16507
rect 29104 16504 29132 16535
rect 29454 16532 29460 16544
rect 29512 16572 29518 16584
rect 29840 16581 29868 16612
rect 30190 16600 30196 16652
rect 30248 16600 30254 16652
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29512 16544 29745 16572
rect 29512 16532 29518 16544
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 29825 16575 29883 16581
rect 29825 16541 29837 16575
rect 29871 16572 29883 16575
rect 30208 16572 30236 16600
rect 29871 16544 30236 16572
rect 30300 16558 30328 16736
rect 33045 16711 33103 16717
rect 33045 16677 33057 16711
rect 33091 16708 33103 16711
rect 33502 16708 33508 16720
rect 33091 16680 33508 16708
rect 33091 16677 33103 16680
rect 33045 16671 33103 16677
rect 33502 16668 33508 16680
rect 33560 16668 33566 16720
rect 34348 16708 34376 16748
rect 34790 16736 34796 16788
rect 34848 16736 34854 16788
rect 34882 16736 34888 16788
rect 34940 16776 34946 16788
rect 35989 16779 36047 16785
rect 35989 16776 36001 16779
rect 34940 16748 36001 16776
rect 34940 16736 34946 16748
rect 35989 16745 36001 16748
rect 36035 16745 36047 16779
rect 35989 16739 36047 16745
rect 38010 16736 38016 16788
rect 38068 16776 38074 16788
rect 38562 16776 38568 16788
rect 38068 16748 38568 16776
rect 38068 16736 38074 16748
rect 38562 16736 38568 16748
rect 38620 16736 38626 16788
rect 36081 16711 36139 16717
rect 36081 16708 36093 16711
rect 34348 16680 36093 16708
rect 36081 16677 36093 16680
rect 36127 16677 36139 16711
rect 36081 16671 36139 16677
rect 38856 16680 40264 16708
rect 31665 16643 31723 16649
rect 31665 16609 31677 16643
rect 31711 16640 31723 16643
rect 31754 16640 31760 16652
rect 31711 16612 31760 16640
rect 31711 16609 31723 16612
rect 31665 16603 31723 16609
rect 31754 16600 31760 16612
rect 31812 16640 31818 16652
rect 31938 16640 31944 16652
rect 31812 16612 31944 16640
rect 31812 16600 31818 16612
rect 31938 16600 31944 16612
rect 31996 16600 32002 16652
rect 32125 16643 32183 16649
rect 32125 16609 32137 16643
rect 32171 16640 32183 16643
rect 32677 16643 32735 16649
rect 32677 16640 32689 16643
rect 32171 16612 32689 16640
rect 32171 16609 32183 16612
rect 32125 16603 32183 16609
rect 32677 16609 32689 16612
rect 32723 16640 32735 16643
rect 33318 16640 33324 16652
rect 32723 16612 33324 16640
rect 32723 16609 32735 16612
rect 32677 16603 32735 16609
rect 33318 16600 33324 16612
rect 33376 16600 33382 16652
rect 34882 16640 34888 16652
rect 33980 16612 34888 16640
rect 33980 16581 34008 16612
rect 34882 16600 34888 16612
rect 34940 16600 34946 16652
rect 35345 16643 35403 16649
rect 35345 16640 35357 16643
rect 35268 16612 35357 16640
rect 35268 16584 35296 16612
rect 35345 16609 35357 16612
rect 35391 16609 35403 16643
rect 35345 16603 35403 16609
rect 37458 16600 37464 16652
rect 37516 16640 37522 16652
rect 38856 16649 38884 16680
rect 40236 16649 40264 16680
rect 38841 16643 38899 16649
rect 38841 16640 38853 16643
rect 37516 16612 38853 16640
rect 37516 16600 37522 16612
rect 38841 16609 38853 16612
rect 38887 16609 38899 16643
rect 38841 16603 38899 16609
rect 39853 16643 39911 16649
rect 39853 16609 39865 16643
rect 39899 16640 39911 16643
rect 40221 16643 40279 16649
rect 39899 16612 39988 16640
rect 39899 16609 39911 16612
rect 39853 16603 39911 16609
rect 32585 16575 32643 16581
rect 29871 16541 29883 16544
rect 29825 16535 29883 16541
rect 32585 16541 32597 16575
rect 32631 16572 32643 16575
rect 33965 16575 34023 16581
rect 32631 16544 32904 16572
rect 32631 16541 32643 16544
rect 32585 16535 32643 16541
rect 29549 16507 29607 16513
rect 29549 16504 29561 16507
rect 29104 16476 29561 16504
rect 28169 16467 28227 16473
rect 29380 16448 29408 16476
rect 29549 16473 29561 16476
rect 29595 16473 29607 16507
rect 29549 16467 29607 16473
rect 31386 16464 31392 16516
rect 31444 16464 31450 16516
rect 31754 16464 31760 16516
rect 31812 16464 31818 16516
rect 31941 16507 31999 16513
rect 31941 16473 31953 16507
rect 31987 16504 31999 16507
rect 32030 16504 32036 16516
rect 31987 16476 32036 16504
rect 31987 16473 31999 16476
rect 31941 16467 31999 16473
rect 32030 16464 32036 16476
rect 32088 16464 32094 16516
rect 22094 16436 22100 16448
rect 20732 16408 22100 16436
rect 22094 16396 22100 16408
rect 22152 16396 22158 16448
rect 22186 16396 22192 16448
rect 22244 16396 22250 16448
rect 25038 16396 25044 16448
rect 25096 16436 25102 16448
rect 26053 16439 26111 16445
rect 26053 16436 26065 16439
rect 25096 16408 26065 16436
rect 25096 16396 25102 16408
rect 26053 16405 26065 16408
rect 26099 16405 26111 16439
rect 26053 16399 26111 16405
rect 27157 16439 27215 16445
rect 27157 16405 27169 16439
rect 27203 16436 27215 16439
rect 27246 16436 27252 16448
rect 27203 16408 27252 16436
rect 27203 16405 27215 16408
rect 27157 16399 27215 16405
rect 27246 16396 27252 16408
rect 27304 16396 27310 16448
rect 29362 16396 29368 16448
rect 29420 16396 29426 16448
rect 29917 16439 29975 16445
rect 29917 16405 29929 16439
rect 29963 16436 29975 16439
rect 30374 16436 30380 16448
rect 29963 16408 30380 16436
rect 29963 16405 29975 16408
rect 29917 16399 29975 16405
rect 30374 16396 30380 16408
rect 30432 16396 30438 16448
rect 32214 16396 32220 16448
rect 32272 16396 32278 16448
rect 32876 16445 32904 16544
rect 33965 16541 33977 16575
rect 34011 16541 34023 16575
rect 33965 16535 34023 16541
rect 34054 16532 34060 16584
rect 34112 16532 34118 16584
rect 34425 16575 34483 16581
rect 34425 16541 34437 16575
rect 34471 16572 34483 16575
rect 34974 16572 34980 16584
rect 34471 16544 34980 16572
rect 34471 16541 34483 16544
rect 34425 16535 34483 16541
rect 34974 16532 34980 16544
rect 35032 16532 35038 16584
rect 35250 16532 35256 16584
rect 35308 16532 35314 16584
rect 35529 16575 35587 16581
rect 35529 16572 35541 16575
rect 35360 16544 35541 16572
rect 33226 16464 33232 16516
rect 33284 16504 33290 16516
rect 33321 16507 33379 16513
rect 33321 16504 33333 16507
rect 33284 16476 33333 16504
rect 33284 16464 33290 16476
rect 33321 16473 33333 16476
rect 33367 16473 33379 16507
rect 33321 16467 33379 16473
rect 34149 16507 34207 16513
rect 34149 16473 34161 16507
rect 34195 16473 34207 16507
rect 34149 16467 34207 16473
rect 34287 16507 34345 16513
rect 34287 16473 34299 16507
rect 34333 16504 34345 16507
rect 34790 16504 34796 16516
rect 34333 16476 34796 16504
rect 34333 16473 34345 16476
rect 34287 16467 34345 16473
rect 32861 16439 32919 16445
rect 32861 16405 32873 16439
rect 32907 16405 32919 16439
rect 32861 16399 32919 16405
rect 33778 16396 33784 16448
rect 33836 16396 33842 16448
rect 34054 16396 34060 16448
rect 34112 16436 34118 16448
rect 34164 16436 34192 16467
rect 34790 16464 34796 16476
rect 34848 16464 34854 16516
rect 35158 16464 35164 16516
rect 35216 16504 35222 16516
rect 35360 16504 35388 16544
rect 35529 16541 35541 16544
rect 35575 16541 35587 16575
rect 35529 16535 35587 16541
rect 35710 16532 35716 16584
rect 35768 16572 35774 16584
rect 35805 16575 35863 16581
rect 35805 16572 35817 16575
rect 35768 16544 35817 16572
rect 35768 16532 35774 16544
rect 35805 16541 35817 16544
rect 35851 16541 35863 16575
rect 35805 16535 35863 16541
rect 36354 16532 36360 16584
rect 36412 16532 36418 16584
rect 36541 16575 36599 16581
rect 36541 16541 36553 16575
rect 36587 16572 36599 16575
rect 36998 16572 37004 16584
rect 36587 16544 37004 16572
rect 36587 16541 36599 16544
rect 36541 16535 36599 16541
rect 35216 16476 35388 16504
rect 35216 16464 35222 16476
rect 35434 16464 35440 16516
rect 35492 16504 35498 16516
rect 35621 16507 35679 16513
rect 35621 16504 35633 16507
rect 35492 16476 35633 16504
rect 35492 16464 35498 16476
rect 35621 16473 35633 16476
rect 35667 16473 35679 16507
rect 36556 16504 36584 16535
rect 36998 16532 37004 16544
rect 37056 16532 37062 16584
rect 37366 16532 37372 16584
rect 37424 16572 37430 16584
rect 38105 16575 38163 16581
rect 38105 16572 38117 16575
rect 37424 16544 38117 16572
rect 37424 16532 37430 16544
rect 38105 16541 38117 16544
rect 38151 16572 38163 16575
rect 38194 16572 38200 16584
rect 38151 16544 38200 16572
rect 38151 16541 38163 16544
rect 38105 16535 38163 16541
rect 38194 16532 38200 16544
rect 38252 16532 38258 16584
rect 35621 16467 35679 16473
rect 36188 16476 36584 16504
rect 34112 16408 34192 16436
rect 34112 16396 34118 16408
rect 34698 16396 34704 16448
rect 34756 16436 34762 16448
rect 36188 16436 36216 16476
rect 34756 16408 36216 16436
rect 36265 16439 36323 16445
rect 34756 16396 34762 16408
rect 36265 16405 36277 16439
rect 36311 16436 36323 16439
rect 37550 16436 37556 16448
rect 36311 16408 37556 16436
rect 36311 16405 36323 16408
rect 36265 16399 36323 16405
rect 37550 16396 37556 16408
rect 37608 16396 37614 16448
rect 39114 16396 39120 16448
rect 39172 16436 39178 16448
rect 39853 16439 39911 16445
rect 39853 16436 39865 16439
rect 39172 16408 39865 16436
rect 39172 16396 39178 16408
rect 39853 16405 39865 16408
rect 39899 16405 39911 16439
rect 39960 16436 39988 16612
rect 40221 16609 40233 16643
rect 40267 16609 40279 16643
rect 40221 16603 40279 16609
rect 40494 16600 40500 16652
rect 40552 16600 40558 16652
rect 40037 16575 40095 16581
rect 40037 16541 40049 16575
rect 40083 16541 40095 16575
rect 40037 16535 40095 16541
rect 40052 16504 40080 16535
rect 40126 16532 40132 16584
rect 40184 16532 40190 16584
rect 41598 16532 41604 16584
rect 41656 16532 41662 16584
rect 40494 16504 40500 16516
rect 40052 16476 40500 16504
rect 40494 16464 40500 16476
rect 40552 16464 40558 16516
rect 40034 16436 40040 16448
rect 39960 16408 40040 16436
rect 39853 16399 39911 16405
rect 40034 16396 40040 16408
rect 40092 16396 40098 16448
rect 41966 16396 41972 16448
rect 42024 16396 42030 16448
rect 1104 16346 42504 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 42504 16346
rect 1104 16272 42504 16294
rect 5445 16235 5503 16241
rect 5445 16201 5457 16235
rect 5491 16232 5503 16235
rect 6362 16232 6368 16244
rect 5491 16204 6368 16232
rect 5491 16201 5503 16204
rect 5445 16195 5503 16201
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 8478 16192 8484 16244
rect 8536 16232 8542 16244
rect 8573 16235 8631 16241
rect 8573 16232 8585 16235
rect 8536 16204 8585 16232
rect 8536 16192 8542 16204
rect 8573 16201 8585 16204
rect 8619 16201 8631 16235
rect 8573 16195 8631 16201
rect 8846 16192 8852 16244
rect 8904 16232 8910 16244
rect 12066 16232 12072 16244
rect 8904 16204 12072 16232
rect 8904 16192 8910 16204
rect 12066 16192 12072 16204
rect 12124 16232 12130 16244
rect 12894 16232 12900 16244
rect 12124 16204 12900 16232
rect 12124 16192 12130 16204
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 13630 16192 13636 16244
rect 13688 16232 13694 16244
rect 15654 16232 15660 16244
rect 13688 16204 15660 16232
rect 13688 16192 13694 16204
rect 15654 16192 15660 16204
rect 15712 16232 15718 16244
rect 17681 16235 17739 16241
rect 17681 16232 17693 16235
rect 15712 16204 17693 16232
rect 15712 16192 15718 16204
rect 17681 16201 17693 16204
rect 17727 16201 17739 16235
rect 17681 16195 17739 16201
rect 18230 16192 18236 16244
rect 18288 16232 18294 16244
rect 20898 16232 20904 16244
rect 18288 16204 20904 16232
rect 18288 16192 18294 16204
rect 3970 16124 3976 16176
rect 4028 16124 4034 16176
rect 5534 16124 5540 16176
rect 5592 16164 5598 16176
rect 5721 16167 5779 16173
rect 5721 16164 5733 16167
rect 5592 16136 5733 16164
rect 5592 16124 5598 16136
rect 5721 16133 5733 16136
rect 5767 16133 5779 16167
rect 5721 16127 5779 16133
rect 8202 16124 8208 16176
rect 8260 16164 8266 16176
rect 8725 16167 8783 16173
rect 8725 16164 8737 16167
rect 8260 16136 8737 16164
rect 8260 16124 8266 16136
rect 8725 16133 8737 16136
rect 8771 16133 8783 16167
rect 8725 16127 8783 16133
rect 8941 16167 8999 16173
rect 8941 16133 8953 16167
rect 8987 16164 8999 16167
rect 9950 16164 9956 16176
rect 8987 16136 9956 16164
rect 8987 16133 8999 16136
rect 8941 16127 8999 16133
rect 9950 16124 9956 16136
rect 10008 16124 10014 16176
rect 11974 16124 11980 16176
rect 12032 16164 12038 16176
rect 12529 16167 12587 16173
rect 12529 16164 12541 16167
rect 12032 16136 12541 16164
rect 12032 16124 12038 16136
rect 12529 16133 12541 16136
rect 12575 16133 12587 16167
rect 12529 16127 12587 16133
rect 12618 16124 12624 16176
rect 12676 16164 12682 16176
rect 15105 16167 15163 16173
rect 12676 16136 13032 16164
rect 12676 16124 12682 16136
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 900 16068 1409 16096
rect 900 16056 906 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 2958 16056 2964 16108
rect 3016 16056 3022 16108
rect 4387 16099 4445 16105
rect 4387 16065 4399 16099
rect 4433 16096 4445 16099
rect 5350 16096 5356 16108
rect 4433 16068 5356 16096
rect 4433 16065 4445 16068
rect 4387 16059 4445 16065
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 5905 16099 5963 16105
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 5994 16096 6000 16108
rect 5951 16068 6000 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 6086 16056 6092 16108
rect 6144 16056 6150 16108
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16096 11759 16099
rect 12345 16099 12403 16105
rect 12345 16096 12357 16099
rect 11747 16068 12357 16096
rect 11747 16065 11759 16068
rect 11701 16059 11759 16065
rect 12345 16065 12357 16068
rect 12391 16065 12403 16099
rect 12345 16059 12403 16065
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16096 12495 16099
rect 12483 16068 12572 16096
rect 12483 16065 12495 16068
rect 12437 16059 12495 16065
rect 1762 15988 1768 16040
rect 1820 16028 1826 16040
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 1820 16000 2605 16028
rect 1820 15988 1826 16000
rect 2593 15997 2605 16000
rect 2639 15997 2651 16031
rect 2593 15991 2651 15997
rect 11054 15988 11060 16040
rect 11112 16028 11118 16040
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 11112 16000 11805 16028
rect 11112 15988 11118 16000
rect 11793 15997 11805 16000
rect 11839 15997 11851 16031
rect 11793 15991 11851 15997
rect 5350 15920 5356 15972
rect 5408 15960 5414 15972
rect 7742 15960 7748 15972
rect 5408 15932 7748 15960
rect 5408 15920 5414 15932
rect 7742 15920 7748 15932
rect 7800 15960 7806 15972
rect 11698 15960 11704 15972
rect 7800 15932 11704 15960
rect 7800 15920 7806 15932
rect 11698 15920 11704 15932
rect 11756 15920 11762 15972
rect 11808 15960 11836 15991
rect 11882 15988 11888 16040
rect 11940 15988 11946 16040
rect 11974 15988 11980 16040
rect 12032 15988 12038 16040
rect 12360 15960 12388 16059
rect 12434 15960 12440 15972
rect 11808 15932 12296 15960
rect 12360 15932 12440 15960
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 1670 15892 1676 15904
rect 1627 15864 1676 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 8757 15895 8815 15901
rect 8757 15861 8769 15895
rect 8803 15892 8815 15895
rect 9398 15892 9404 15904
rect 8803 15864 9404 15892
rect 8803 15861 8815 15864
rect 8757 15855 8815 15861
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 10744 15864 11529 15892
rect 10744 15852 10750 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 11606 15852 11612 15904
rect 11664 15892 11670 15904
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 11664 15864 12173 15892
rect 11664 15852 11670 15864
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 12268 15892 12296 15932
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 12544 15892 12572 16068
rect 12710 16056 12716 16108
rect 12768 16096 12774 16108
rect 13004 16105 13032 16136
rect 15105 16133 15117 16167
rect 15151 16164 15163 16167
rect 19628 16164 19656 16204
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 21085 16235 21143 16241
rect 21085 16201 21097 16235
rect 21131 16232 21143 16235
rect 21174 16232 21180 16244
rect 21131 16204 21180 16232
rect 21131 16201 21143 16204
rect 21085 16195 21143 16201
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 24118 16192 24124 16244
rect 24176 16192 24182 16244
rect 24210 16192 24216 16244
rect 24268 16192 24274 16244
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25590 16232 25596 16244
rect 24912 16204 25596 16232
rect 24912 16192 24918 16204
rect 25590 16192 25596 16204
rect 25648 16232 25654 16244
rect 28994 16232 29000 16244
rect 25648 16204 29000 16232
rect 25648 16192 25654 16204
rect 28994 16192 29000 16204
rect 29052 16192 29058 16244
rect 29362 16192 29368 16244
rect 29420 16192 29426 16244
rect 30926 16192 30932 16244
rect 30984 16232 30990 16244
rect 31113 16235 31171 16241
rect 31113 16232 31125 16235
rect 30984 16204 31125 16232
rect 30984 16192 30990 16204
rect 31113 16201 31125 16204
rect 31159 16201 31171 16235
rect 31113 16195 31171 16201
rect 31205 16235 31263 16241
rect 31205 16201 31217 16235
rect 31251 16232 31263 16235
rect 31386 16232 31392 16244
rect 31251 16204 31392 16232
rect 31251 16201 31263 16204
rect 31205 16195 31263 16201
rect 15151 16136 17540 16164
rect 19366 16136 19656 16164
rect 15151 16133 15163 16136
rect 15105 16127 15163 16133
rect 12805 16099 12863 16105
rect 12805 16096 12817 16099
rect 12768 16068 12817 16096
rect 12768 16056 12774 16068
rect 12805 16065 12817 16068
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 13262 16096 13268 16108
rect 13035 16068 13268 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 12820 15960 12848 16059
rect 13262 16056 13268 16068
rect 13320 16056 13326 16108
rect 13814 16056 13820 16108
rect 13872 16096 13878 16108
rect 14194 16099 14252 16105
rect 14194 16096 14206 16099
rect 13872 16068 14206 16096
rect 13872 16056 13878 16068
rect 14194 16065 14206 16068
rect 14240 16065 14252 16099
rect 14194 16059 14252 16065
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15378 16096 15384 16108
rect 15243 16068 15384 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15378 16056 15384 16068
rect 15436 16056 15442 16108
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16096 15807 16099
rect 15838 16096 15844 16108
rect 15795 16068 15844 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 14461 16031 14519 16037
rect 14461 15997 14473 16031
rect 14507 15997 14519 16031
rect 14461 15991 14519 15997
rect 13081 15963 13139 15969
rect 13081 15960 13093 15963
rect 12820 15932 13093 15960
rect 13081 15929 13093 15932
rect 13127 15960 13139 15963
rect 13354 15960 13360 15972
rect 13127 15932 13360 15960
rect 13127 15929 13139 15932
rect 13081 15923 13139 15929
rect 13354 15920 13360 15932
rect 13412 15920 13418 15972
rect 14476 15960 14504 15991
rect 15194 15960 15200 15972
rect 14476 15932 15200 15960
rect 15194 15920 15200 15932
rect 15252 15920 15258 15972
rect 15488 15960 15516 16059
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 16482 15988 16488 16040
rect 16540 15988 16546 16040
rect 17052 15960 17080 16059
rect 17126 16056 17132 16108
rect 17184 16056 17190 16108
rect 17512 16105 17540 16136
rect 19702 16124 19708 16176
rect 19760 16164 19766 16176
rect 20191 16167 20249 16173
rect 20191 16164 20203 16167
rect 19760 16136 20203 16164
rect 19760 16124 19766 16136
rect 20191 16133 20203 16136
rect 20237 16133 20249 16167
rect 20191 16127 20249 16133
rect 20806 16124 20812 16176
rect 20864 16164 20870 16176
rect 23750 16164 23756 16176
rect 20864 16136 23756 16164
rect 20864 16124 20870 16136
rect 23750 16124 23756 16136
rect 23808 16124 23814 16176
rect 17497 16099 17555 16105
rect 17497 16065 17509 16099
rect 17543 16065 17555 16099
rect 17497 16059 17555 16065
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 19484 16068 19901 16096
rect 19484 16056 19490 16068
rect 19889 16065 19901 16068
rect 19935 16065 19947 16099
rect 19889 16059 19947 16065
rect 19978 16056 19984 16108
rect 20036 16056 20042 16108
rect 20073 16099 20131 16105
rect 20073 16065 20085 16099
rect 20119 16065 20131 16099
rect 20073 16059 20131 16065
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 17310 15988 17316 16040
rect 17368 15988 17374 16040
rect 17402 15988 17408 16040
rect 17460 16028 17466 16040
rect 17865 16031 17923 16037
rect 17865 16028 17877 16031
rect 17460 16000 17877 16028
rect 17460 15988 17466 16000
rect 17865 15997 17877 16000
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 18141 16031 18199 16037
rect 18141 15997 18153 16031
rect 18187 16028 18199 16031
rect 20088 16028 20116 16059
rect 20162 16028 20168 16040
rect 18187 16000 19196 16028
rect 20088 16000 20168 16028
rect 18187 15997 18199 16000
rect 18141 15991 18199 15997
rect 19168 15960 19196 16000
rect 20162 15988 20168 16000
rect 20220 15988 20226 16040
rect 20349 16031 20407 16037
rect 20349 15997 20361 16031
rect 20395 15997 20407 16031
rect 20349 15991 20407 15997
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20732 16028 20760 16059
rect 21818 16056 21824 16108
rect 21876 16056 21882 16108
rect 22002 16056 22008 16108
rect 22060 16056 22066 16108
rect 23934 16056 23940 16108
rect 23992 16056 23998 16108
rect 24136 16096 24164 16192
rect 27246 16124 27252 16176
rect 27304 16124 27310 16176
rect 29086 16164 29092 16176
rect 28474 16136 29092 16164
rect 29086 16124 29092 16136
rect 29144 16124 29150 16176
rect 31128 16164 31156 16195
rect 31386 16192 31392 16204
rect 31444 16192 31450 16244
rect 34698 16192 34704 16244
rect 34756 16232 34762 16244
rect 34756 16204 35112 16232
rect 34756 16192 34762 16204
rect 31481 16167 31539 16173
rect 31481 16164 31493 16167
rect 31128 16136 31493 16164
rect 31481 16133 31493 16136
rect 31527 16133 31539 16167
rect 31481 16127 31539 16133
rect 31573 16167 31631 16173
rect 31573 16133 31585 16167
rect 31619 16164 31631 16167
rect 32214 16164 32220 16176
rect 31619 16136 32220 16164
rect 31619 16133 31631 16136
rect 31573 16127 31631 16133
rect 32214 16124 32220 16136
rect 32272 16124 32278 16176
rect 33778 16124 33784 16176
rect 33836 16124 33842 16176
rect 35084 16164 35112 16204
rect 35250 16192 35256 16244
rect 35308 16192 35314 16244
rect 37734 16192 37740 16244
rect 37792 16192 37798 16244
rect 35084 16136 35388 16164
rect 24857 16099 24915 16105
rect 24857 16096 24869 16099
rect 24136 16068 24869 16096
rect 24857 16065 24869 16068
rect 24903 16065 24915 16099
rect 24857 16059 24915 16065
rect 25038 16056 25044 16108
rect 25096 16056 25102 16108
rect 29641 16099 29699 16105
rect 29641 16096 29653 16099
rect 29288 16068 29653 16096
rect 29288 16040 29316 16068
rect 29641 16065 29653 16068
rect 29687 16065 29699 16099
rect 29641 16059 29699 16065
rect 30374 16056 30380 16108
rect 30432 16096 30438 16108
rect 30469 16099 30527 16105
rect 30469 16096 30481 16099
rect 30432 16068 30481 16096
rect 30432 16056 30438 16068
rect 30469 16065 30481 16068
rect 30515 16065 30527 16099
rect 30469 16059 30527 16065
rect 31389 16099 31447 16105
rect 31389 16065 31401 16099
rect 31435 16065 31447 16099
rect 31389 16059 31447 16065
rect 21177 16031 21235 16037
rect 21177 16028 21189 16031
rect 20732 16000 21189 16028
rect 20625 15991 20683 15997
rect 21177 15997 21189 16000
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 21637 16031 21695 16037
rect 21637 15997 21649 16031
rect 21683 16028 21695 16031
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21683 16000 21925 16028
rect 21683 15997 21695 16000
rect 21637 15991 21695 15997
rect 21913 15997 21925 16000
rect 21959 16028 21971 16031
rect 22186 16028 22192 16040
rect 21959 16000 22192 16028
rect 21959 15997 21971 16000
rect 21913 15991 21971 15997
rect 19705 15963 19763 15969
rect 19705 15960 19717 15963
rect 15488 15932 16804 15960
rect 17052 15932 17816 15960
rect 19168 15932 19717 15960
rect 12802 15892 12808 15904
rect 12268 15864 12808 15892
rect 12161 15855 12219 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 12986 15892 12992 15904
rect 12943 15864 12992 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 15289 15895 15347 15901
rect 15289 15861 15301 15895
rect 15335 15892 15347 15895
rect 15378 15892 15384 15904
rect 15335 15864 15384 15892
rect 15335 15861 15347 15864
rect 15289 15855 15347 15861
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 15838 15852 15844 15904
rect 15896 15852 15902 15904
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 16776 15892 16804 15932
rect 17310 15892 17316 15904
rect 16776 15864 17316 15892
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 17788 15892 17816 15932
rect 19705 15929 19717 15932
rect 19751 15929 19763 15963
rect 19705 15923 19763 15929
rect 18138 15892 18144 15904
rect 17788 15864 18144 15892
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 19613 15895 19671 15901
rect 19613 15861 19625 15895
rect 19659 15892 19671 15895
rect 20254 15892 20260 15904
rect 19659 15864 20260 15892
rect 19659 15861 19671 15864
rect 19613 15855 19671 15861
rect 20254 15852 20260 15864
rect 20312 15852 20318 15904
rect 20364 15892 20392 15991
rect 20640 15960 20668 15991
rect 22186 15988 22192 16000
rect 22244 15988 22250 16040
rect 24673 16031 24731 16037
rect 24673 15997 24685 16031
rect 24719 16028 24731 16031
rect 24762 16028 24768 16040
rect 24719 16000 24768 16028
rect 24719 15997 24731 16000
rect 24673 15991 24731 15997
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 26973 16031 27031 16037
rect 26973 15997 26985 16031
rect 27019 15997 27031 16031
rect 26973 15991 27031 15997
rect 20898 15960 20904 15972
rect 20640 15932 20904 15960
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 21358 15920 21364 15972
rect 21416 15920 21422 15972
rect 24397 15963 24455 15969
rect 24397 15929 24409 15963
rect 24443 15960 24455 15963
rect 25038 15960 25044 15972
rect 24443 15932 25044 15960
rect 24443 15929 24455 15932
rect 24397 15923 24455 15929
rect 25038 15920 25044 15932
rect 25096 15920 25102 15972
rect 26786 15960 26792 15972
rect 25148 15932 26792 15960
rect 20714 15892 20720 15904
rect 20364 15864 20720 15892
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 22922 15892 22928 15904
rect 22152 15864 22928 15892
rect 22152 15852 22158 15864
rect 22922 15852 22928 15864
rect 22980 15892 22986 15904
rect 25148 15892 25176 15932
rect 26786 15920 26792 15932
rect 26844 15920 26850 15972
rect 22980 15864 25176 15892
rect 25225 15895 25283 15901
rect 22980 15852 22986 15864
rect 25225 15861 25237 15895
rect 25271 15892 25283 15895
rect 26418 15892 26424 15904
rect 25271 15864 26424 15892
rect 25271 15861 25283 15864
rect 25225 15855 25283 15861
rect 26418 15852 26424 15864
rect 26476 15852 26482 15904
rect 26988 15892 27016 15991
rect 27798 15988 27804 16040
rect 27856 16028 27862 16040
rect 28718 16028 28724 16040
rect 27856 16000 28724 16028
rect 27856 15988 27862 16000
rect 28718 15988 28724 16000
rect 28776 16028 28782 16040
rect 28776 16000 29040 16028
rect 28776 15988 28782 16000
rect 28626 15920 28632 15972
rect 28684 15960 28690 15972
rect 28905 15963 28963 15969
rect 28905 15960 28917 15963
rect 28684 15932 28917 15960
rect 28684 15920 28690 15932
rect 28905 15929 28917 15932
rect 28951 15929 28963 15963
rect 29012 15960 29040 16000
rect 29270 15988 29276 16040
rect 29328 15988 29334 16040
rect 29365 16031 29423 16037
rect 29365 15997 29377 16031
rect 29411 16028 29423 16031
rect 29411 16000 29684 16028
rect 29411 15997 29423 16000
rect 29365 15991 29423 15997
rect 29549 15963 29607 15969
rect 29549 15960 29561 15963
rect 29012 15932 29561 15960
rect 28905 15923 28963 15929
rect 29549 15929 29561 15932
rect 29595 15929 29607 15963
rect 29549 15923 29607 15929
rect 27614 15892 27620 15904
rect 26988 15864 27620 15892
rect 27614 15852 27620 15864
rect 27672 15852 27678 15904
rect 28534 15852 28540 15904
rect 28592 15892 28598 15904
rect 28721 15895 28779 15901
rect 28721 15892 28733 15895
rect 28592 15864 28733 15892
rect 28592 15852 28598 15864
rect 28721 15861 28733 15864
rect 28767 15861 28779 15895
rect 28721 15855 28779 15861
rect 28810 15852 28816 15904
rect 28868 15852 28874 15904
rect 28920 15892 28948 15923
rect 29656 15892 29684 16000
rect 28920 15864 29684 15892
rect 31404 15892 31432 16059
rect 31662 16056 31668 16108
rect 31720 16096 31726 16108
rect 31757 16099 31815 16105
rect 31757 16096 31769 16099
rect 31720 16068 31769 16096
rect 31720 16056 31726 16068
rect 31757 16065 31769 16068
rect 31803 16096 31815 16099
rect 31803 16068 31892 16096
rect 31803 16065 31815 16068
rect 31757 16059 31815 16065
rect 31864 16028 31892 16068
rect 31938 16056 31944 16108
rect 31996 16096 32002 16108
rect 33505 16099 33563 16105
rect 33505 16096 33517 16099
rect 31996 16068 33517 16096
rect 31996 16056 32002 16068
rect 33505 16065 33517 16068
rect 33551 16065 33563 16099
rect 35250 16096 35256 16108
rect 34914 16068 35256 16096
rect 33505 16059 33563 16065
rect 35250 16056 35256 16068
rect 35308 16056 35314 16108
rect 35360 16105 35388 16136
rect 37458 16124 37464 16176
rect 37516 16164 37522 16176
rect 39761 16167 39819 16173
rect 37516 16136 38240 16164
rect 37516 16124 37522 16136
rect 35345 16099 35403 16105
rect 35345 16065 35357 16099
rect 35391 16065 35403 16099
rect 35345 16059 35403 16065
rect 35529 16099 35587 16105
rect 35529 16065 35541 16099
rect 35575 16096 35587 16099
rect 36354 16096 36360 16108
rect 35575 16068 36360 16096
rect 35575 16065 35587 16068
rect 35529 16059 35587 16065
rect 36354 16056 36360 16068
rect 36412 16056 36418 16108
rect 38212 16105 38240 16136
rect 39761 16133 39773 16167
rect 39807 16164 39819 16167
rect 41966 16164 41972 16176
rect 39807 16136 40632 16164
rect 39807 16133 39819 16136
rect 39761 16127 39819 16133
rect 37645 16099 37703 16105
rect 37645 16065 37657 16099
rect 37691 16096 37703 16099
rect 38197 16099 38255 16105
rect 37691 16068 38148 16096
rect 37691 16065 37703 16068
rect 37645 16059 37703 16065
rect 33870 16028 33876 16040
rect 31864 16000 33876 16028
rect 33870 15988 33876 16000
rect 33928 15988 33934 16040
rect 34422 15988 34428 16040
rect 34480 16028 34486 16040
rect 35158 16028 35164 16040
rect 34480 16000 35164 16028
rect 34480 15988 34486 16000
rect 35158 15988 35164 16000
rect 35216 16028 35222 16040
rect 35437 16031 35495 16037
rect 35437 16028 35449 16031
rect 35216 16000 35449 16028
rect 35216 15988 35222 16000
rect 35437 15997 35449 16000
rect 35483 15997 35495 16031
rect 35437 15991 35495 15997
rect 37921 16031 37979 16037
rect 37921 15997 37933 16031
rect 37967 15997 37979 16031
rect 38120 16028 38148 16068
rect 38197 16065 38209 16099
rect 38243 16065 38255 16099
rect 38197 16059 38255 16065
rect 40034 16056 40040 16108
rect 40092 16056 40098 16108
rect 40126 16056 40132 16108
rect 40184 16056 40190 16108
rect 40604 16105 40632 16136
rect 41616 16136 41972 16164
rect 40589 16099 40647 16105
rect 40589 16065 40601 16099
rect 40635 16065 40647 16099
rect 40589 16059 40647 16065
rect 41233 16099 41291 16105
rect 41233 16065 41245 16099
rect 41279 16096 41291 16099
rect 41322 16096 41328 16108
rect 41279 16068 41328 16096
rect 41279 16065 41291 16068
rect 41233 16059 41291 16065
rect 41322 16056 41328 16068
rect 41380 16056 41386 16108
rect 41616 16105 41644 16136
rect 41966 16124 41972 16136
rect 42024 16124 42030 16176
rect 41601 16099 41659 16105
rect 41601 16065 41613 16099
rect 41647 16065 41659 16099
rect 41601 16059 41659 16065
rect 41785 16099 41843 16105
rect 41785 16065 41797 16099
rect 41831 16096 41843 16099
rect 42058 16096 42064 16108
rect 41831 16068 42064 16096
rect 41831 16065 41843 16068
rect 41785 16059 41843 16065
rect 42058 16056 42064 16068
rect 42116 16056 42122 16108
rect 38933 16031 38991 16037
rect 38933 16028 38945 16031
rect 38120 16000 38945 16028
rect 37921 15991 37979 15997
rect 38933 15997 38945 16000
rect 38979 15997 38991 16031
rect 38933 15991 38991 15997
rect 34974 15920 34980 15972
rect 35032 15960 35038 15972
rect 36998 15960 37004 15972
rect 35032 15932 37004 15960
rect 35032 15920 35038 15932
rect 36998 15920 37004 15932
rect 37056 15920 37062 15972
rect 37936 15960 37964 15991
rect 39482 15988 39488 16040
rect 39540 15988 39546 16040
rect 38102 15960 38108 15972
rect 37936 15932 38108 15960
rect 38102 15920 38108 15932
rect 38160 15920 38166 15972
rect 40052 15960 40080 16056
rect 40218 15988 40224 16040
rect 40276 15988 40282 16040
rect 40494 15988 40500 16040
rect 40552 16028 40558 16040
rect 41049 16031 41107 16037
rect 41049 16028 41061 16031
rect 40552 16000 41061 16028
rect 40552 15988 40558 16000
rect 41049 15997 41061 16000
rect 41095 15997 41107 16031
rect 41049 15991 41107 15997
rect 41509 16031 41567 16037
rect 41509 15997 41521 16031
rect 41555 16028 41567 16031
rect 42242 16028 42248 16040
rect 41555 16000 42248 16028
rect 41555 15997 41567 16000
rect 41509 15991 41567 15997
rect 42242 15988 42248 16000
rect 42300 15988 42306 16040
rect 41693 15963 41751 15969
rect 41693 15960 41705 15963
rect 40052 15932 41705 15960
rect 41693 15929 41705 15932
rect 41739 15929 41751 15963
rect 41693 15923 41751 15929
rect 34992 15892 35020 15920
rect 31404 15864 35020 15892
rect 35250 15852 35256 15904
rect 35308 15892 35314 15904
rect 36538 15892 36544 15904
rect 35308 15864 36544 15892
rect 35308 15852 35314 15864
rect 36538 15852 36544 15864
rect 36596 15852 36602 15904
rect 37274 15852 37280 15904
rect 37332 15852 37338 15904
rect 37550 15852 37556 15904
rect 37608 15892 37614 15904
rect 41417 15895 41475 15901
rect 41417 15892 41429 15895
rect 37608 15864 41429 15892
rect 37608 15852 37614 15864
rect 41417 15861 41429 15864
rect 41463 15861 41475 15895
rect 41417 15855 41475 15861
rect 1104 15802 42504 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 42504 15802
rect 1104 15728 42504 15750
rect 3559 15691 3617 15697
rect 3559 15657 3571 15691
rect 3605 15688 3617 15691
rect 4798 15688 4804 15700
rect 3605 15660 4804 15688
rect 3605 15657 3617 15660
rect 3559 15651 3617 15657
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 5718 15648 5724 15700
rect 5776 15648 5782 15700
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 7653 15691 7711 15697
rect 7653 15688 7665 15691
rect 6512 15660 7665 15688
rect 6512 15648 6518 15660
rect 7653 15657 7665 15660
rect 7699 15657 7711 15691
rect 7653 15651 7711 15657
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 8389 15691 8447 15697
rect 8389 15688 8401 15691
rect 8260 15660 8401 15688
rect 8260 15648 8266 15660
rect 8389 15657 8401 15660
rect 8435 15657 8447 15691
rect 11606 15688 11612 15700
rect 8389 15651 8447 15657
rect 10336 15660 11612 15688
rect 5629 15623 5687 15629
rect 5629 15589 5641 15623
rect 5675 15589 5687 15623
rect 5629 15583 5687 15589
rect 8297 15623 8355 15629
rect 8297 15589 8309 15623
rect 8343 15620 8355 15623
rect 9030 15620 9036 15632
rect 8343 15592 9036 15620
rect 8343 15589 8355 15592
rect 8297 15583 8355 15589
rect 1762 15512 1768 15564
rect 1820 15512 1826 15564
rect 5350 15512 5356 15564
rect 5408 15512 5414 15564
rect 5644 15552 5672 15583
rect 9030 15580 9036 15592
rect 9088 15580 9094 15632
rect 9122 15580 9128 15632
rect 9180 15620 9186 15632
rect 10336 15620 10364 15660
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 11790 15648 11796 15700
rect 11848 15648 11854 15700
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 12253 15691 12311 15697
rect 12253 15688 12265 15691
rect 12032 15660 12265 15688
rect 12032 15648 12038 15660
rect 12253 15657 12265 15660
rect 12299 15657 12311 15691
rect 12253 15651 12311 15657
rect 13814 15648 13820 15700
rect 13872 15648 13878 15700
rect 16761 15691 16819 15697
rect 16761 15657 16773 15691
rect 16807 15688 16819 15691
rect 17494 15688 17500 15700
rect 16807 15660 17500 15688
rect 16807 15657 16819 15660
rect 16761 15651 16819 15657
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 18874 15688 18880 15700
rect 18472 15660 18880 15688
rect 18472 15648 18478 15660
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 18969 15691 19027 15697
rect 18969 15657 18981 15691
rect 19015 15688 19027 15691
rect 19426 15688 19432 15700
rect 19015 15660 19432 15688
rect 19015 15657 19027 15660
rect 18969 15651 19027 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19886 15648 19892 15700
rect 19944 15648 19950 15700
rect 19981 15691 20039 15697
rect 19981 15657 19993 15691
rect 20027 15688 20039 15691
rect 20346 15688 20352 15700
rect 20027 15660 20352 15688
rect 20027 15657 20039 15660
rect 19981 15651 20039 15657
rect 20346 15648 20352 15660
rect 20404 15688 20410 15700
rect 20404 15660 20576 15688
rect 20404 15648 20410 15660
rect 9180 15592 10364 15620
rect 9180 15580 9186 15592
rect 7193 15555 7251 15561
rect 7193 15552 7205 15555
rect 5644 15524 7205 15552
rect 7193 15521 7205 15524
rect 7239 15521 7251 15555
rect 9140 15552 9168 15580
rect 7193 15515 7251 15521
rect 8588 15524 9168 15552
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15484 2191 15487
rect 2222 15484 2228 15496
rect 2179 15456 2228 15484
rect 2179 15453 2191 15456
rect 2133 15447 2191 15453
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 5258 15444 5264 15496
rect 5316 15444 5322 15496
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 7558 15484 7564 15496
rect 7515 15456 7564 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 8202 15484 8208 15496
rect 8159 15456 8208 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 8588 15493 8616 15524
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15453 8355 15487
rect 8297 15447 8355 15453
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 9582 15484 9588 15496
rect 8803 15456 9588 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 3970 15416 3976 15428
rect 3174 15388 3976 15416
rect 3970 15376 3976 15388
rect 4028 15376 4034 15428
rect 6638 15376 6644 15428
rect 6696 15376 6702 15428
rect 7926 15376 7932 15428
rect 7984 15376 7990 15428
rect 8312 15416 8340 15447
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 9692 15484 9720 15592
rect 9769 15555 9827 15561
rect 9769 15521 9781 15555
rect 9815 15552 9827 15555
rect 9950 15552 9956 15564
rect 9815 15524 9956 15552
rect 9815 15521 9827 15524
rect 9769 15515 9827 15521
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 10336 15561 10364 15592
rect 10686 15580 10692 15632
rect 10744 15580 10750 15632
rect 11808 15620 11836 15648
rect 19150 15620 19156 15632
rect 11808 15592 13492 15620
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 9861 15487 9919 15493
rect 9861 15484 9873 15487
rect 9692 15456 9873 15484
rect 9861 15453 9873 15456
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 10042 15444 10048 15496
rect 10100 15444 10106 15496
rect 10873 15487 10931 15493
rect 10873 15453 10885 15487
rect 10919 15484 10931 15487
rect 10919 15456 12434 15484
rect 10919 15453 10931 15456
rect 10873 15447 10931 15453
rect 9953 15419 10011 15425
rect 9953 15416 9965 15419
rect 8312 15388 9965 15416
rect 9953 15385 9965 15388
rect 9999 15385 10011 15419
rect 11118 15419 11176 15425
rect 11118 15416 11130 15419
rect 9953 15379 10011 15385
rect 10796 15388 11130 15416
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 10796 15357 10824 15388
rect 11118 15385 11130 15388
rect 11164 15385 11176 15419
rect 12406 15416 12434 15456
rect 12802 15444 12808 15496
rect 12860 15484 12866 15496
rect 12897 15487 12955 15493
rect 12897 15484 12909 15487
rect 12860 15456 12909 15484
rect 12860 15444 12866 15456
rect 12897 15453 12909 15456
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 12912 15416 12940 15447
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 13044 15456 13093 15484
rect 13044 15444 13050 15456
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 13262 15444 13268 15496
rect 13320 15444 13326 15496
rect 13354 15444 13360 15496
rect 13412 15444 13418 15496
rect 13464 15493 13492 15592
rect 18156 15592 19156 15620
rect 17129 15555 17187 15561
rect 17129 15521 17141 15555
rect 17175 15552 17187 15555
rect 18156 15552 18184 15592
rect 19150 15580 19156 15592
rect 19208 15580 19214 15632
rect 19242 15580 19248 15632
rect 19300 15620 19306 15632
rect 19300 15592 20392 15620
rect 19300 15580 19306 15592
rect 17175 15524 18184 15552
rect 18601 15555 18659 15561
rect 17175 15521 17187 15524
rect 17129 15515 17187 15521
rect 18601 15521 18613 15555
rect 18647 15552 18659 15555
rect 18690 15552 18696 15564
rect 18647 15524 18696 15552
rect 18647 15521 18659 15524
rect 18601 15515 18659 15521
rect 18690 15512 18696 15524
rect 18748 15552 18754 15564
rect 18748 15524 19012 15552
rect 18748 15512 18754 15524
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 13630 15444 13636 15496
rect 13688 15444 13694 15496
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 15252 15456 15393 15484
rect 15252 15444 15258 15456
rect 15381 15453 15393 15456
rect 15427 15484 15439 15487
rect 16853 15487 16911 15493
rect 16853 15484 16865 15487
rect 15427 15456 16865 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 16853 15453 16865 15456
rect 16899 15453 16911 15487
rect 16853 15447 16911 15453
rect 13538 15416 13544 15428
rect 12406 15388 12848 15416
rect 12912 15388 13544 15416
rect 11118 15379 11176 15385
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 8536 15320 9137 15348
rect 8536 15308 8542 15320
rect 9125 15317 9137 15320
rect 9171 15317 9183 15351
rect 9125 15311 9183 15317
rect 10781 15351 10839 15357
rect 10781 15317 10793 15351
rect 10827 15317 10839 15351
rect 10781 15311 10839 15317
rect 12345 15351 12403 15357
rect 12345 15317 12357 15351
rect 12391 15348 12403 15351
rect 12618 15348 12624 15360
rect 12391 15320 12624 15348
rect 12391 15317 12403 15320
rect 12345 15311 12403 15317
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 12820 15348 12848 15388
rect 13538 15376 13544 15388
rect 13596 15376 13602 15428
rect 15648 15419 15706 15425
rect 15648 15385 15660 15419
rect 15694 15416 15706 15419
rect 16666 15416 16672 15428
rect 15694 15388 16672 15416
rect 15694 15385 15706 15388
rect 15648 15379 15706 15385
rect 16666 15376 16672 15388
rect 16724 15376 16730 15428
rect 16868 15416 16896 15447
rect 18230 15444 18236 15496
rect 18288 15444 18294 15496
rect 18782 15444 18788 15496
rect 18840 15444 18846 15496
rect 18984 15484 19012 15524
rect 19058 15512 19064 15564
rect 19116 15512 19122 15564
rect 20364 15493 20392 15592
rect 20548 15552 20576 15660
rect 20806 15648 20812 15700
rect 20864 15648 20870 15700
rect 20898 15648 20904 15700
rect 20956 15688 20962 15700
rect 22281 15691 22339 15697
rect 22281 15688 22293 15691
rect 20956 15660 22293 15688
rect 20956 15648 20962 15660
rect 22281 15657 22293 15660
rect 22327 15657 22339 15691
rect 22281 15651 22339 15657
rect 24397 15691 24455 15697
rect 24397 15657 24409 15691
rect 24443 15688 24455 15691
rect 24443 15660 26924 15688
rect 24443 15657 24455 15660
rect 24397 15651 24455 15657
rect 21085 15623 21143 15629
rect 21085 15589 21097 15623
rect 21131 15620 21143 15623
rect 22186 15620 22192 15632
rect 21131 15592 22192 15620
rect 21131 15589 21143 15592
rect 21085 15583 21143 15589
rect 22186 15580 22192 15592
rect 22244 15620 22250 15632
rect 22244 15592 22416 15620
rect 22244 15580 22250 15592
rect 21177 15555 21235 15561
rect 21177 15552 21189 15555
rect 20548 15524 21189 15552
rect 21177 15521 21189 15524
rect 21223 15521 21235 15555
rect 21177 15515 21235 15521
rect 21358 15512 21364 15564
rect 21416 15552 21422 15564
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21416 15524 22109 15552
rect 21416 15512 21422 15524
rect 21468 15493 21496 15524
rect 22097 15521 22109 15524
rect 22143 15521 22155 15555
rect 22097 15515 22155 15521
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 18984 15456 19349 15484
rect 19337 15453 19349 15456
rect 19383 15484 19395 15487
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 19383 15456 20177 15484
rect 19383 15453 19395 15456
rect 19337 15447 19395 15453
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20354 15487 20412 15493
rect 20354 15453 20366 15487
rect 20400 15453 20412 15487
rect 20993 15487 21051 15493
rect 20993 15484 21005 15487
rect 20354 15447 20412 15453
rect 20640 15456 21005 15484
rect 17034 15416 17040 15428
rect 16868 15388 17040 15416
rect 17034 15376 17040 15388
rect 17092 15416 17098 15428
rect 17402 15416 17408 15428
rect 17092 15388 17408 15416
rect 17092 15376 17098 15388
rect 17402 15376 17408 15388
rect 17460 15376 17466 15428
rect 18966 15376 18972 15428
rect 19024 15416 19030 15428
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 19024 15388 19993 15416
rect 19024 15376 19030 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 20257 15419 20315 15425
rect 20257 15385 20269 15419
rect 20303 15416 20315 15419
rect 20530 15416 20536 15428
rect 20303 15388 20536 15416
rect 20303 15385 20315 15388
rect 20257 15379 20315 15385
rect 20530 15376 20536 15388
rect 20588 15376 20594 15428
rect 14366 15348 14372 15360
rect 12820 15320 14372 15348
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 18874 15308 18880 15360
rect 18932 15348 18938 15360
rect 19886 15348 19892 15360
rect 18932 15320 19892 15348
rect 18932 15308 18938 15320
rect 19886 15308 19892 15320
rect 19944 15348 19950 15360
rect 20438 15348 20444 15360
rect 19944 15320 20444 15348
rect 19944 15308 19950 15320
rect 20438 15308 20444 15320
rect 20496 15348 20502 15360
rect 20640 15348 20668 15456
rect 20993 15453 21005 15456
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21269 15487 21327 15493
rect 21269 15453 21281 15487
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 21453 15487 21511 15493
rect 21453 15453 21465 15487
rect 21499 15484 21511 15487
rect 21499 15456 21533 15484
rect 21499 15453 21511 15456
rect 21453 15447 21511 15453
rect 21284 15416 21312 15447
rect 21818 15444 21824 15496
rect 21876 15493 21882 15496
rect 21876 15487 21909 15493
rect 21897 15453 21909 15487
rect 21876 15447 21909 15453
rect 22005 15487 22063 15493
rect 22005 15453 22017 15487
rect 22051 15484 22063 15487
rect 22278 15484 22284 15496
rect 22051 15456 22284 15484
rect 22051 15453 22063 15456
rect 22005 15447 22063 15453
rect 21876 15444 21882 15447
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 22388 15493 22416 15592
rect 22462 15580 22468 15632
rect 22520 15620 22526 15632
rect 22649 15623 22707 15629
rect 22649 15620 22661 15623
rect 22520 15592 22661 15620
rect 22520 15580 22526 15592
rect 22649 15589 22661 15592
rect 22695 15589 22707 15623
rect 22649 15583 22707 15589
rect 24673 15623 24731 15629
rect 24673 15589 24685 15623
rect 24719 15620 24731 15623
rect 24762 15620 24768 15632
rect 24719 15592 24768 15620
rect 24719 15589 24731 15592
rect 24673 15583 24731 15589
rect 24762 15580 24768 15592
rect 24820 15580 24826 15632
rect 25869 15623 25927 15629
rect 25869 15620 25881 15623
rect 25516 15592 25881 15620
rect 22572 15524 22968 15552
rect 22373 15487 22431 15493
rect 22373 15453 22385 15487
rect 22419 15453 22431 15487
rect 22373 15447 22431 15453
rect 22462 15444 22468 15496
rect 22520 15484 22526 15496
rect 22572 15493 22600 15524
rect 22940 15493 22968 15524
rect 23750 15512 23756 15564
rect 23808 15552 23814 15564
rect 25516 15552 25544 15592
rect 25869 15589 25881 15592
rect 25915 15589 25927 15623
rect 26326 15620 26332 15632
rect 25869 15583 25927 15589
rect 25976 15592 26332 15620
rect 25976 15552 26004 15592
rect 26326 15580 26332 15592
rect 26384 15580 26390 15632
rect 26896 15620 26924 15660
rect 28534 15648 28540 15700
rect 28592 15688 28598 15700
rect 37001 15691 37059 15697
rect 28592 15660 29684 15688
rect 28592 15648 28598 15660
rect 27430 15620 27436 15632
rect 26896 15592 27436 15620
rect 27430 15580 27436 15592
rect 27488 15620 27494 15632
rect 28905 15623 28963 15629
rect 28905 15620 28917 15623
rect 27488 15592 28917 15620
rect 27488 15580 27494 15592
rect 28905 15589 28917 15592
rect 28951 15589 28963 15623
rect 28905 15583 28963 15589
rect 28997 15623 29055 15629
rect 28997 15589 29009 15623
rect 29043 15620 29055 15623
rect 29270 15620 29276 15632
rect 29043 15592 29276 15620
rect 29043 15589 29055 15592
rect 28997 15583 29055 15589
rect 29270 15580 29276 15592
rect 29328 15620 29334 15632
rect 29549 15623 29607 15629
rect 29549 15620 29561 15623
rect 29328 15592 29561 15620
rect 29328 15580 29334 15592
rect 29549 15589 29561 15592
rect 29595 15589 29607 15623
rect 29549 15583 29607 15589
rect 23808 15524 24808 15552
rect 23808 15512 23814 15524
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 22520 15456 22569 15484
rect 22520 15444 22526 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 23109 15487 23167 15493
rect 23109 15453 23121 15487
rect 23155 15484 23167 15487
rect 23658 15484 23664 15496
rect 23155 15456 23664 15484
rect 23155 15453 23167 15456
rect 23109 15447 23167 15453
rect 21836 15416 21864 15444
rect 21284 15388 21864 15416
rect 22756 15416 22784 15447
rect 23124 15416 23152 15447
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 23934 15444 23940 15496
rect 23992 15484 23998 15496
rect 24780 15493 24808 15524
rect 24872 15524 25544 15552
rect 24872 15493 24900 15524
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 23992 15456 24593 15484
rect 23992 15444 23998 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 24857 15487 24915 15493
rect 24857 15453 24869 15487
rect 24903 15453 24915 15487
rect 24857 15447 24915 15453
rect 25038 15444 25044 15496
rect 25096 15444 25102 15496
rect 25516 15493 25544 15524
rect 25792 15524 26004 15552
rect 25792 15493 25820 15524
rect 26050 15512 26056 15564
rect 26108 15552 26114 15564
rect 26510 15552 26516 15564
rect 26108 15524 26516 15552
rect 26108 15512 26114 15524
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 29454 15552 29460 15564
rect 28828 15524 29460 15552
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15453 25559 15487
rect 25501 15447 25559 15453
rect 25685 15487 25743 15493
rect 25685 15453 25697 15487
rect 25731 15453 25743 15487
rect 25685 15447 25743 15453
rect 25777 15487 25835 15493
rect 25777 15453 25789 15487
rect 25823 15453 25835 15487
rect 25777 15447 25835 15453
rect 25954 15487 26012 15493
rect 25954 15453 25966 15487
rect 26000 15453 26012 15487
rect 25954 15447 26012 15453
rect 26145 15487 26203 15493
rect 26145 15453 26157 15487
rect 26191 15484 26203 15487
rect 26789 15487 26847 15493
rect 26789 15484 26801 15487
rect 26191 15456 26801 15484
rect 26191 15453 26203 15456
rect 26145 15447 26203 15453
rect 22756 15388 23152 15416
rect 20496 15320 20668 15348
rect 20496 15308 20502 15320
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 21637 15351 21695 15357
rect 21637 15348 21649 15351
rect 21048 15320 21649 15348
rect 21048 15308 21054 15320
rect 21637 15317 21649 15320
rect 21683 15317 21695 15351
rect 21637 15311 21695 15317
rect 22097 15351 22155 15357
rect 22097 15317 22109 15351
rect 22143 15348 22155 15351
rect 22186 15348 22192 15360
rect 22143 15320 22192 15348
rect 22143 15317 22155 15320
rect 22097 15311 22155 15317
rect 22186 15308 22192 15320
rect 22244 15308 22250 15360
rect 22278 15308 22284 15360
rect 22336 15348 22342 15360
rect 23017 15351 23075 15357
rect 23017 15348 23029 15351
rect 22336 15320 23029 15348
rect 22336 15308 22342 15320
rect 23017 15317 23029 15320
rect 23063 15348 23075 15351
rect 23934 15348 23940 15360
rect 23063 15320 23940 15348
rect 23063 15317 23075 15320
rect 23017 15311 23075 15317
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 25590 15308 25596 15360
rect 25648 15308 25654 15360
rect 25700 15348 25728 15447
rect 25976 15416 26004 15447
rect 26050 15416 26056 15428
rect 25976 15388 26056 15416
rect 26050 15376 26056 15388
rect 26108 15376 26114 15428
rect 26252 15348 26280 15456
rect 26789 15453 26801 15456
rect 26835 15453 26847 15487
rect 26789 15447 26847 15453
rect 26881 15487 26939 15493
rect 26881 15453 26893 15487
rect 26927 15484 26939 15487
rect 26927 15456 27568 15484
rect 26927 15453 26939 15456
rect 26881 15447 26939 15453
rect 26326 15376 26332 15428
rect 26384 15376 26390 15428
rect 26510 15376 26516 15428
rect 26568 15376 26574 15428
rect 27246 15376 27252 15428
rect 27304 15376 27310 15428
rect 27540 15416 27568 15456
rect 27614 15444 27620 15496
rect 27672 15444 27678 15496
rect 28626 15444 28632 15496
rect 28684 15444 28690 15496
rect 28828 15493 28856 15524
rect 29454 15512 29460 15524
rect 29512 15512 29518 15564
rect 28813 15487 28871 15493
rect 28813 15453 28825 15487
rect 28859 15453 28871 15487
rect 28813 15447 28871 15453
rect 29089 15487 29147 15493
rect 29089 15453 29101 15487
rect 29135 15453 29147 15487
rect 29089 15447 29147 15453
rect 29549 15487 29607 15493
rect 29549 15453 29561 15487
rect 29595 15484 29607 15487
rect 29656 15484 29684 15660
rect 37001 15657 37013 15691
rect 37047 15688 37059 15691
rect 37090 15688 37096 15700
rect 37047 15660 37096 15688
rect 37047 15657 37059 15660
rect 37001 15651 37059 15657
rect 37090 15648 37096 15660
rect 37148 15648 37154 15700
rect 37274 15648 37280 15700
rect 37332 15688 37338 15700
rect 37442 15691 37500 15697
rect 37442 15688 37454 15691
rect 37332 15660 37454 15688
rect 37332 15648 37338 15660
rect 37442 15657 37454 15660
rect 37488 15657 37500 15691
rect 37442 15651 37500 15657
rect 38654 15648 38660 15700
rect 38712 15688 38718 15700
rect 41598 15688 41604 15700
rect 38712 15660 41604 15688
rect 38712 15648 38718 15660
rect 41598 15648 41604 15660
rect 41656 15648 41662 15700
rect 38764 15592 40908 15620
rect 31294 15512 31300 15564
rect 31352 15552 31358 15564
rect 31481 15555 31539 15561
rect 31481 15552 31493 15555
rect 31352 15524 31493 15552
rect 31352 15512 31358 15524
rect 31481 15521 31493 15524
rect 31527 15521 31539 15555
rect 31481 15515 31539 15521
rect 31665 15555 31723 15561
rect 31665 15521 31677 15555
rect 31711 15552 31723 15555
rect 33042 15552 33048 15564
rect 31711 15524 33048 15552
rect 31711 15521 31723 15524
rect 31665 15515 31723 15521
rect 33042 15512 33048 15524
rect 33100 15512 33106 15564
rect 35250 15512 35256 15564
rect 35308 15552 35314 15564
rect 37185 15555 37243 15561
rect 37185 15552 37197 15555
rect 35308 15524 37197 15552
rect 35308 15512 35314 15524
rect 37185 15521 37197 15524
rect 37231 15552 37243 15555
rect 37458 15552 37464 15564
rect 37231 15524 37464 15552
rect 37231 15521 37243 15524
rect 37185 15515 37243 15521
rect 37458 15512 37464 15524
rect 37516 15512 37522 15564
rect 38654 15512 38660 15564
rect 38712 15512 38718 15564
rect 29595 15456 29684 15484
rect 29595 15453 29607 15456
rect 29549 15447 29607 15453
rect 27706 15416 27712 15428
rect 27540 15388 27712 15416
rect 27706 15376 27712 15388
rect 27764 15416 27770 15428
rect 29104 15416 29132 15447
rect 29730 15444 29736 15496
rect 29788 15444 29794 15496
rect 31754 15484 31760 15496
rect 31312 15456 31760 15484
rect 27764 15388 29132 15416
rect 29273 15419 29331 15425
rect 27764 15376 27770 15388
rect 29273 15385 29285 15419
rect 29319 15416 29331 15419
rect 31312 15416 31340 15456
rect 31754 15444 31760 15456
rect 31812 15444 31818 15496
rect 31846 15444 31852 15496
rect 31904 15444 31910 15496
rect 38672 15484 38700 15512
rect 38594 15456 38700 15484
rect 29319 15388 31340 15416
rect 31389 15419 31447 15425
rect 29319 15385 29331 15388
rect 29273 15379 29331 15385
rect 31389 15385 31401 15419
rect 31435 15416 31447 15419
rect 32493 15419 32551 15425
rect 32493 15416 32505 15419
rect 31435 15388 32505 15416
rect 31435 15385 31447 15388
rect 31389 15379 31447 15385
rect 32493 15385 32505 15388
rect 32539 15416 32551 15419
rect 32766 15416 32772 15428
rect 32539 15388 32772 15416
rect 32539 15385 32551 15388
rect 32493 15379 32551 15385
rect 32766 15376 32772 15388
rect 32824 15376 32830 15428
rect 35434 15376 35440 15428
rect 35492 15416 35498 15428
rect 35529 15419 35587 15425
rect 35529 15416 35541 15419
rect 35492 15388 35541 15416
rect 35492 15376 35498 15388
rect 35529 15385 35541 15388
rect 35575 15385 35587 15419
rect 36754 15388 36860 15416
rect 35529 15379 35587 15385
rect 25700 15320 26280 15348
rect 26344 15348 26372 15376
rect 26694 15348 26700 15360
rect 26344 15320 26700 15348
rect 26694 15308 26700 15320
rect 26752 15308 26758 15360
rect 26786 15308 26792 15360
rect 26844 15348 26850 15360
rect 27157 15351 27215 15357
rect 27157 15348 27169 15351
rect 26844 15320 27169 15348
rect 26844 15308 26850 15320
rect 27157 15317 27169 15320
rect 27203 15348 27215 15351
rect 27522 15348 27528 15360
rect 27203 15320 27528 15348
rect 27203 15317 27215 15320
rect 27157 15311 27215 15317
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 28350 15308 28356 15360
rect 28408 15348 28414 15360
rect 29730 15348 29736 15360
rect 28408 15320 29736 15348
rect 28408 15308 28414 15320
rect 29730 15308 29736 15320
rect 29788 15308 29794 15360
rect 31018 15308 31024 15360
rect 31076 15308 31082 15360
rect 36538 15308 36544 15360
rect 36596 15348 36602 15360
rect 36832 15348 36860 15388
rect 38764 15348 38792 15592
rect 38933 15555 38991 15561
rect 38933 15521 38945 15555
rect 38979 15552 38991 15555
rect 39482 15552 39488 15564
rect 38979 15524 39488 15552
rect 38979 15521 38991 15524
rect 38933 15515 38991 15521
rect 39482 15512 39488 15524
rect 39540 15512 39546 15564
rect 39850 15512 39856 15564
rect 39908 15552 39914 15564
rect 39908 15524 40172 15552
rect 39908 15512 39914 15524
rect 39114 15444 39120 15496
rect 39172 15444 39178 15496
rect 39574 15444 39580 15496
rect 39632 15444 39638 15496
rect 39022 15376 39028 15428
rect 39080 15416 39086 15428
rect 39868 15416 39896 15512
rect 40034 15444 40040 15496
rect 40092 15444 40098 15496
rect 40144 15493 40172 15524
rect 40129 15487 40187 15493
rect 40129 15453 40141 15487
rect 40175 15453 40187 15487
rect 40129 15447 40187 15453
rect 40402 15444 40408 15496
rect 40460 15444 40466 15496
rect 39080 15388 39896 15416
rect 40221 15419 40279 15425
rect 39080 15376 39086 15388
rect 40221 15385 40233 15419
rect 40267 15416 40279 15419
rect 40773 15419 40831 15425
rect 40773 15416 40785 15419
rect 40267 15388 40785 15416
rect 40267 15385 40279 15388
rect 40221 15379 40279 15385
rect 40773 15385 40785 15388
rect 40819 15385 40831 15419
rect 40773 15379 40831 15385
rect 36596 15320 38792 15348
rect 36596 15308 36602 15320
rect 39206 15308 39212 15360
rect 39264 15308 39270 15360
rect 39298 15308 39304 15360
rect 39356 15308 39362 15360
rect 39853 15351 39911 15357
rect 39853 15317 39865 15351
rect 39899 15348 39911 15351
rect 40034 15348 40040 15360
rect 39899 15320 40040 15348
rect 39899 15317 39911 15320
rect 39853 15311 39911 15317
rect 40034 15308 40040 15320
rect 40092 15308 40098 15360
rect 40880 15348 40908 15592
rect 41414 15444 41420 15496
rect 41472 15444 41478 15496
rect 41782 15376 41788 15428
rect 41840 15416 41846 15428
rect 41877 15419 41935 15425
rect 41877 15416 41889 15419
rect 41840 15388 41889 15416
rect 41840 15376 41846 15388
rect 41877 15385 41889 15388
rect 41923 15385 41935 15419
rect 41877 15379 41935 15385
rect 41800 15348 41828 15376
rect 40880 15320 41828 15348
rect 1104 15258 42504 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 42504 15258
rect 1104 15184 42504 15206
rect 4479 15147 4537 15153
rect 4479 15113 4491 15147
rect 4525 15144 4537 15147
rect 4614 15144 4620 15156
rect 4525 15116 4620 15144
rect 4525 15113 4537 15116
rect 4479 15107 4537 15113
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 5166 15144 5172 15156
rect 4755 15116 5172 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 5166 15104 5172 15116
rect 5224 15104 5230 15156
rect 5429 15147 5487 15153
rect 5429 15113 5441 15147
rect 5475 15144 5487 15147
rect 5534 15144 5540 15156
rect 5475 15116 5540 15144
rect 5475 15113 5487 15116
rect 5429 15107 5487 15113
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 7098 15144 7104 15156
rect 6687 15116 7104 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 7098 15104 7104 15116
rect 7156 15144 7162 15156
rect 7926 15144 7932 15156
rect 7156 15116 7932 15144
rect 7156 15104 7162 15116
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10100 15116 10149 15144
rect 10100 15104 10106 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 12989 15147 13047 15153
rect 12989 15113 13001 15147
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 3970 15036 3976 15088
rect 4028 15036 4034 15088
rect 5258 15036 5264 15088
rect 5316 15076 5322 15088
rect 5629 15079 5687 15085
rect 5629 15076 5641 15079
rect 5316 15048 5641 15076
rect 5316 15036 5322 15048
rect 5629 15045 5641 15048
rect 5675 15076 5687 15079
rect 5718 15076 5724 15088
rect 5675 15048 5724 15076
rect 5675 15045 5687 15048
rect 5629 15039 5687 15045
rect 5718 15036 5724 15048
rect 5776 15036 5782 15088
rect 8294 15076 8300 15088
rect 6840 15048 8300 15076
rect 6840 15020 6868 15048
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 13004 15076 13032 15107
rect 13538 15104 13544 15156
rect 13596 15104 13602 15156
rect 16482 15104 16488 15156
rect 16540 15104 16546 15156
rect 18138 15104 18144 15156
rect 18196 15104 18202 15156
rect 19058 15104 19064 15156
rect 19116 15104 19122 15156
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 19702 15144 19708 15156
rect 19392 15116 19708 15144
rect 19392 15104 19398 15116
rect 19702 15104 19708 15116
rect 19760 15144 19766 15156
rect 19797 15147 19855 15153
rect 19797 15144 19809 15147
rect 19760 15116 19809 15144
rect 19760 15104 19766 15116
rect 19797 15113 19809 15116
rect 19843 15113 19855 15147
rect 19797 15107 19855 15113
rect 19978 15104 19984 15156
rect 20036 15144 20042 15156
rect 20257 15147 20315 15153
rect 20257 15144 20269 15147
rect 20036 15116 20269 15144
rect 20036 15104 20042 15116
rect 20257 15113 20269 15116
rect 20303 15113 20315 15147
rect 20257 15107 20315 15113
rect 20717 15147 20775 15153
rect 20717 15113 20729 15147
rect 20763 15144 20775 15147
rect 20898 15144 20904 15156
rect 20763 15116 20904 15144
rect 20763 15113 20775 15116
rect 20717 15107 20775 15113
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 26513 15147 26571 15153
rect 26513 15144 26525 15147
rect 24688 15116 26525 15144
rect 14654 15079 14712 15085
rect 14654 15076 14666 15079
rect 13004 15048 14666 15076
rect 14654 15045 14666 15048
rect 14700 15045 14712 15079
rect 19076 15076 19104 15104
rect 19076 15048 20024 15076
rect 14654 15039 14712 15045
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 15008 4951 15011
rect 5902 15008 5908 15020
rect 4939 14980 5908 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 2682 14900 2688 14952
rect 2740 14900 2746 14952
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3786 14940 3792 14952
rect 3099 14912 3792 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 3786 14900 3792 14912
rect 3844 14900 3850 14952
rect 4632 14940 4660 14971
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 6089 15011 6147 15017
rect 6089 14977 6101 15011
rect 6135 14977 6147 15011
rect 6089 14971 6147 14977
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 4632 14912 5304 14940
rect 5276 14816 5304 14912
rect 5810 14900 5816 14952
rect 5868 14940 5874 14952
rect 6104 14940 6132 14971
rect 5868 14912 6132 14940
rect 5868 14900 5874 14912
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 5905 14875 5963 14881
rect 5905 14872 5917 14875
rect 5776 14844 5917 14872
rect 5776 14832 5782 14844
rect 5905 14841 5917 14844
rect 5951 14841 5963 14875
rect 6564 14872 6592 14971
rect 6822 14968 6828 15020
rect 6880 14968 6886 15020
rect 8205 15011 8263 15017
rect 8205 14977 8217 15011
rect 8251 15008 8263 15011
rect 8478 15008 8484 15020
rect 8251 14980 8484 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8921 15011 8979 15017
rect 8921 15008 8933 15011
rect 8588 14980 8933 15008
rect 7558 14900 7564 14952
rect 7616 14900 7622 14952
rect 8110 14900 8116 14952
rect 8168 14900 8174 14952
rect 8588 14949 8616 14980
rect 8921 14977 8933 14980
rect 8967 14977 8979 15011
rect 8921 14971 8979 14977
rect 12618 14968 12624 15020
rect 12676 14968 12682 15020
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 15105 15011 15163 15017
rect 15105 15008 15117 15011
rect 14967 14980 15117 15008
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 15105 14977 15117 14980
rect 15151 15008 15163 15011
rect 15194 15008 15200 15020
rect 15151 14980 15200 15008
rect 15151 14977 15163 14980
rect 15105 14971 15163 14977
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 15378 15017 15384 15020
rect 15372 15008 15384 15017
rect 15339 14980 15384 15008
rect 15372 14971 15384 14980
rect 15378 14968 15384 14971
rect 15436 14968 15442 15020
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16632 14980 16681 15008
rect 16632 14968 16638 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18049 15011 18107 15017
rect 18049 15008 18061 15011
rect 18012 14980 18061 15008
rect 18012 14968 18018 14980
rect 18049 14977 18061 14980
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 18874 14968 18880 15020
rect 18932 14968 18938 15020
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 15008 19119 15011
rect 19107 14980 19840 15008
rect 19107 14977 19119 14980
rect 19061 14971 19119 14977
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 8665 14943 8723 14949
rect 8665 14909 8677 14943
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 7576 14872 7604 14900
rect 8680 14872 8708 14903
rect 10318 14900 10324 14952
rect 10376 14940 10382 14952
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 10376 14912 10701 14940
rect 10376 14900 10382 14912
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14940 12771 14943
rect 12986 14940 12992 14952
rect 12759 14912 12992 14940
rect 12759 14909 12771 14912
rect 12713 14903 12771 14909
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 17034 14900 17040 14952
rect 17092 14940 17098 14952
rect 17405 14943 17463 14949
rect 17405 14940 17417 14943
rect 17092 14912 17417 14940
rect 17092 14900 17098 14912
rect 17405 14909 17417 14912
rect 17451 14909 17463 14943
rect 17405 14903 17463 14909
rect 18322 14900 18328 14952
rect 18380 14900 18386 14952
rect 18414 14900 18420 14952
rect 18472 14940 18478 14952
rect 19153 14943 19211 14949
rect 19153 14940 19165 14943
rect 18472 14912 19165 14940
rect 18472 14900 18478 14912
rect 19153 14909 19165 14912
rect 19199 14909 19211 14943
rect 19812 14940 19840 14980
rect 19886 14968 19892 15020
rect 19944 14968 19950 15020
rect 19996 15017 20024 15048
rect 20346 15036 20352 15088
rect 20404 15036 20410 15088
rect 20438 15036 20444 15088
rect 20496 15076 20502 15088
rect 20533 15079 20591 15085
rect 20533 15076 20545 15079
rect 20496 15048 20545 15076
rect 20496 15036 20502 15048
rect 20533 15045 20545 15048
rect 20579 15045 20591 15079
rect 20533 15039 20591 15045
rect 20622 15036 20628 15088
rect 20680 15076 20686 15088
rect 22373 15079 22431 15085
rect 22373 15076 22385 15079
rect 20680 15048 22385 15076
rect 20680 15036 20686 15048
rect 22373 15045 22385 15048
rect 22419 15076 22431 15079
rect 22830 15076 22836 15088
rect 22419 15048 22836 15076
rect 22419 15045 22431 15048
rect 22373 15039 22431 15045
rect 22830 15036 22836 15048
rect 22888 15036 22894 15088
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 22094 14968 22100 15020
rect 22152 14968 22158 15020
rect 22278 14968 22284 15020
rect 22336 14968 22342 15020
rect 24688 15017 24716 15116
rect 26513 15113 26525 15116
rect 26559 15113 26571 15147
rect 26513 15107 26571 15113
rect 29086 15104 29092 15156
rect 29144 15144 29150 15156
rect 29454 15144 29460 15156
rect 29144 15116 29460 15144
rect 29144 15104 29150 15116
rect 29454 15104 29460 15116
rect 29512 15144 29518 15156
rect 31662 15144 31668 15156
rect 29512 15116 31668 15144
rect 29512 15104 29518 15116
rect 31662 15104 31668 15116
rect 31720 15104 31726 15156
rect 31846 15104 31852 15156
rect 31904 15104 31910 15156
rect 32766 15104 32772 15156
rect 32824 15104 32830 15156
rect 34348 15116 35388 15144
rect 24765 15079 24823 15085
rect 24765 15045 24777 15079
rect 24811 15076 24823 15079
rect 26053 15079 26111 15085
rect 26053 15076 26065 15079
rect 24811 15048 26065 15076
rect 24811 15045 24823 15048
rect 24765 15039 24823 15045
rect 26053 15045 26065 15048
rect 26099 15045 26111 15079
rect 26053 15039 26111 15045
rect 26234 15036 26240 15088
rect 26292 15076 26298 15088
rect 26292 15048 26556 15076
rect 26292 15036 26298 15048
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 24673 15011 24731 15017
rect 24673 14977 24685 15011
rect 24719 14977 24731 15011
rect 24673 14971 24731 14977
rect 24857 15011 24915 15017
rect 24857 14977 24869 15011
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 24995 15011 25053 15017
rect 24995 14977 25007 15011
rect 25041 15008 25053 15011
rect 25866 15008 25872 15020
rect 25041 14980 25872 15008
rect 25041 14977 25053 14980
rect 24995 14971 25053 14977
rect 20438 14940 20444 14952
rect 19812 14912 20444 14940
rect 19153 14903 19211 14909
rect 20438 14900 20444 14912
rect 20496 14900 20502 14952
rect 21085 14943 21143 14949
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 22186 14940 22192 14952
rect 21131 14912 22192 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 12342 14872 12348 14884
rect 6564 14844 7512 14872
rect 7576 14844 8708 14872
rect 9968 14844 12348 14872
rect 5905 14835 5963 14841
rect 4890 14764 4896 14816
rect 4948 14764 4954 14816
rect 5258 14764 5264 14816
rect 5316 14764 5322 14816
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 6270 14804 6276 14816
rect 5500 14776 6276 14804
rect 5500 14764 5506 14776
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 7484 14804 7512 14844
rect 9968 14804 9996 14844
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 18782 14832 18788 14884
rect 18840 14872 18846 14884
rect 18840 14844 19932 14872
rect 18840 14832 18846 14844
rect 7484 14776 9996 14804
rect 10042 14764 10048 14816
rect 10100 14764 10106 14816
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 16264 14776 17693 14804
rect 16264 14764 16270 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 17681 14767 17739 14773
rect 18874 14764 18880 14816
rect 18932 14804 18938 14816
rect 19242 14804 19248 14816
rect 18932 14776 19248 14804
rect 18932 14764 18938 14776
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 19904 14813 19932 14844
rect 21634 14832 21640 14884
rect 21692 14872 21698 14884
rect 22480 14872 22508 14971
rect 24486 14900 24492 14952
rect 24544 14940 24550 14952
rect 24872 14940 24900 14971
rect 25866 14968 25872 14980
rect 25924 14968 25930 15020
rect 26418 14968 26424 15020
rect 26476 14968 26482 15020
rect 26528 15017 26556 15048
rect 27614 15036 27620 15088
rect 27672 15076 27678 15088
rect 28169 15079 28227 15085
rect 28169 15076 28181 15079
rect 27672 15048 28181 15076
rect 27672 15036 27678 15048
rect 28169 15045 28181 15048
rect 28215 15076 28227 15079
rect 30736 15079 30794 15085
rect 28215 15048 30512 15076
rect 28215 15045 28227 15048
rect 28169 15039 28227 15045
rect 26513 15011 26571 15017
rect 26513 14977 26525 15011
rect 26559 14977 26571 15011
rect 26513 14971 26571 14977
rect 26697 15011 26755 15017
rect 26697 14977 26709 15011
rect 26743 14977 26755 15011
rect 26697 14971 26755 14977
rect 27249 15011 27307 15017
rect 27249 14977 27261 15011
rect 27295 14977 27307 15011
rect 27249 14971 27307 14977
rect 24544 14912 24900 14940
rect 24544 14900 24550 14912
rect 24504 14872 24532 14900
rect 21692 14844 22508 14872
rect 22572 14844 24532 14872
rect 24872 14872 24900 14912
rect 25133 14943 25191 14949
rect 25133 14909 25145 14943
rect 25179 14940 25191 14943
rect 25314 14940 25320 14952
rect 25179 14912 25320 14940
rect 25179 14909 25191 14912
rect 25133 14903 25191 14909
rect 25314 14900 25320 14912
rect 25372 14900 25378 14952
rect 25409 14943 25467 14949
rect 25409 14909 25421 14943
rect 25455 14940 25467 14943
rect 25590 14940 25596 14952
rect 25455 14912 25596 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 25590 14900 25596 14912
rect 25648 14900 25654 14952
rect 26436 14940 26464 14968
rect 26712 14940 26740 14971
rect 26436 14912 26740 14940
rect 27264 14940 27292 14971
rect 27430 14968 27436 15020
rect 27488 14968 27494 15020
rect 28629 15011 28687 15017
rect 28629 14977 28641 15011
rect 28675 15008 28687 15011
rect 28810 15008 28816 15020
rect 28675 14980 28816 15008
rect 28675 14977 28687 14980
rect 28629 14971 28687 14977
rect 28810 14968 28816 14980
rect 28868 14968 28874 15020
rect 29086 14968 29092 15020
rect 29144 14968 29150 15020
rect 29273 15011 29331 15017
rect 29273 14977 29285 15011
rect 29319 14977 29331 15011
rect 29273 14971 29331 14977
rect 28166 14940 28172 14952
rect 27264 14912 28172 14940
rect 28166 14900 28172 14912
rect 28224 14900 28230 14952
rect 28718 14900 28724 14952
rect 28776 14900 28782 14952
rect 26418 14872 26424 14884
rect 24872 14844 26424 14872
rect 21692 14832 21698 14844
rect 19889 14807 19947 14813
rect 19889 14773 19901 14807
rect 19935 14773 19947 14807
rect 19889 14767 19947 14773
rect 21269 14807 21327 14813
rect 21269 14773 21281 14807
rect 21315 14804 21327 14807
rect 21450 14804 21456 14816
rect 21315 14776 21456 14804
rect 21315 14773 21327 14776
rect 21269 14767 21327 14773
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 21726 14764 21732 14816
rect 21784 14804 21790 14816
rect 22572 14804 22600 14844
rect 26418 14832 26424 14844
rect 26476 14832 26482 14884
rect 26786 14832 26792 14884
rect 26844 14872 26850 14884
rect 28534 14872 28540 14884
rect 26844 14844 28540 14872
rect 26844 14832 26850 14844
rect 28534 14832 28540 14844
rect 28592 14832 28598 14884
rect 28997 14875 29055 14881
rect 28997 14841 29009 14875
rect 29043 14872 29055 14875
rect 29288 14872 29316 14971
rect 29362 14968 29368 15020
rect 29420 14968 29426 15020
rect 30484 15017 30512 15048
rect 30736 15045 30748 15079
rect 30782 15076 30794 15079
rect 31018 15076 31024 15088
rect 30782 15048 31024 15076
rect 30782 15045 30794 15048
rect 30736 15039 30794 15045
rect 31018 15036 31024 15048
rect 31076 15036 31082 15088
rect 34348 15076 34376 15116
rect 31726 15048 34376 15076
rect 29457 15011 29515 15017
rect 29457 14977 29469 15011
rect 29503 15008 29515 15011
rect 30469 15011 30527 15017
rect 29503 14980 30420 15008
rect 29503 14977 29515 14980
rect 29457 14971 29515 14977
rect 29380 14940 29408 14968
rect 29733 14943 29791 14949
rect 29733 14940 29745 14943
rect 29380 14912 29745 14940
rect 29733 14909 29745 14912
rect 29779 14909 29791 14943
rect 29733 14903 29791 14909
rect 30285 14943 30343 14949
rect 30285 14909 30297 14943
rect 30331 14909 30343 14943
rect 30392 14940 30420 14980
rect 30469 14977 30481 15011
rect 30515 14977 30527 15011
rect 31726 15008 31754 15048
rect 34422 15036 34428 15088
rect 34480 15076 34486 15088
rect 35253 15079 35311 15085
rect 35253 15076 35265 15079
rect 34480 15048 35265 15076
rect 34480 15036 34486 15048
rect 35253 15045 35265 15048
rect 35299 15045 35311 15079
rect 35253 15039 35311 15045
rect 30469 14971 30527 14977
rect 30576 14980 31754 15008
rect 32677 15011 32735 15017
rect 30576 14940 30604 14980
rect 32677 14977 32689 15011
rect 32723 15008 32735 15011
rect 33229 15011 33287 15017
rect 33229 15008 33241 15011
rect 32723 14980 33241 15008
rect 32723 14977 32735 14980
rect 32677 14971 32735 14977
rect 33229 14977 33241 14980
rect 33275 14977 33287 15011
rect 33229 14971 33287 14977
rect 34057 15011 34115 15017
rect 34057 14977 34069 15011
rect 34103 14977 34115 15011
rect 34057 14971 34115 14977
rect 34241 15011 34299 15017
rect 34241 14977 34253 15011
rect 34287 15008 34299 15011
rect 34514 15008 34520 15020
rect 34287 14980 34520 15008
rect 34287 14977 34299 14980
rect 34241 14971 34299 14977
rect 30392 14912 30604 14940
rect 32953 14943 33011 14949
rect 30285 14903 30343 14909
rect 32953 14909 32965 14943
rect 32999 14940 33011 14943
rect 33134 14940 33140 14952
rect 32999 14912 33140 14940
rect 32999 14909 33011 14912
rect 32953 14903 33011 14909
rect 29043 14844 29316 14872
rect 29641 14875 29699 14881
rect 29043 14841 29055 14844
rect 28997 14835 29055 14841
rect 29641 14841 29653 14875
rect 29687 14872 29699 14875
rect 29822 14872 29828 14884
rect 29687 14844 29828 14872
rect 29687 14841 29699 14844
rect 29641 14835 29699 14841
rect 29822 14832 29828 14844
rect 29880 14832 29886 14884
rect 30300 14872 30328 14903
rect 33134 14900 33140 14912
rect 33192 14900 33198 14952
rect 33870 14900 33876 14952
rect 33928 14900 33934 14952
rect 30466 14872 30472 14884
rect 30300 14844 30472 14872
rect 30466 14832 30472 14844
rect 30524 14832 30530 14884
rect 31570 14832 31576 14884
rect 31628 14872 31634 14884
rect 34072 14872 34100 14971
rect 34514 14968 34520 14980
rect 34572 14968 34578 15020
rect 35360 15017 35388 15116
rect 35434 15104 35440 15156
rect 35492 15144 35498 15156
rect 35989 15147 36047 15153
rect 35989 15144 36001 15147
rect 35492 15116 36001 15144
rect 35492 15104 35498 15116
rect 35989 15113 36001 15116
rect 36035 15113 36047 15147
rect 35989 15107 36047 15113
rect 36357 15147 36415 15153
rect 36357 15113 36369 15147
rect 36403 15144 36415 15147
rect 37090 15144 37096 15156
rect 36403 15116 37096 15144
rect 36403 15113 36415 15116
rect 36357 15107 36415 15113
rect 37090 15104 37096 15116
rect 37148 15104 37154 15156
rect 37458 15104 37464 15156
rect 37516 15144 37522 15156
rect 37516 15116 40172 15144
rect 37516 15104 37522 15116
rect 38010 15076 38016 15088
rect 37292 15048 38016 15076
rect 37292 15020 37320 15048
rect 38010 15036 38016 15048
rect 38068 15036 38074 15088
rect 38746 15036 38752 15088
rect 38804 15036 38810 15088
rect 39206 15036 39212 15088
rect 39264 15076 39270 15088
rect 39850 15076 39856 15088
rect 39264 15048 39856 15076
rect 39264 15036 39270 15048
rect 39850 15036 39856 15048
rect 39908 15036 39914 15088
rect 34977 15011 35035 15017
rect 34977 14977 34989 15011
rect 35023 14977 35035 15011
rect 34977 14971 35035 14977
rect 35161 15011 35219 15017
rect 35161 14977 35173 15011
rect 35207 14977 35219 15011
rect 35161 14971 35219 14977
rect 35345 15011 35403 15017
rect 35345 14977 35357 15011
rect 35391 15008 35403 15011
rect 37274 15008 37280 15020
rect 35391 14980 37280 15008
rect 35391 14977 35403 14980
rect 35345 14971 35403 14977
rect 31628 14844 34100 14872
rect 34992 14872 35020 14971
rect 35176 14940 35204 14971
rect 37274 14968 37280 14980
rect 37332 14968 37338 15020
rect 37458 14968 37464 15020
rect 37516 14968 37522 15020
rect 40144 15017 40172 15116
rect 41414 15104 41420 15156
rect 41472 15144 41478 15156
rect 41877 15147 41935 15153
rect 41877 15144 41889 15147
rect 41472 15116 41889 15144
rect 41472 15104 41478 15116
rect 41877 15113 41889 15116
rect 41923 15113 41935 15147
rect 41877 15107 41935 15113
rect 40129 15011 40187 15017
rect 40129 14977 40141 15011
rect 40175 14977 40187 15011
rect 41538 14980 41644 15008
rect 40129 14971 40187 14977
rect 41616 14952 41644 14980
rect 35434 14940 35440 14952
rect 35176 14912 35440 14940
rect 35434 14900 35440 14912
rect 35492 14900 35498 14952
rect 36449 14943 36507 14949
rect 36449 14909 36461 14943
rect 36495 14909 36507 14943
rect 36449 14903 36507 14909
rect 35342 14872 35348 14884
rect 34992 14844 35348 14872
rect 31628 14832 31634 14844
rect 21784 14776 22600 14804
rect 22649 14807 22707 14813
rect 21784 14764 21790 14776
rect 22649 14773 22661 14807
rect 22695 14804 22707 14807
rect 23106 14804 23112 14816
rect 22695 14776 23112 14804
rect 22695 14773 22707 14776
rect 22649 14767 22707 14773
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 24118 14764 24124 14816
rect 24176 14804 24182 14816
rect 24489 14807 24547 14813
rect 24489 14804 24501 14807
rect 24176 14776 24501 14804
rect 24176 14764 24182 14776
rect 24489 14773 24501 14776
rect 24535 14773 24547 14807
rect 24489 14767 24547 14773
rect 25866 14764 25872 14816
rect 25924 14804 25930 14816
rect 25961 14807 26019 14813
rect 25961 14804 25973 14807
rect 25924 14776 25973 14804
rect 25924 14764 25930 14776
rect 25961 14773 25973 14776
rect 26007 14773 26019 14807
rect 25961 14767 26019 14773
rect 26234 14764 26240 14816
rect 26292 14804 26298 14816
rect 27157 14807 27215 14813
rect 27157 14804 27169 14807
rect 26292 14776 27169 14804
rect 26292 14764 26298 14776
rect 27157 14773 27169 14776
rect 27203 14804 27215 14807
rect 27246 14804 27252 14816
rect 27203 14776 27252 14804
rect 27203 14773 27215 14776
rect 27157 14767 27215 14773
rect 27246 14764 27252 14776
rect 27304 14764 27310 14816
rect 32214 14764 32220 14816
rect 32272 14804 32278 14816
rect 32309 14807 32367 14813
rect 32309 14804 32321 14807
rect 32272 14776 32321 14804
rect 32272 14764 32278 14776
rect 32309 14773 32321 14776
rect 32355 14773 32367 14807
rect 32309 14767 32367 14773
rect 34054 14764 34060 14816
rect 34112 14804 34118 14816
rect 34992 14804 35020 14844
rect 35342 14832 35348 14844
rect 35400 14832 35406 14884
rect 36464 14872 36492 14903
rect 36538 14900 36544 14952
rect 36596 14900 36602 14952
rect 37734 14900 37740 14952
rect 37792 14900 37798 14952
rect 39209 14943 39267 14949
rect 39209 14909 39221 14943
rect 39255 14940 39267 14943
rect 39853 14943 39911 14949
rect 39853 14940 39865 14943
rect 39255 14912 39865 14940
rect 39255 14909 39267 14912
rect 39209 14903 39267 14909
rect 39853 14909 39865 14912
rect 39899 14909 39911 14943
rect 39853 14903 39911 14909
rect 40405 14943 40463 14949
rect 40405 14909 40417 14943
rect 40451 14940 40463 14943
rect 40862 14940 40868 14952
rect 40451 14912 40868 14940
rect 40451 14909 40463 14912
rect 40405 14903 40463 14909
rect 39868 14872 39896 14903
rect 40862 14900 40868 14912
rect 40920 14900 40926 14952
rect 41598 14900 41604 14952
rect 41656 14900 41662 14952
rect 40126 14872 40132 14884
rect 36464 14844 37596 14872
rect 39868 14844 40132 14872
rect 34112 14776 35020 14804
rect 35529 14807 35587 14813
rect 34112 14764 34118 14776
rect 35529 14773 35541 14807
rect 35575 14804 35587 14807
rect 36446 14804 36452 14816
rect 35575 14776 36452 14804
rect 35575 14773 35587 14776
rect 35529 14767 35587 14773
rect 36446 14764 36452 14776
rect 36504 14764 36510 14816
rect 37568 14804 37596 14844
rect 40126 14832 40132 14844
rect 40184 14832 40190 14884
rect 38470 14804 38476 14816
rect 37568 14776 38476 14804
rect 38470 14764 38476 14776
rect 38528 14804 38534 14816
rect 39301 14807 39359 14813
rect 39301 14804 39313 14807
rect 38528 14776 39313 14804
rect 38528 14764 38534 14776
rect 39301 14773 39313 14776
rect 39347 14773 39359 14807
rect 39301 14767 39359 14773
rect 1104 14714 42504 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 42504 14714
rect 1104 14640 42504 14662
rect 3786 14560 3792 14612
rect 3844 14560 3850 14612
rect 4890 14560 4896 14612
rect 4948 14600 4954 14612
rect 5058 14603 5116 14609
rect 5058 14600 5070 14603
rect 4948 14572 5070 14600
rect 4948 14560 4954 14572
rect 5058 14569 5070 14572
rect 5104 14569 5116 14603
rect 5058 14563 5116 14569
rect 10318 14560 10324 14612
rect 10376 14560 10382 14612
rect 17954 14560 17960 14612
rect 18012 14560 18018 14612
rect 21913 14603 21971 14609
rect 21913 14569 21925 14603
rect 21959 14600 21971 14603
rect 22370 14600 22376 14612
rect 21959 14572 22376 14600
rect 21959 14569 21971 14572
rect 21913 14563 21971 14569
rect 22370 14560 22376 14572
rect 22428 14560 22434 14612
rect 26881 14603 26939 14609
rect 26881 14569 26893 14603
rect 26927 14600 26939 14603
rect 28626 14600 28632 14612
rect 26927 14572 28632 14600
rect 26927 14569 26939 14572
rect 26881 14563 26939 14569
rect 28626 14560 28632 14572
rect 28684 14560 28690 14612
rect 37734 14560 37740 14612
rect 37792 14600 37798 14612
rect 38013 14603 38071 14609
rect 38013 14600 38025 14603
rect 37792 14572 38025 14600
rect 37792 14560 37798 14572
rect 38013 14569 38025 14572
rect 38059 14569 38071 14603
rect 38013 14563 38071 14569
rect 39574 14560 39580 14612
rect 39632 14560 39638 14612
rect 40862 14560 40868 14612
rect 40920 14560 40926 14612
rect 41782 14560 41788 14612
rect 41840 14560 41846 14612
rect 18322 14492 18328 14544
rect 18380 14532 18386 14544
rect 19426 14532 19432 14544
rect 18380 14504 19432 14532
rect 18380 14492 18386 14504
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 20254 14492 20260 14544
rect 20312 14532 20318 14544
rect 21726 14532 21732 14544
rect 20312 14504 21732 14532
rect 20312 14492 20318 14504
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2682 14464 2688 14476
rect 1443 14436 2688 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2682 14424 2688 14436
rect 2740 14464 2746 14476
rect 4801 14467 4859 14473
rect 4801 14464 4813 14467
rect 2740 14436 4813 14464
rect 2740 14424 2746 14436
rect 4801 14433 4813 14436
rect 4847 14464 4859 14467
rect 7558 14464 7564 14476
rect 4847 14436 7564 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 6932 14405 6960 14436
rect 7558 14424 7564 14436
rect 7616 14464 7622 14476
rect 8294 14464 8300 14476
rect 7616 14436 8300 14464
rect 7616 14424 7622 14436
rect 8294 14424 8300 14436
rect 8352 14464 8358 14476
rect 8941 14467 8999 14473
rect 8941 14464 8953 14467
rect 8352 14436 8953 14464
rect 8352 14424 8358 14436
rect 8941 14433 8953 14436
rect 8987 14433 8999 14467
rect 8941 14427 8999 14433
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 12158 14464 12164 14476
rect 10551 14436 12164 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 15933 14467 15991 14473
rect 15933 14433 15945 14467
rect 15979 14464 15991 14467
rect 16942 14464 16948 14476
rect 15979 14436 16948 14464
rect 15979 14433 15991 14436
rect 15933 14427 15991 14433
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17681 14467 17739 14473
rect 17681 14433 17693 14467
rect 17727 14464 17739 14467
rect 20530 14464 20536 14476
rect 17727 14436 18644 14464
rect 17727 14433 17739 14436
rect 17681 14427 17739 14433
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1728 14368 1777 14396
rect 1728 14356 1734 14368
rect 1765 14365 1777 14368
rect 1811 14365 1823 14399
rect 1765 14359 1823 14365
rect 3191 14399 3249 14405
rect 3191 14365 3203 14399
rect 3237 14396 3249 14399
rect 4341 14399 4399 14405
rect 4341 14396 4353 14399
rect 3237 14368 4353 14396
rect 3237 14365 3249 14368
rect 3191 14359 3249 14365
rect 4341 14365 4353 14368
rect 4387 14365 4399 14399
rect 4341 14359 4399 14365
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 9030 14356 9036 14408
rect 9088 14396 9094 14408
rect 9197 14399 9255 14405
rect 9197 14396 9209 14399
rect 9088 14368 9209 14396
rect 9088 14356 9094 14368
rect 9197 14365 9209 14368
rect 9243 14365 9255 14399
rect 9197 14359 9255 14365
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14396 10839 14399
rect 11974 14396 11980 14408
rect 10827 14368 11980 14396
rect 10827 14365 10839 14368
rect 10781 14359 10839 14365
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 18616 14405 18644 14436
rect 18892 14436 20536 14464
rect 18601 14399 18659 14405
rect 18601 14365 18613 14399
rect 18647 14396 18659 14399
rect 18693 14399 18751 14405
rect 18693 14396 18705 14399
rect 18647 14368 18705 14396
rect 18647 14365 18659 14368
rect 18601 14359 18659 14365
rect 18693 14365 18705 14368
rect 18739 14396 18751 14399
rect 18782 14396 18788 14408
rect 18739 14368 18788 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 18892 14405 18920 14436
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14365 18935 14399
rect 18877 14359 18935 14365
rect 19061 14399 19119 14405
rect 19061 14365 19073 14399
rect 19107 14396 19119 14399
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 19107 14368 19441 14396
rect 19107 14365 19119 14368
rect 19061 14359 19119 14365
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19702 14356 19708 14408
rect 19760 14405 19766 14408
rect 19760 14399 19789 14405
rect 19777 14365 19789 14399
rect 19760 14359 19789 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20714 14396 20720 14408
rect 19935 14368 20720 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 19760 14356 19766 14359
rect 20714 14356 20720 14368
rect 20772 14396 20778 14408
rect 21266 14396 21272 14408
rect 20772 14368 21272 14396
rect 20772 14356 20778 14368
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 21652 14405 21680 14504
rect 21726 14492 21732 14504
rect 21784 14492 21790 14544
rect 34517 14535 34575 14541
rect 34517 14501 34529 14535
rect 34563 14532 34575 14535
rect 35434 14532 35440 14544
rect 34563 14504 35440 14532
rect 34563 14501 34575 14504
rect 34517 14495 34575 14501
rect 35434 14492 35440 14504
rect 35492 14492 35498 14544
rect 39853 14535 39911 14541
rect 39853 14532 39865 14535
rect 39040 14504 39865 14532
rect 23661 14467 23719 14473
rect 23661 14433 23673 14467
rect 23707 14464 23719 14467
rect 24949 14467 25007 14473
rect 24949 14464 24961 14467
rect 23707 14436 24961 14464
rect 23707 14433 23719 14436
rect 23661 14427 23719 14433
rect 24949 14433 24961 14436
rect 24995 14464 25007 14467
rect 27614 14464 27620 14476
rect 24995 14436 27620 14464
rect 24995 14433 25007 14436
rect 24949 14427 25007 14433
rect 27614 14424 27620 14436
rect 27672 14464 27678 14476
rect 28905 14467 28963 14473
rect 28905 14464 28917 14467
rect 27672 14436 28917 14464
rect 27672 14424 27678 14436
rect 28905 14433 28917 14436
rect 28951 14464 28963 14467
rect 29549 14467 29607 14473
rect 29549 14464 29561 14467
rect 28951 14436 29561 14464
rect 28951 14433 28963 14436
rect 28905 14427 28963 14433
rect 29549 14433 29561 14436
rect 29595 14433 29607 14467
rect 29549 14427 29607 14433
rect 29822 14424 29828 14476
rect 29880 14424 29886 14476
rect 29914 14424 29920 14476
rect 29972 14464 29978 14476
rect 29972 14436 31524 14464
rect 29972 14424 29978 14436
rect 21361 14399 21419 14405
rect 21361 14365 21373 14399
rect 21407 14396 21419 14399
rect 21637 14399 21695 14405
rect 21407 14368 21588 14396
rect 21407 14365 21419 14368
rect 21361 14359 21419 14365
rect 2774 14288 2780 14340
rect 2832 14328 2838 14340
rect 3970 14328 3976 14340
rect 2832 14300 3976 14328
rect 2832 14288 2838 14300
rect 3970 14288 3976 14300
rect 4028 14288 4034 14340
rect 4614 14288 4620 14340
rect 4672 14328 4678 14340
rect 4672 14300 5566 14328
rect 4672 14288 4678 14300
rect 9858 14288 9864 14340
rect 9916 14328 9922 14340
rect 10505 14331 10563 14337
rect 10505 14328 10517 14331
rect 9916 14300 10517 14328
rect 9916 14288 9922 14300
rect 10505 14297 10517 14300
rect 10551 14297 10563 14331
rect 10505 14291 10563 14297
rect 16206 14288 16212 14340
rect 16264 14288 16270 14340
rect 18506 14328 18512 14340
rect 17434 14300 18512 14328
rect 18506 14288 18512 14300
rect 18564 14288 18570 14340
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19521 14331 19579 14337
rect 19521 14328 19533 14331
rect 19208 14300 19533 14328
rect 19208 14288 19214 14300
rect 19521 14297 19533 14300
rect 19567 14297 19579 14331
rect 19521 14291 19579 14297
rect 19613 14331 19671 14337
rect 19613 14297 19625 14331
rect 19659 14328 19671 14331
rect 20254 14328 20260 14340
rect 19659 14300 20260 14328
rect 19659 14297 19671 14300
rect 19613 14291 19671 14297
rect 20254 14288 20260 14300
rect 20312 14288 20318 14340
rect 21450 14288 21456 14340
rect 21508 14288 21514 14340
rect 21560 14328 21588 14368
rect 21637 14365 21649 14399
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 26786 14356 26792 14408
rect 26844 14356 26850 14408
rect 31496 14405 31524 14436
rect 31938 14424 31944 14476
rect 31996 14424 32002 14476
rect 32214 14424 32220 14476
rect 32272 14424 32278 14476
rect 34241 14467 34299 14473
rect 34241 14433 34253 14467
rect 34287 14464 34299 14467
rect 38102 14464 38108 14476
rect 34287 14436 38108 14464
rect 34287 14433 34299 14436
rect 34241 14427 34299 14433
rect 38102 14424 38108 14436
rect 38160 14424 38166 14476
rect 38933 14467 38991 14473
rect 38933 14464 38945 14467
rect 38304 14436 38945 14464
rect 26973 14399 27031 14405
rect 26973 14365 26985 14399
rect 27019 14396 27031 14399
rect 31481 14399 31539 14405
rect 27019 14368 27200 14396
rect 27019 14365 27031 14368
rect 26973 14359 27031 14365
rect 22094 14328 22100 14340
rect 21560 14300 22100 14328
rect 22094 14288 22100 14300
rect 22152 14288 22158 14340
rect 22830 14288 22836 14340
rect 22888 14288 22894 14340
rect 23385 14331 23443 14337
rect 23385 14297 23397 14331
rect 23431 14328 23443 14331
rect 23750 14328 23756 14340
rect 23431 14300 23756 14328
rect 23431 14297 23443 14300
rect 23385 14291 23443 14297
rect 23750 14288 23756 14300
rect 23808 14288 23814 14340
rect 25225 14331 25283 14337
rect 25225 14297 25237 14331
rect 25271 14328 25283 14331
rect 25314 14328 25320 14340
rect 25271 14300 25320 14328
rect 25271 14297 25283 14300
rect 25225 14291 25283 14297
rect 25314 14288 25320 14300
rect 25372 14288 25378 14340
rect 25424 14300 25714 14328
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 6549 14263 6607 14269
rect 6549 14260 6561 14263
rect 6052 14232 6561 14260
rect 6052 14220 6058 14232
rect 6549 14229 6561 14232
rect 6595 14229 6607 14263
rect 6549 14223 6607 14229
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 12802 14260 12808 14272
rect 11756 14232 12808 14260
rect 11756 14220 11762 14232
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 18012 14232 19257 14260
rect 18012 14220 18018 14232
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 19978 14220 19984 14272
rect 20036 14220 20042 14272
rect 21082 14220 21088 14272
rect 21140 14220 21146 14272
rect 24762 14220 24768 14272
rect 24820 14260 24826 14272
rect 25424 14260 25452 14300
rect 26510 14288 26516 14340
rect 26568 14328 26574 14340
rect 26878 14328 26884 14340
rect 26568 14300 26884 14328
rect 26568 14288 26574 14300
rect 26878 14288 26884 14300
rect 26936 14288 26942 14340
rect 24820 14232 25452 14260
rect 24820 14220 24826 14232
rect 26694 14220 26700 14272
rect 26752 14220 26758 14272
rect 27172 14269 27200 14368
rect 31481 14365 31493 14399
rect 31527 14365 31539 14399
rect 31481 14359 31539 14365
rect 34149 14399 34207 14405
rect 34149 14365 34161 14399
rect 34195 14396 34207 14399
rect 34330 14396 34336 14408
rect 34195 14368 34336 14396
rect 34195 14365 34207 14368
rect 34149 14359 34207 14365
rect 34330 14356 34336 14368
rect 34388 14356 34394 14408
rect 35158 14356 35164 14408
rect 35216 14356 35222 14408
rect 38197 14399 38255 14405
rect 38197 14365 38209 14399
rect 38243 14398 38255 14399
rect 38304 14398 38332 14436
rect 38933 14433 38945 14436
rect 38979 14433 38991 14467
rect 38933 14427 38991 14433
rect 38243 14370 38332 14398
rect 38243 14365 38255 14370
rect 38197 14359 38255 14365
rect 38378 14356 38384 14408
rect 38436 14356 38442 14408
rect 38470 14356 38476 14408
rect 38528 14405 38534 14408
rect 38528 14399 38557 14405
rect 38545 14365 38557 14399
rect 38528 14359 38557 14365
rect 38528 14356 38534 14359
rect 38654 14356 38660 14408
rect 38712 14356 38718 14408
rect 28629 14331 28687 14337
rect 28198 14300 28580 14328
rect 27157 14263 27215 14269
rect 27157 14229 27169 14263
rect 27203 14260 27215 14263
rect 28350 14260 28356 14272
rect 27203 14232 28356 14260
rect 27203 14229 27215 14232
rect 27157 14223 27215 14229
rect 28350 14220 28356 14232
rect 28408 14220 28414 14272
rect 28552 14260 28580 14300
rect 28629 14297 28641 14331
rect 28675 14328 28687 14331
rect 29086 14328 29092 14340
rect 28675 14300 29092 14328
rect 28675 14297 28687 14300
rect 28629 14291 28687 14297
rect 29086 14288 29092 14300
rect 29144 14288 29150 14340
rect 30374 14288 30380 14340
rect 30432 14288 30438 14340
rect 31846 14288 31852 14340
rect 31904 14288 31910 14340
rect 32950 14288 32956 14340
rect 33008 14288 33014 14340
rect 34422 14288 34428 14340
rect 34480 14328 34486 14340
rect 35805 14331 35863 14337
rect 35805 14328 35817 14331
rect 34480 14300 35817 14328
rect 34480 14288 34486 14300
rect 35805 14297 35817 14300
rect 35851 14297 35863 14331
rect 35805 14291 35863 14297
rect 38289 14331 38347 14337
rect 38289 14297 38301 14331
rect 38335 14328 38347 14331
rect 39040 14328 39068 14504
rect 39853 14501 39865 14504
rect 39899 14501 39911 14535
rect 39853 14495 39911 14501
rect 39574 14464 39580 14476
rect 39408 14436 39580 14464
rect 39114 14356 39120 14408
rect 39172 14356 39178 14408
rect 39206 14356 39212 14408
rect 39264 14396 39270 14408
rect 39408 14405 39436 14436
rect 39574 14424 39580 14436
rect 39632 14464 39638 14476
rect 39632 14436 39988 14464
rect 39632 14424 39638 14436
rect 39301 14399 39359 14405
rect 39301 14396 39313 14399
rect 39264 14368 39313 14396
rect 39264 14356 39270 14368
rect 39301 14365 39313 14368
rect 39347 14365 39359 14399
rect 39301 14359 39359 14365
rect 39393 14399 39451 14405
rect 39393 14365 39405 14399
rect 39439 14365 39451 14399
rect 39393 14359 39451 14365
rect 39482 14356 39488 14408
rect 39540 14356 39546 14408
rect 39669 14399 39727 14405
rect 39669 14365 39681 14399
rect 39715 14396 39727 14399
rect 39758 14396 39764 14408
rect 39715 14368 39764 14396
rect 39715 14365 39727 14368
rect 39669 14359 39727 14365
rect 39758 14356 39764 14368
rect 39816 14356 39822 14408
rect 39850 14356 39856 14408
rect 39908 14356 39914 14408
rect 39960 14405 39988 14436
rect 40034 14424 40040 14476
rect 40092 14464 40098 14476
rect 40221 14467 40279 14473
rect 40221 14464 40233 14467
rect 40092 14436 40233 14464
rect 40092 14424 40098 14436
rect 40221 14433 40233 14436
rect 40267 14433 40279 14467
rect 40221 14427 40279 14433
rect 39945 14399 40003 14405
rect 39945 14365 39957 14399
rect 39991 14365 40003 14399
rect 39945 14359 40003 14365
rect 41506 14356 41512 14408
rect 41564 14356 41570 14408
rect 38335 14300 39068 14328
rect 40129 14331 40187 14337
rect 38335 14297 38347 14300
rect 38289 14291 38347 14297
rect 40129 14297 40141 14331
rect 40175 14297 40187 14331
rect 40129 14291 40187 14297
rect 28810 14260 28816 14272
rect 28552 14232 28816 14260
rect 28810 14220 28816 14232
rect 28868 14260 28874 14272
rect 29270 14260 29276 14272
rect 28868 14232 29276 14260
rect 28868 14220 28874 14232
rect 29270 14220 29276 14232
rect 29328 14220 29334 14272
rect 30558 14220 30564 14272
rect 30616 14260 30622 14272
rect 31297 14263 31355 14269
rect 31297 14260 31309 14263
rect 30616 14232 31309 14260
rect 30616 14220 30622 14232
rect 31297 14229 31309 14232
rect 31343 14229 31355 14263
rect 31297 14223 31355 14229
rect 33689 14263 33747 14269
rect 33689 14229 33701 14263
rect 33735 14260 33747 14263
rect 33870 14260 33876 14272
rect 33735 14232 33876 14260
rect 33735 14229 33747 14232
rect 33689 14223 33747 14229
rect 33870 14220 33876 14232
rect 33928 14260 33934 14272
rect 34606 14260 34612 14272
rect 33928 14232 34612 14260
rect 33928 14220 33934 14232
rect 34606 14220 34612 14232
rect 34664 14220 34670 14272
rect 35342 14220 35348 14272
rect 35400 14260 35406 14272
rect 37918 14260 37924 14272
rect 35400 14232 37924 14260
rect 35400 14220 35406 14232
rect 37918 14220 37924 14232
rect 37976 14260 37982 14272
rect 38378 14260 38384 14272
rect 37976 14232 38384 14260
rect 37976 14220 37982 14232
rect 38378 14220 38384 14232
rect 38436 14220 38442 14272
rect 39114 14220 39120 14272
rect 39172 14260 39178 14272
rect 40144 14260 40172 14291
rect 39172 14232 40172 14260
rect 39172 14220 39178 14232
rect 1104 14170 42504 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 42504 14170
rect 1104 14096 42504 14118
rect 2222 14016 2228 14068
rect 2280 14056 2286 14068
rect 2317 14059 2375 14065
rect 2317 14056 2329 14059
rect 2280 14028 2329 14056
rect 2280 14016 2286 14028
rect 2317 14025 2329 14028
rect 2363 14025 2375 14059
rect 4798 14056 4804 14068
rect 2317 14019 2375 14025
rect 2746 14028 4804 14056
rect 2746 13988 2774 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 5813 14059 5871 14065
rect 5813 14056 5825 14059
rect 5684 14028 5825 14056
rect 5684 14016 5690 14028
rect 5813 14025 5825 14028
rect 5859 14056 5871 14059
rect 6733 14059 6791 14065
rect 6733 14056 6745 14059
rect 5859 14028 6745 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 6733 14025 6745 14028
rect 6779 14025 6791 14059
rect 11698 14056 11704 14068
rect 6733 14019 6791 14025
rect 11164 14028 11704 14056
rect 4614 13988 4620 14000
rect 1688 13960 2774 13988
rect 4554 13960 4620 13988
rect 1688 13929 1716 13960
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 4706 13948 4712 14000
rect 4764 13988 4770 14000
rect 5261 13991 5319 13997
rect 5261 13988 5273 13991
rect 4764 13960 5273 13988
rect 4764 13948 4770 13960
rect 5261 13957 5273 13960
rect 5307 13957 5319 13991
rect 5261 13951 5319 13957
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 5276 13920 5304 13951
rect 5350 13948 5356 14000
rect 5408 13988 5414 14000
rect 5461 13991 5519 13997
rect 5461 13988 5473 13991
rect 5408 13960 5473 13988
rect 5408 13948 5414 13960
rect 5461 13957 5473 13960
rect 5507 13957 5519 13991
rect 5461 13951 5519 13957
rect 5994 13948 6000 14000
rect 6052 13948 6058 14000
rect 6086 13948 6092 14000
rect 6144 13988 6150 14000
rect 6546 13988 6552 14000
rect 6144 13960 6552 13988
rect 6144 13948 6150 13960
rect 6546 13948 6552 13960
rect 6604 13988 6610 14000
rect 6641 13991 6699 13997
rect 6641 13988 6653 13991
rect 6604 13960 6653 13988
rect 6604 13948 6610 13960
rect 6641 13957 6653 13960
rect 6687 13957 6699 13991
rect 6641 13951 6699 13957
rect 9858 13948 9864 14000
rect 9916 13948 9922 14000
rect 10318 13948 10324 14000
rect 10376 13948 10382 14000
rect 5626 13920 5632 13932
rect 5276 13892 5632 13920
rect 1673 13883 1731 13889
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 2958 13812 2964 13864
rect 3016 13812 3022 13864
rect 3050 13812 3056 13864
rect 3108 13812 3114 13864
rect 3326 13812 3332 13864
rect 3384 13812 3390 13864
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5442 13852 5448 13864
rect 5123 13824 5448 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 1486 13676 1492 13728
rect 1544 13676 1550 13728
rect 5442 13676 5448 13728
rect 5500 13676 5506 13728
rect 5629 13719 5687 13725
rect 5629 13685 5641 13719
rect 5675 13716 5687 13719
rect 5736 13716 5764 13883
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 9398 13920 9404 13932
rect 8352 13892 9404 13920
rect 8352 13880 8358 13892
rect 9398 13880 9404 13892
rect 9456 13920 9462 13932
rect 9585 13923 9643 13929
rect 9585 13920 9597 13923
rect 9456 13892 9597 13920
rect 9456 13880 9462 13892
rect 9585 13889 9597 13892
rect 9631 13889 9643 13923
rect 11164 13920 11192 14028
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 11974 14016 11980 14068
rect 12032 14016 12038 14068
rect 12158 14016 12164 14068
rect 12216 14016 12222 14068
rect 12342 14016 12348 14068
rect 12400 14056 12406 14068
rect 12400 14028 18092 14056
rect 12400 14016 12406 14028
rect 12250 13948 12256 14000
rect 12308 13988 12314 14000
rect 12713 13991 12771 13997
rect 12713 13988 12725 13991
rect 12308 13960 12725 13988
rect 12308 13948 12314 13960
rect 12713 13957 12725 13960
rect 12759 13957 12771 13991
rect 12713 13951 12771 13957
rect 18064 13932 18092 14028
rect 18414 14016 18420 14068
rect 18472 14016 18478 14068
rect 19794 14056 19800 14068
rect 19168 14028 19800 14056
rect 18506 13948 18512 14000
rect 18564 13988 18570 14000
rect 19168 13988 19196 14028
rect 19794 14016 19800 14028
rect 19852 14016 19858 14068
rect 20257 14059 20315 14065
rect 20257 14025 20269 14059
rect 20303 14056 20315 14059
rect 20530 14056 20536 14068
rect 20303 14028 20536 14056
rect 20303 14025 20315 14028
rect 20257 14019 20315 14025
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 22097 14059 22155 14065
rect 22097 14025 22109 14059
rect 22143 14056 22155 14059
rect 22278 14056 22284 14068
rect 22143 14028 22284 14056
rect 22143 14025 22155 14028
rect 22097 14019 22155 14025
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 23750 14016 23756 14068
rect 23808 14016 23814 14068
rect 25130 14056 25136 14068
rect 23860 14028 25136 14056
rect 18564 13960 19274 13988
rect 18564 13948 18570 13960
rect 9585 13883 9643 13889
rect 11072 13892 11192 13920
rect 11517 13923 11575 13929
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 11072 13852 11100 13892
rect 11517 13889 11529 13923
rect 11563 13920 11575 13923
rect 11790 13920 11796 13932
rect 11563 13892 11796 13920
rect 11563 13889 11575 13892
rect 11517 13883 11575 13889
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 11974 13920 11980 13932
rect 11931 13892 11980 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 11974 13880 11980 13892
rect 12032 13880 12038 13932
rect 12069 13923 12127 13929
rect 12069 13889 12081 13923
rect 12115 13920 12127 13923
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 12115 13892 12173 13920
rect 12115 13889 12127 13892
rect 12069 13883 12127 13889
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13920 12403 13923
rect 12802 13920 12808 13932
rect 12391 13892 12808 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 12084 13852 12112 13883
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 5960 13824 6040 13852
rect 5960 13812 5966 13824
rect 6012 13793 6040 13824
rect 9692 13824 11100 13852
rect 11348 13824 12112 13852
rect 5997 13787 6055 13793
rect 5997 13753 6009 13787
rect 6043 13753 6055 13787
rect 5997 13747 6055 13753
rect 8754 13744 8760 13796
rect 8812 13784 8818 13796
rect 9692 13784 9720 13824
rect 8812 13756 9720 13784
rect 8812 13744 8818 13756
rect 11348 13728 11376 13824
rect 11974 13744 11980 13796
rect 12032 13784 12038 13796
rect 12912 13784 12940 13883
rect 18046 13880 18052 13932
rect 18104 13880 18110 13932
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13920 21051 13923
rect 22094 13920 22100 13932
rect 21039 13892 22100 13920
rect 21039 13889 21051 13892
rect 20993 13883 21051 13889
rect 22094 13880 22100 13892
rect 22152 13920 22158 13932
rect 22922 13920 22928 13932
rect 22152 13892 22928 13920
rect 22152 13880 22158 13892
rect 22922 13880 22928 13892
rect 22980 13880 22986 13932
rect 23106 13880 23112 13932
rect 23164 13880 23170 13932
rect 23860 13929 23888 14028
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 25590 14016 25596 14068
rect 25648 14016 25654 14068
rect 25685 14059 25743 14065
rect 25685 14025 25697 14059
rect 25731 14025 25743 14059
rect 25685 14019 25743 14025
rect 24118 13948 24124 14000
rect 24176 13948 24182 14000
rect 24762 13948 24768 14000
rect 24820 13948 24826 14000
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13889 23903 13923
rect 23845 13883 23903 13889
rect 25590 13880 25596 13932
rect 25648 13920 25654 13932
rect 25700 13920 25728 14019
rect 25774 14016 25780 14068
rect 25832 14056 25838 14068
rect 26053 14059 26111 14065
rect 26053 14056 26065 14059
rect 25832 14028 26065 14056
rect 25832 14016 25838 14028
rect 26053 14025 26065 14028
rect 26099 14056 26111 14059
rect 26878 14056 26884 14068
rect 26099 14028 26884 14056
rect 26099 14025 26111 14028
rect 26053 14019 26111 14025
rect 26878 14016 26884 14028
rect 26936 14016 26942 14068
rect 27430 14016 27436 14068
rect 27488 14056 27494 14068
rect 32398 14056 32404 14068
rect 27488 14028 32404 14056
rect 27488 14016 27494 14028
rect 32398 14016 32404 14028
rect 32456 14016 32462 14068
rect 32493 14059 32551 14065
rect 32493 14025 32505 14059
rect 32539 14056 32551 14059
rect 33042 14056 33048 14068
rect 32539 14028 33048 14056
rect 32539 14025 32551 14028
rect 32493 14019 32551 14025
rect 33042 14016 33048 14028
rect 33100 14056 33106 14068
rect 33100 14028 34744 14056
rect 33100 14016 33106 14028
rect 29086 13948 29092 14000
rect 29144 13948 29150 14000
rect 29270 13948 29276 14000
rect 29328 13988 29334 14000
rect 29328 13960 30958 13988
rect 29328 13948 29334 13960
rect 32950 13948 32956 14000
rect 33008 13948 33014 14000
rect 25648 13892 25728 13920
rect 25648 13880 25654 13892
rect 26694 13880 26700 13932
rect 26752 13920 26758 13932
rect 27525 13923 27583 13929
rect 27525 13920 27537 13923
rect 26752 13892 27537 13920
rect 26752 13880 26758 13892
rect 27525 13889 27537 13892
rect 27571 13889 27583 13923
rect 27525 13883 27583 13889
rect 27890 13880 27896 13932
rect 27948 13920 27954 13932
rect 34716 13929 34744 14028
rect 34790 14016 34796 14068
rect 34848 14056 34854 14068
rect 34977 14059 35035 14065
rect 34977 14056 34989 14059
rect 34848 14028 34989 14056
rect 34848 14016 34854 14028
rect 34977 14025 34989 14028
rect 35023 14056 35035 14059
rect 35158 14056 35164 14068
rect 35023 14028 35164 14056
rect 35023 14025 35035 14028
rect 34977 14019 35035 14025
rect 35158 14016 35164 14028
rect 35216 14016 35222 14068
rect 37274 14016 37280 14068
rect 37332 14056 37338 14068
rect 38289 14059 38347 14065
rect 38289 14056 38301 14059
rect 37332 14028 38301 14056
rect 37332 14016 37338 14028
rect 38289 14025 38301 14028
rect 38335 14056 38347 14059
rect 38378 14056 38384 14068
rect 38335 14028 38384 14056
rect 38335 14025 38347 14028
rect 38289 14019 38347 14025
rect 38378 14016 38384 14028
rect 38436 14056 38442 14068
rect 38562 14056 38568 14068
rect 38436 14028 38568 14056
rect 38436 14016 38442 14028
rect 38562 14016 38568 14028
rect 38620 14016 38626 14068
rect 38933 14059 38991 14065
rect 38933 14025 38945 14059
rect 38979 14056 38991 14059
rect 39942 14056 39948 14068
rect 38979 14028 39948 14056
rect 38979 14025 38991 14028
rect 38933 14019 38991 14025
rect 39942 14016 39948 14028
rect 40000 14016 40006 14068
rect 41049 14059 41107 14065
rect 41049 14025 41061 14059
rect 41095 14056 41107 14059
rect 41138 14056 41144 14068
rect 41095 14028 41144 14056
rect 41095 14025 41107 14028
rect 41049 14019 41107 14025
rect 41138 14016 41144 14028
rect 41196 14016 41202 14068
rect 36446 13948 36452 14000
rect 36504 13948 36510 14000
rect 39758 13948 39764 14000
rect 39816 13988 39822 14000
rect 40037 13991 40095 13997
rect 40037 13988 40049 13991
rect 39816 13960 40049 13988
rect 39816 13948 39822 13960
rect 40037 13957 40049 13960
rect 40083 13988 40095 13991
rect 41414 13988 41420 14000
rect 40083 13960 41420 13988
rect 40083 13957 40095 13960
rect 40037 13951 40095 13957
rect 41414 13948 41420 13960
rect 41472 13948 41478 14000
rect 30193 13923 30251 13929
rect 30193 13920 30205 13923
rect 27948 13892 30205 13920
rect 27948 13880 27954 13892
rect 30193 13889 30205 13892
rect 30239 13889 30251 13923
rect 30193 13883 30251 13889
rect 34701 13923 34759 13929
rect 34701 13889 34713 13923
rect 34747 13889 34759 13923
rect 34701 13883 34759 13889
rect 35342 13880 35348 13932
rect 35400 13880 35406 13932
rect 38197 13923 38255 13929
rect 38197 13889 38209 13923
rect 38243 13920 38255 13923
rect 38286 13920 38292 13932
rect 38243 13892 38292 13920
rect 38243 13889 38255 13892
rect 38197 13883 38255 13889
rect 38286 13880 38292 13892
rect 38344 13880 38350 13932
rect 38657 13923 38715 13929
rect 38657 13889 38669 13923
rect 38703 13920 38715 13923
rect 39114 13920 39120 13932
rect 38703 13892 39120 13920
rect 38703 13889 38715 13892
rect 38657 13883 38715 13889
rect 39114 13880 39120 13892
rect 39172 13880 39178 13932
rect 39298 13880 39304 13932
rect 39356 13880 39362 13932
rect 39482 13880 39488 13932
rect 39540 13920 39546 13932
rect 39853 13923 39911 13929
rect 39853 13920 39865 13923
rect 39540 13892 39865 13920
rect 39540 13880 39546 13892
rect 39853 13889 39865 13892
rect 39899 13889 39911 13923
rect 39853 13883 39911 13889
rect 40957 13923 41015 13929
rect 40957 13889 40969 13923
rect 41003 13920 41015 13923
rect 41509 13923 41567 13929
rect 41509 13920 41521 13923
rect 41003 13892 41521 13920
rect 41003 13889 41015 13892
rect 40957 13883 41015 13889
rect 41509 13889 41521 13892
rect 41555 13889 41567 13923
rect 41509 13883 41567 13889
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16500 13824 16681 13852
rect 16500 13796 16528 13824
rect 16669 13821 16681 13824
rect 16715 13852 16727 13855
rect 17034 13852 17040 13864
rect 16715 13824 17040 13852
rect 16715 13821 16727 13824
rect 16669 13815 16727 13821
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 18506 13812 18512 13864
rect 18564 13812 18570 13864
rect 18782 13812 18788 13864
rect 18840 13812 18846 13864
rect 21634 13812 21640 13864
rect 21692 13812 21698 13864
rect 22370 13812 22376 13864
rect 22428 13852 22434 13864
rect 22649 13855 22707 13861
rect 22649 13852 22661 13855
rect 22428 13824 22661 13852
rect 22428 13812 22434 13824
rect 22649 13821 22661 13824
rect 22695 13821 22707 13855
rect 22649 13815 22707 13821
rect 22830 13812 22836 13864
rect 22888 13852 22894 13864
rect 25682 13852 25688 13864
rect 22888 13824 25688 13852
rect 22888 13812 22894 13824
rect 25682 13812 25688 13824
rect 25740 13852 25746 13864
rect 25740 13824 25820 13852
rect 25740 13812 25746 13824
rect 12032 13756 12940 13784
rect 12032 13744 12038 13756
rect 16482 13744 16488 13796
rect 16540 13744 16546 13796
rect 25792 13784 25820 13824
rect 25866 13812 25872 13864
rect 25924 13852 25930 13864
rect 26145 13855 26203 13861
rect 26145 13852 26157 13855
rect 25924 13824 26157 13852
rect 25924 13812 25930 13824
rect 26145 13821 26157 13824
rect 26191 13821 26203 13855
rect 26145 13815 26203 13821
rect 26329 13855 26387 13861
rect 26329 13821 26341 13855
rect 26375 13821 26387 13855
rect 26329 13815 26387 13821
rect 26050 13784 26056 13796
rect 25792 13756 26056 13784
rect 26050 13744 26056 13756
rect 26108 13744 26114 13796
rect 26344 13784 26372 13815
rect 28350 13812 28356 13864
rect 28408 13812 28414 13864
rect 28442 13812 28448 13864
rect 28500 13812 28506 13864
rect 30466 13812 30472 13864
rect 30524 13812 30530 13864
rect 31941 13855 31999 13861
rect 31941 13821 31953 13855
rect 31987 13852 31999 13855
rect 32122 13852 32128 13864
rect 31987 13824 32128 13852
rect 31987 13821 31999 13824
rect 31941 13815 31999 13821
rect 32122 13812 32128 13824
rect 32180 13812 32186 13864
rect 33962 13812 33968 13864
rect 34020 13812 34026 13864
rect 34241 13855 34299 13861
rect 34241 13821 34253 13855
rect 34287 13852 34299 13855
rect 34287 13824 34560 13852
rect 34287 13821 34299 13824
rect 34241 13815 34299 13821
rect 28258 13784 28264 13796
rect 26344 13756 28264 13784
rect 5810 13716 5816 13728
rect 5675 13688 5816 13716
rect 5675 13685 5687 13688
rect 5629 13679 5687 13685
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 11330 13676 11336 13728
rect 11388 13676 11394 13728
rect 12526 13676 12532 13728
rect 12584 13676 12590 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 16390 13716 16396 13728
rect 15344 13688 16396 13716
rect 15344 13676 15350 13688
rect 16390 13676 16396 13688
rect 16448 13676 16454 13728
rect 16932 13719 16990 13725
rect 16932 13685 16944 13719
rect 16978 13716 16990 13719
rect 17954 13716 17960 13728
rect 16978 13688 17960 13716
rect 16978 13685 16990 13688
rect 16932 13679 16990 13685
rect 17954 13676 17960 13688
rect 18012 13676 18018 13728
rect 23474 13676 23480 13728
rect 23532 13716 23538 13728
rect 26344 13716 26372 13756
rect 28258 13744 28264 13756
rect 28316 13744 28322 13796
rect 32306 13744 32312 13796
rect 32364 13784 32370 13796
rect 32950 13784 32956 13796
rect 32364 13756 32956 13784
rect 32364 13744 32370 13756
rect 32950 13744 32956 13756
rect 33008 13744 33014 13796
rect 34330 13744 34336 13796
rect 34388 13744 34394 13796
rect 34532 13784 34560 13824
rect 34606 13812 34612 13864
rect 34664 13812 34670 13864
rect 36725 13855 36783 13861
rect 36725 13852 36737 13855
rect 35452 13824 36737 13852
rect 35452 13796 35480 13824
rect 36725 13821 36737 13824
rect 36771 13852 36783 13855
rect 38933 13855 38991 13861
rect 36771 13824 37228 13852
rect 36771 13821 36783 13824
rect 36725 13815 36783 13821
rect 35434 13784 35440 13796
rect 34532 13756 35440 13784
rect 35434 13744 35440 13756
rect 35492 13744 35498 13796
rect 37200 13784 37228 13824
rect 38933 13821 38945 13855
rect 38979 13852 38991 13855
rect 39206 13852 39212 13864
rect 38979 13824 39212 13852
rect 38979 13821 38991 13824
rect 38933 13815 38991 13821
rect 39206 13812 39212 13824
rect 39264 13852 39270 13864
rect 39316 13852 39344 13880
rect 39264 13824 39344 13852
rect 39264 13812 39270 13824
rect 39758 13812 39764 13864
rect 39816 13852 39822 13864
rect 40221 13855 40279 13861
rect 40221 13852 40233 13855
rect 39816 13824 40233 13852
rect 39816 13812 39822 13824
rect 40221 13821 40233 13824
rect 40267 13821 40279 13855
rect 40221 13815 40279 13821
rect 41141 13855 41199 13861
rect 41141 13821 41153 13855
rect 41187 13821 41199 13855
rect 41141 13815 41199 13821
rect 37458 13784 37464 13796
rect 37200 13756 37464 13784
rect 37458 13744 37464 13756
rect 37516 13744 37522 13796
rect 37642 13744 37648 13796
rect 37700 13784 37706 13796
rect 38194 13784 38200 13796
rect 37700 13756 38200 13784
rect 37700 13744 37706 13756
rect 38194 13744 38200 13756
rect 38252 13784 38258 13796
rect 40770 13784 40776 13796
rect 38252 13756 40776 13784
rect 38252 13744 38258 13756
rect 40770 13744 40776 13756
rect 40828 13784 40834 13796
rect 41156 13784 41184 13815
rect 42150 13812 42156 13864
rect 42208 13812 42214 13864
rect 40828 13756 41184 13784
rect 40828 13744 40834 13756
rect 23532 13688 26372 13716
rect 23532 13676 23538 13688
rect 26970 13676 26976 13728
rect 27028 13676 27034 13728
rect 27706 13676 27712 13728
rect 27764 13676 27770 13728
rect 38749 13719 38807 13725
rect 38749 13685 38761 13719
rect 38795 13716 38807 13719
rect 39390 13716 39396 13728
rect 38795 13688 39396 13716
rect 38795 13685 38807 13688
rect 38749 13679 38807 13685
rect 39390 13676 39396 13688
rect 39448 13676 39454 13728
rect 40589 13719 40647 13725
rect 40589 13685 40601 13719
rect 40635 13716 40647 13719
rect 40678 13716 40684 13728
rect 40635 13688 40684 13716
rect 40635 13685 40647 13688
rect 40589 13679 40647 13685
rect 40678 13676 40684 13688
rect 40736 13676 40742 13728
rect 1104 13626 42504 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 42504 13626
rect 1104 13552 42504 13574
rect 2958 13472 2964 13524
rect 3016 13512 3022 13524
rect 3191 13515 3249 13521
rect 3191 13512 3203 13515
rect 3016 13484 3203 13512
rect 3016 13472 3022 13484
rect 3191 13481 3203 13484
rect 3237 13481 3249 13515
rect 3191 13475 3249 13481
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 5261 13515 5319 13521
rect 5261 13512 5273 13515
rect 3384 13484 5273 13512
rect 3384 13472 3390 13484
rect 5261 13481 5273 13484
rect 5307 13481 5319 13515
rect 5261 13475 5319 13481
rect 6546 13472 6552 13524
rect 6604 13472 6610 13524
rect 8481 13515 8539 13521
rect 8481 13512 8493 13515
rect 6656 13484 8493 13512
rect 4985 13447 5043 13453
rect 4985 13413 4997 13447
rect 5031 13413 5043 13447
rect 4985 13407 5043 13413
rect 1578 13336 1584 13388
rect 1636 13376 1642 13388
rect 1765 13379 1823 13385
rect 1765 13376 1777 13379
rect 1636 13348 1777 13376
rect 1636 13336 1642 13348
rect 1765 13345 1777 13348
rect 1811 13345 1823 13379
rect 1765 13339 1823 13345
rect 1394 13268 1400 13320
rect 1452 13268 1458 13320
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 5000 13308 5028 13407
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 6656 13444 6684 13484
rect 8481 13481 8493 13484
rect 8527 13512 8539 13515
rect 8527 13484 9260 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 5408 13416 6684 13444
rect 9232 13444 9260 13484
rect 10686 13472 10692 13524
rect 10744 13512 10750 13524
rect 10965 13515 11023 13521
rect 10965 13512 10977 13515
rect 10744 13484 10977 13512
rect 10744 13472 10750 13484
rect 10965 13481 10977 13484
rect 11011 13481 11023 13515
rect 10965 13475 11023 13481
rect 15286 13472 15292 13524
rect 15344 13472 15350 13524
rect 21910 13512 21916 13524
rect 15764 13484 21916 13512
rect 11606 13444 11612 13456
rect 9232 13416 11612 13444
rect 5408 13404 5414 13416
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 5718 13376 5724 13388
rect 5592 13348 5724 13376
rect 5592 13336 5598 13348
rect 5718 13336 5724 13348
rect 5776 13376 5782 13388
rect 5776 13348 6040 13376
rect 5776 13336 5782 13348
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4755 13280 4936 13308
rect 5000 13280 5089 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 2774 13200 2780 13252
rect 2832 13200 2838 13252
rect 4706 13132 4712 13184
rect 4764 13172 4770 13184
rect 4801 13175 4859 13181
rect 4801 13172 4813 13175
rect 4764 13144 4813 13172
rect 4764 13132 4770 13144
rect 4801 13141 4813 13144
rect 4847 13141 4859 13175
rect 4908 13172 4936 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5810 13308 5816 13320
rect 5307 13280 5816 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6012 13317 6040 13348
rect 8294 13336 8300 13388
rect 8352 13336 8358 13388
rect 15764 13376 15792 13484
rect 21910 13472 21916 13484
rect 21968 13512 21974 13524
rect 21968 13484 31156 13512
rect 21968 13472 21974 13484
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 19245 13447 19303 13453
rect 19245 13444 19257 13447
rect 18840 13416 19257 13444
rect 18840 13404 18846 13416
rect 19245 13413 19257 13416
rect 19291 13413 19303 13447
rect 19245 13407 19303 13413
rect 21634 13404 21640 13456
rect 21692 13444 21698 13456
rect 22005 13447 22063 13453
rect 22005 13444 22017 13447
rect 21692 13416 22017 13444
rect 21692 13404 21698 13416
rect 22005 13413 22017 13416
rect 22051 13413 22063 13447
rect 22005 13407 22063 13413
rect 23566 13404 23572 13456
rect 23624 13444 23630 13456
rect 23845 13447 23903 13453
rect 23845 13444 23857 13447
rect 23624 13416 23857 13444
rect 23624 13404 23630 13416
rect 23845 13413 23857 13416
rect 23891 13413 23903 13447
rect 23845 13407 23903 13413
rect 25222 13404 25228 13456
rect 25280 13404 25286 13456
rect 26878 13404 26884 13456
rect 26936 13444 26942 13456
rect 27065 13447 27123 13453
rect 27065 13444 27077 13447
rect 26936 13416 27077 13444
rect 26936 13404 26942 13416
rect 27065 13413 27077 13416
rect 27111 13413 27123 13447
rect 27065 13407 27123 13413
rect 28077 13447 28135 13453
rect 28077 13413 28089 13447
rect 28123 13444 28135 13447
rect 28442 13444 28448 13456
rect 28123 13416 28448 13444
rect 28123 13413 28135 13416
rect 28077 13407 28135 13413
rect 28442 13404 28448 13416
rect 28500 13404 28506 13456
rect 28534 13404 28540 13456
rect 28592 13444 28598 13456
rect 28994 13444 29000 13456
rect 28592 13416 29000 13444
rect 28592 13404 28598 13416
rect 28994 13404 29000 13416
rect 29052 13444 29058 13456
rect 29914 13444 29920 13456
rect 29052 13416 29920 13444
rect 29052 13404 29058 13416
rect 29914 13404 29920 13416
rect 29972 13404 29978 13456
rect 10888 13348 15792 13376
rect 5997 13311 6055 13317
rect 5997 13277 6009 13311
rect 6043 13308 6055 13311
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6043 13280 6285 13308
rect 6043 13277 6055 13280
rect 5997 13271 6055 13277
rect 6273 13277 6285 13280
rect 6319 13308 6331 13311
rect 6730 13308 6736 13320
rect 6319 13280 6736 13308
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 6730 13268 6736 13280
rect 6788 13268 6794 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8754 13308 8760 13320
rect 8435 13280 8760 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 10888 13317 10916 13348
rect 16390 13336 16396 13388
rect 16448 13376 16454 13388
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 16448 13348 17601 13376
rect 16448 13336 16454 13348
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 17773 13379 17831 13385
rect 17773 13345 17785 13379
rect 17819 13376 17831 13379
rect 18414 13376 18420 13388
rect 17819 13348 18420 13376
rect 17819 13345 17831 13348
rect 17773 13339 17831 13345
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 20257 13379 20315 13385
rect 20257 13376 20269 13379
rect 18564 13348 20269 13376
rect 18564 13336 18570 13348
rect 20257 13345 20269 13348
rect 20303 13345 20315 13379
rect 20257 13339 20315 13345
rect 20533 13379 20591 13385
rect 20533 13345 20545 13379
rect 20579 13376 20591 13379
rect 21082 13376 21088 13388
rect 20579 13348 21088 13376
rect 20579 13345 20591 13348
rect 20533 13339 20591 13345
rect 21082 13336 21088 13348
rect 21140 13336 21146 13388
rect 22097 13379 22155 13385
rect 22097 13345 22109 13379
rect 22143 13376 22155 13379
rect 22370 13376 22376 13388
rect 22143 13348 22376 13376
rect 22143 13345 22155 13348
rect 22097 13339 22155 13345
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 24854 13336 24860 13388
rect 24912 13376 24918 13388
rect 24912 13348 24992 13376
rect 24912 13336 24918 13348
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 11146 13268 11152 13320
rect 11204 13268 11210 13320
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 11330 13308 11336 13320
rect 11287 13280 11336 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11572 13280 11897 13308
rect 11572 13268 11578 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 14550 13308 14556 13320
rect 13294 13280 14556 13308
rect 11885 13271 11943 13277
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 4985 13243 5043 13249
rect 4985 13209 4997 13243
rect 5031 13240 5043 13243
rect 5442 13240 5448 13252
rect 5031 13212 5448 13240
rect 5031 13209 5043 13212
rect 4985 13203 5043 13209
rect 5442 13200 5448 13212
rect 5500 13200 5506 13252
rect 5828 13240 5856 13268
rect 6089 13243 6147 13249
rect 6089 13240 6101 13243
rect 5828 13212 6101 13240
rect 6089 13209 6101 13212
rect 6135 13209 6147 13243
rect 7590 13212 7972 13240
rect 6089 13203 6147 13209
rect 5350 13172 5356 13184
rect 4908 13144 5356 13172
rect 4801 13135 4859 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 5994 13132 6000 13184
rect 6052 13132 6058 13184
rect 6454 13132 6460 13184
rect 6512 13132 6518 13184
rect 7944 13172 7972 13212
rect 8018 13200 8024 13252
rect 8076 13200 8082 13252
rect 10318 13240 10324 13252
rect 8404 13212 10324 13240
rect 8404 13172 8432 13212
rect 10318 13200 10324 13212
rect 10376 13200 10382 13252
rect 12158 13200 12164 13252
rect 12216 13200 12222 13252
rect 14660 13240 14688 13271
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 18524 13308 18552 13336
rect 17092 13280 18552 13308
rect 19429 13311 19487 13317
rect 17092 13268 17098 13280
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 19702 13308 19708 13320
rect 19475 13280 19708 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13308 19855 13311
rect 19886 13308 19892 13320
rect 19843 13280 19892 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 24210 13268 24216 13320
rect 24268 13308 24274 13320
rect 24670 13308 24676 13320
rect 24268 13280 24676 13308
rect 24268 13268 24274 13280
rect 24670 13268 24676 13280
rect 24728 13268 24734 13320
rect 24964 13317 24992 13348
rect 25590 13336 25596 13388
rect 25648 13336 25654 13388
rect 30558 13376 30564 13388
rect 27908 13348 30564 13376
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13277 25099 13311
rect 25041 13271 25099 13277
rect 13648 13212 14688 13240
rect 7944 13144 8432 13172
rect 9582 13132 9588 13184
rect 9640 13132 9646 13184
rect 11422 13132 11428 13184
rect 11480 13172 11486 13184
rect 11609 13175 11667 13181
rect 11609 13172 11621 13175
rect 11480 13144 11621 13172
rect 11480 13132 11486 13144
rect 11609 13141 11621 13144
rect 11655 13172 11667 13175
rect 12986 13172 12992 13184
rect 11655 13144 12992 13172
rect 11655 13141 11667 13144
rect 11609 13135 11667 13141
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 13446 13132 13452 13184
rect 13504 13172 13510 13184
rect 13648 13181 13676 13212
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 16761 13243 16819 13249
rect 14976 13212 15594 13240
rect 14976 13200 14982 13212
rect 16761 13209 16773 13243
rect 16807 13240 16819 13243
rect 16807 13212 17172 13240
rect 16807 13209 16819 13212
rect 16761 13203 16819 13209
rect 13633 13175 13691 13181
rect 13633 13172 13645 13175
rect 13504 13144 13645 13172
rect 13504 13132 13510 13144
rect 13633 13141 13645 13144
rect 13679 13141 13691 13175
rect 13633 13135 13691 13141
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 17144 13181 17172 13212
rect 19518 13200 19524 13252
rect 19576 13200 19582 13252
rect 19613 13243 19671 13249
rect 19613 13209 19625 13243
rect 19659 13240 19671 13243
rect 19978 13240 19984 13252
rect 19659 13212 19984 13240
rect 19659 13209 19671 13212
rect 19613 13203 19671 13209
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 22373 13243 22431 13249
rect 21758 13212 22094 13240
rect 14093 13175 14151 13181
rect 14093 13172 14105 13175
rect 13780 13144 14105 13172
rect 13780 13132 13786 13144
rect 14093 13141 14105 13144
rect 14139 13141 14151 13175
rect 14093 13135 14151 13141
rect 17129 13175 17187 13181
rect 17129 13141 17141 13175
rect 17175 13141 17187 13175
rect 17129 13135 17187 13141
rect 17497 13175 17555 13181
rect 17497 13141 17509 13175
rect 17543 13172 17555 13175
rect 17862 13172 17868 13184
rect 17543 13144 17868 13172
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 22066 13172 22094 13212
rect 22373 13209 22385 13243
rect 22419 13240 22431 13243
rect 22462 13240 22468 13252
rect 22419 13212 22468 13240
rect 22419 13209 22431 13212
rect 22373 13203 22431 13209
rect 22462 13200 22468 13212
rect 22520 13200 22526 13252
rect 22830 13200 22836 13252
rect 22888 13200 22894 13252
rect 24857 13243 24915 13249
rect 24857 13209 24869 13243
rect 24903 13209 24915 13243
rect 25056 13240 25084 13271
rect 25130 13268 25136 13320
rect 25188 13308 25194 13320
rect 25317 13311 25375 13317
rect 25317 13308 25329 13311
rect 25188 13280 25329 13308
rect 25188 13268 25194 13280
rect 25317 13277 25329 13280
rect 25363 13277 25375 13311
rect 25317 13271 25375 13277
rect 27522 13268 27528 13320
rect 27580 13268 27586 13320
rect 27706 13268 27712 13320
rect 27764 13268 27770 13320
rect 27908 13317 27936 13348
rect 30558 13336 30564 13348
rect 30616 13336 30622 13388
rect 27893 13311 27951 13317
rect 27893 13277 27905 13311
rect 27939 13277 27951 13311
rect 27893 13271 27951 13277
rect 28184 13280 28672 13308
rect 25866 13240 25872 13252
rect 25056 13212 25872 13240
rect 24857 13203 24915 13209
rect 23750 13172 23756 13184
rect 22066 13144 23756 13172
rect 23750 13132 23756 13144
rect 23808 13132 23814 13184
rect 24872 13172 24900 13203
rect 25866 13200 25872 13212
rect 25924 13200 25930 13252
rect 26050 13200 26056 13252
rect 26108 13200 26114 13252
rect 27246 13200 27252 13252
rect 27304 13240 27310 13252
rect 27801 13243 27859 13249
rect 27801 13240 27813 13243
rect 27304 13212 27813 13240
rect 27304 13200 27310 13212
rect 27801 13209 27813 13212
rect 27847 13209 27859 13243
rect 27801 13203 27859 13209
rect 26970 13172 26976 13184
rect 24872 13144 26976 13172
rect 26970 13132 26976 13144
rect 27028 13132 27034 13184
rect 27614 13132 27620 13184
rect 27672 13172 27678 13184
rect 28184 13172 28212 13280
rect 28534 13200 28540 13252
rect 28592 13200 28598 13252
rect 28644 13240 28672 13280
rect 28718 13268 28724 13320
rect 28776 13268 28782 13320
rect 31128 13317 31156 13484
rect 32398 13472 32404 13524
rect 32456 13512 32462 13524
rect 32585 13515 32643 13521
rect 32585 13512 32597 13515
rect 32456 13484 32597 13512
rect 32456 13472 32462 13484
rect 32585 13481 32597 13484
rect 32631 13512 32643 13515
rect 37366 13512 37372 13524
rect 32631 13484 37372 13512
rect 32631 13481 32643 13484
rect 32585 13475 32643 13481
rect 37366 13472 37372 13484
rect 37424 13472 37430 13524
rect 38102 13472 38108 13524
rect 38160 13512 38166 13524
rect 38473 13515 38531 13521
rect 38473 13512 38485 13515
rect 38160 13484 38485 13512
rect 38160 13472 38166 13484
rect 38473 13481 38485 13484
rect 38519 13481 38531 13515
rect 39022 13512 39028 13524
rect 38473 13475 38531 13481
rect 38580 13484 39028 13512
rect 33689 13447 33747 13453
rect 33689 13413 33701 13447
rect 33735 13444 33747 13447
rect 33962 13444 33968 13456
rect 33735 13416 33968 13444
rect 33735 13413 33747 13416
rect 33689 13407 33747 13413
rect 33962 13404 33968 13416
rect 34020 13404 34026 13456
rect 34701 13447 34759 13453
rect 34701 13444 34713 13447
rect 34348 13416 34713 13444
rect 33042 13336 33048 13388
rect 33100 13336 33106 13388
rect 34348 13385 34376 13416
rect 34701 13413 34713 13416
rect 34747 13413 34759 13447
rect 34701 13407 34759 13413
rect 34992 13416 35664 13444
rect 34333 13379 34391 13385
rect 34333 13345 34345 13379
rect 34379 13345 34391 13379
rect 34333 13339 34391 13345
rect 31113 13311 31171 13317
rect 31113 13277 31125 13311
rect 31159 13277 31171 13311
rect 31113 13271 31171 13277
rect 34882 13268 34888 13320
rect 34940 13268 34946 13320
rect 34992 13317 35020 13416
rect 35434 13336 35440 13388
rect 35492 13376 35498 13388
rect 35529 13379 35587 13385
rect 35529 13376 35541 13379
rect 35492 13348 35541 13376
rect 35492 13336 35498 13348
rect 35529 13345 35541 13348
rect 35575 13345 35587 13379
rect 35636 13376 35664 13416
rect 36814 13404 36820 13456
rect 36872 13444 36878 13456
rect 37277 13447 37335 13453
rect 37277 13444 37289 13447
rect 36872 13416 37289 13444
rect 36872 13404 36878 13416
rect 37277 13413 37289 13416
rect 37323 13413 37335 13447
rect 37277 13407 37335 13413
rect 38580 13376 38608 13484
rect 39022 13472 39028 13484
rect 39080 13472 39086 13524
rect 39390 13472 39396 13524
rect 39448 13472 39454 13524
rect 42150 13472 42156 13524
rect 42208 13472 42214 13524
rect 39408 13444 39436 13472
rect 35636 13348 38608 13376
rect 38672 13416 39436 13444
rect 35529 13339 35587 13345
rect 34977 13311 35035 13317
rect 34977 13277 34989 13311
rect 35023 13277 35035 13311
rect 34977 13271 35035 13277
rect 35066 13268 35072 13320
rect 35124 13268 35130 13320
rect 35253 13311 35311 13317
rect 35253 13277 35265 13311
rect 35299 13277 35311 13311
rect 35253 13271 35311 13277
rect 30098 13240 30104 13252
rect 28644 13212 30104 13240
rect 30098 13200 30104 13212
rect 30156 13200 30162 13252
rect 30650 13200 30656 13252
rect 30708 13240 30714 13252
rect 35268 13240 35296 13271
rect 37458 13268 37464 13320
rect 37516 13268 37522 13320
rect 38672 13317 38700 13416
rect 40405 13379 40463 13385
rect 40405 13376 40417 13379
rect 38764 13348 40417 13376
rect 38657 13311 38715 13317
rect 38657 13277 38669 13311
rect 38703 13277 38715 13311
rect 38657 13271 38715 13277
rect 30708 13212 35296 13240
rect 30708 13200 30714 13212
rect 27672 13144 28212 13172
rect 27672 13132 27678 13144
rect 28258 13132 28264 13184
rect 28316 13132 28322 13184
rect 28902 13132 28908 13184
rect 28960 13172 28966 13184
rect 32122 13172 32128 13184
rect 28960 13144 32128 13172
rect 28960 13132 28966 13144
rect 32122 13132 32128 13144
rect 32180 13132 32186 13184
rect 33597 13175 33655 13181
rect 33597 13141 33609 13175
rect 33643 13172 33655 13175
rect 35066 13172 35072 13184
rect 33643 13144 35072 13172
rect 33643 13141 33655 13144
rect 33597 13135 33655 13141
rect 35066 13132 35072 13144
rect 35124 13132 35130 13184
rect 35268 13172 35296 13212
rect 35805 13243 35863 13249
rect 35805 13209 35817 13243
rect 35851 13240 35863 13243
rect 36078 13240 36084 13252
rect 35851 13212 36084 13240
rect 35851 13209 35863 13212
rect 35805 13203 35863 13209
rect 36078 13200 36084 13212
rect 36136 13200 36142 13252
rect 36262 13200 36268 13252
rect 36320 13200 36326 13252
rect 38470 13200 38476 13252
rect 38528 13240 38534 13252
rect 38764 13240 38792 13348
rect 40405 13345 40417 13348
rect 40451 13345 40463 13379
rect 40405 13339 40463 13345
rect 40678 13336 40684 13388
rect 40736 13336 40742 13388
rect 38933 13311 38991 13317
rect 38933 13277 38945 13311
rect 38979 13277 38991 13311
rect 38933 13271 38991 13277
rect 38528 13212 38792 13240
rect 38948 13240 38976 13271
rect 39114 13268 39120 13320
rect 39172 13268 39178 13320
rect 39206 13268 39212 13320
rect 39264 13268 39270 13320
rect 39393 13311 39451 13317
rect 39393 13277 39405 13311
rect 39439 13308 39451 13311
rect 39482 13308 39488 13320
rect 39439 13280 39488 13308
rect 39439 13277 39451 13280
rect 39393 13271 39451 13277
rect 39224 13240 39252 13268
rect 38948 13212 39252 13240
rect 38528 13200 38534 13212
rect 37274 13172 37280 13184
rect 35268 13144 37280 13172
rect 37274 13132 37280 13144
rect 37332 13132 37338 13184
rect 39114 13132 39120 13184
rect 39172 13172 39178 13184
rect 39408 13172 39436 13271
rect 39482 13268 39488 13280
rect 39540 13268 39546 13320
rect 41138 13200 41144 13252
rect 41196 13200 41202 13252
rect 39172 13144 39436 13172
rect 39577 13175 39635 13181
rect 39172 13132 39178 13144
rect 39577 13141 39589 13175
rect 39623 13172 39635 13175
rect 40218 13172 40224 13184
rect 39623 13144 40224 13172
rect 39623 13141 39635 13144
rect 39577 13135 39635 13141
rect 40218 13132 40224 13144
rect 40276 13132 40282 13184
rect 1104 13082 42504 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 42504 13082
rect 1104 13008 42504 13030
rect 4798 12928 4804 12980
rect 4856 12928 4862 12980
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6749 12971 6807 12977
rect 6749 12968 6761 12971
rect 6052 12940 6761 12968
rect 6052 12928 6058 12940
rect 6749 12937 6761 12940
rect 6795 12937 6807 12971
rect 6749 12931 6807 12937
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12968 6975 12971
rect 8018 12968 8024 12980
rect 6963 12940 8024 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 10410 12968 10416 12980
rect 9640 12940 10416 12968
rect 9640 12928 9674 12940
rect 10410 12928 10416 12940
rect 10468 12968 10474 12980
rect 16574 12968 16580 12980
rect 10468 12940 16580 12968
rect 10468 12928 10474 12940
rect 16574 12928 16580 12940
rect 16632 12968 16638 12980
rect 18138 12968 18144 12980
rect 16632 12940 18144 12968
rect 16632 12928 16638 12940
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 18414 12928 18420 12980
rect 18472 12968 18478 12980
rect 18601 12971 18659 12977
rect 18601 12968 18613 12971
rect 18472 12940 18613 12968
rect 18472 12928 18478 12940
rect 18601 12937 18613 12940
rect 18647 12937 18659 12971
rect 19886 12968 19892 12980
rect 18601 12931 18659 12937
rect 18800 12940 19892 12968
rect 3234 12900 3240 12912
rect 2990 12872 3240 12900
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 6549 12903 6607 12909
rect 6549 12869 6561 12903
rect 6595 12869 6607 12903
rect 9125 12903 9183 12909
rect 9125 12900 9137 12903
rect 6549 12863 6607 12869
rect 6840 12872 9137 12900
rect 4062 12792 4068 12844
rect 4120 12792 4126 12844
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 4614 12832 4620 12844
rect 4295 12804 4620 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5442 12832 5448 12844
rect 5399 12804 5448 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 6564 12776 6592 12863
rect 6840 12844 6868 12872
rect 9125 12869 9137 12872
rect 9171 12900 9183 12903
rect 9646 12900 9674 12928
rect 9171 12872 9674 12900
rect 9171 12869 9183 12872
rect 9125 12863 9183 12869
rect 12526 12860 12532 12912
rect 12584 12860 12590 12912
rect 13249 12903 13307 12909
rect 13249 12869 13261 12903
rect 13295 12900 13307 12903
rect 13354 12900 13360 12912
rect 13295 12872 13360 12900
rect 13295 12869 13307 12872
rect 13249 12863 13307 12869
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 13446 12860 13452 12912
rect 13504 12860 13510 12912
rect 14550 12860 14556 12912
rect 14608 12900 14614 12912
rect 14918 12900 14924 12912
rect 14608 12872 14924 12900
rect 14608 12860 14614 12872
rect 14918 12860 14924 12872
rect 14976 12900 14982 12912
rect 15102 12900 15108 12912
rect 14976 12872 15108 12900
rect 14976 12860 14982 12872
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 6822 12792 6828 12844
rect 6880 12792 6886 12844
rect 8846 12792 8852 12844
rect 8904 12792 8910 12844
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9950 12832 9956 12844
rect 9079 12804 9956 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9950 12792 9956 12804
rect 10008 12832 10014 12844
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 10008 12804 10057 12832
rect 10008 12792 10014 12804
rect 10045 12801 10057 12804
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 10199 12835 10257 12841
rect 10199 12801 10211 12835
rect 10245 12832 10257 12835
rect 10686 12832 10692 12844
rect 10245 12804 10692 12832
rect 10245 12801 10257 12804
rect 10199 12795 10257 12801
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 11238 12832 11244 12844
rect 10919 12804 11244 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 12544 12832 12572 12860
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 11940 12804 12480 12832
rect 12544 12804 12633 12832
rect 11940 12792 11946 12804
rect 1394 12724 1400 12776
rect 1452 12764 1458 12776
rect 1489 12767 1547 12773
rect 1489 12764 1501 12767
rect 1452 12736 1501 12764
rect 1452 12724 1458 12736
rect 1489 12733 1501 12736
rect 1535 12733 1547 12767
rect 1489 12727 1547 12733
rect 1504 12628 1532 12727
rect 1762 12724 1768 12776
rect 1820 12724 1826 12776
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3283 12736 3893 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 3881 12733 3893 12736
rect 3927 12764 3939 12767
rect 3970 12764 3976 12776
rect 3927 12736 3976 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5626 12764 5632 12776
rect 5123 12736 5632 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5626 12724 5632 12736
rect 5684 12764 5690 12776
rect 6546 12764 6552 12776
rect 5684 12736 6552 12764
rect 5684 12724 5690 12736
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 10413 12767 10471 12773
rect 10413 12733 10425 12767
rect 10459 12764 10471 12767
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10459 12736 10977 12764
rect 10459 12733 10471 12736
rect 10413 12727 10471 12733
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 11149 12767 11207 12773
rect 11149 12733 11161 12767
rect 11195 12764 11207 12767
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 11195 12736 11529 12764
rect 11195 12733 11207 12736
rect 11149 12727 11207 12733
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 12066 12724 12072 12776
rect 12124 12724 12130 12776
rect 12452 12764 12480 12804
rect 12621 12801 12633 12804
rect 12667 12801 12679 12835
rect 12621 12795 12679 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13722 12832 13728 12844
rect 13035 12804 13728 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 16482 12832 16488 12844
rect 15335 12804 16488 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 18800 12841 18828 12940
rect 19886 12928 19892 12940
rect 19944 12928 19950 12980
rect 22462 12928 22468 12980
rect 22520 12928 22526 12980
rect 22922 12928 22928 12980
rect 22980 12928 22986 12980
rect 28718 12968 28724 12980
rect 25056 12940 28724 12968
rect 19061 12903 19119 12909
rect 19061 12869 19073 12903
rect 19107 12900 19119 12903
rect 20162 12900 20168 12912
rect 19107 12872 20168 12900
rect 19107 12869 19119 12872
rect 19061 12863 19119 12869
rect 20162 12860 20168 12872
rect 20220 12900 20226 12912
rect 25056 12900 25084 12940
rect 28718 12928 28724 12940
rect 28776 12928 28782 12980
rect 28997 12971 29055 12977
rect 28997 12937 29009 12971
rect 29043 12968 29055 12971
rect 29086 12968 29092 12980
rect 29043 12940 29092 12968
rect 29043 12937 29055 12940
rect 28997 12931 29055 12937
rect 29086 12928 29092 12940
rect 29144 12928 29150 12980
rect 29454 12928 29460 12980
rect 29512 12928 29518 12980
rect 30466 12928 30472 12980
rect 30524 12968 30530 12980
rect 32125 12971 32183 12977
rect 32125 12968 32137 12971
rect 30524 12940 32137 12968
rect 30524 12928 30530 12940
rect 32125 12937 32137 12940
rect 32171 12937 32183 12971
rect 32125 12931 32183 12937
rect 32214 12928 32220 12980
rect 32272 12968 32278 12980
rect 32493 12971 32551 12977
rect 32493 12968 32505 12971
rect 32272 12940 32505 12968
rect 32272 12928 32278 12940
rect 32493 12937 32505 12940
rect 32539 12937 32551 12971
rect 32493 12931 32551 12937
rect 33410 12928 33416 12980
rect 33468 12928 33474 12980
rect 35342 12928 35348 12980
rect 35400 12968 35406 12980
rect 35437 12971 35495 12977
rect 35437 12968 35449 12971
rect 35400 12940 35449 12968
rect 35400 12928 35406 12940
rect 35437 12937 35449 12940
rect 35483 12968 35495 12971
rect 35526 12968 35532 12980
rect 35483 12940 35532 12968
rect 35483 12937 35495 12940
rect 35437 12931 35495 12937
rect 35526 12928 35532 12940
rect 35584 12928 35590 12980
rect 36078 12928 36084 12980
rect 36136 12968 36142 12980
rect 36173 12971 36231 12977
rect 36173 12968 36185 12971
rect 36136 12940 36185 12968
rect 36136 12928 36142 12940
rect 36173 12937 36185 12940
rect 36219 12937 36231 12971
rect 36173 12931 36231 12937
rect 36541 12971 36599 12977
rect 36541 12937 36553 12971
rect 36587 12968 36599 12971
rect 36814 12968 36820 12980
rect 36587 12940 36820 12968
rect 36587 12937 36599 12940
rect 36541 12931 36599 12937
rect 36814 12928 36820 12940
rect 36872 12928 36878 12980
rect 38562 12968 38568 12980
rect 37568 12940 38568 12968
rect 20220 12872 25084 12900
rect 20220 12860 20226 12872
rect 25130 12860 25136 12912
rect 25188 12900 25194 12912
rect 26053 12903 26111 12909
rect 26053 12900 26065 12903
rect 25188 12872 26065 12900
rect 25188 12860 25194 12872
rect 26053 12869 26065 12872
rect 26099 12900 26111 12903
rect 26142 12900 26148 12912
rect 26099 12872 26148 12900
rect 26099 12869 26111 12872
rect 26053 12863 26111 12869
rect 26142 12860 26148 12872
rect 26200 12860 26206 12912
rect 28902 12900 28908 12912
rect 27724 12872 28908 12900
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 18785 12835 18843 12841
rect 18785 12801 18797 12835
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 12529 12767 12587 12773
rect 12529 12764 12541 12767
rect 12452 12736 12541 12764
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3329 12699 3387 12705
rect 3329 12696 3341 12699
rect 2924 12668 3341 12696
rect 2924 12656 2930 12668
rect 3329 12665 3341 12668
rect 3375 12665 3387 12699
rect 3329 12659 3387 12665
rect 3418 12656 3424 12708
rect 3476 12696 3482 12708
rect 6822 12696 6828 12708
rect 3476 12668 6828 12696
rect 3476 12656 3482 12668
rect 6822 12656 6828 12668
rect 6880 12656 6886 12708
rect 8570 12656 8576 12708
rect 8628 12696 8634 12708
rect 8757 12699 8815 12705
rect 8757 12696 8769 12699
rect 8628 12668 8769 12696
rect 8628 12656 8634 12668
rect 8757 12665 8769 12668
rect 8803 12696 8815 12699
rect 9858 12696 9864 12708
rect 8803 12668 9864 12696
rect 8803 12665 8815 12668
rect 8757 12659 8815 12665
rect 9858 12656 9864 12668
rect 9916 12696 9922 12708
rect 11422 12696 11428 12708
rect 9916 12668 11428 12696
rect 9916 12656 9922 12668
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 12158 12656 12164 12708
rect 12216 12696 12222 12708
rect 12345 12699 12403 12705
rect 12345 12696 12357 12699
rect 12216 12668 12357 12696
rect 12216 12656 12222 12668
rect 12345 12665 12357 12668
rect 12391 12665 12403 12699
rect 12452 12696 12480 12736
rect 12529 12733 12541 12736
rect 12575 12733 12587 12767
rect 12529 12727 12587 12733
rect 12894 12724 12900 12776
rect 12952 12724 12958 12776
rect 15010 12724 15016 12776
rect 15068 12724 15074 12776
rect 18616 12764 18644 12795
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 19484 12804 19533 12832
rect 19484 12792 19490 12804
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 20070 12832 20076 12844
rect 19935 12804 20076 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 20070 12792 20076 12804
rect 20128 12792 20134 12844
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12832 22891 12835
rect 23566 12832 23572 12844
rect 22879 12804 23572 12832
rect 22879 12801 22891 12804
rect 22833 12795 22891 12801
rect 23566 12792 23572 12804
rect 23624 12792 23630 12844
rect 25225 12835 25283 12841
rect 25225 12801 25237 12835
rect 25271 12832 25283 12835
rect 25314 12832 25320 12844
rect 25271 12804 25320 12832
rect 25271 12801 25283 12804
rect 25225 12795 25283 12801
rect 25314 12792 25320 12804
rect 25372 12832 25378 12844
rect 27338 12832 27344 12844
rect 25372 12804 27344 12832
rect 25372 12792 25378 12804
rect 27338 12792 27344 12804
rect 27396 12792 27402 12844
rect 27433 12835 27491 12841
rect 27433 12801 27445 12835
rect 27479 12801 27491 12835
rect 27433 12795 27491 12801
rect 19334 12764 19340 12776
rect 18616 12736 19340 12764
rect 19334 12724 19340 12736
rect 19392 12724 19398 12776
rect 23109 12767 23167 12773
rect 23109 12764 23121 12767
rect 22066 12736 23121 12764
rect 13630 12696 13636 12708
rect 12452 12668 13636 12696
rect 12345 12659 12403 12665
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 17862 12656 17868 12708
rect 17920 12696 17926 12708
rect 19610 12696 19616 12708
rect 17920 12668 19616 12696
rect 17920 12656 17926 12668
rect 19610 12656 19616 12668
rect 19668 12696 19674 12708
rect 22066 12696 22094 12736
rect 23109 12733 23121 12736
rect 23155 12764 23167 12767
rect 23474 12764 23480 12776
rect 23155 12736 23480 12764
rect 23155 12733 23167 12736
rect 23109 12727 23167 12733
rect 23474 12724 23480 12736
rect 23532 12724 23538 12776
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 27448 12764 27476 12795
rect 27614 12792 27620 12844
rect 27672 12792 27678 12844
rect 27724 12841 27752 12872
rect 28902 12860 28908 12872
rect 28960 12860 28966 12912
rect 29362 12900 29368 12912
rect 29012 12872 29368 12900
rect 27709 12835 27767 12841
rect 27709 12801 27721 12835
rect 27755 12801 27767 12835
rect 27709 12795 27767 12801
rect 27985 12835 28043 12841
rect 27985 12801 27997 12835
rect 28031 12832 28043 12835
rect 28074 12832 28080 12844
rect 28031 12804 28080 12832
rect 28031 12801 28043 12804
rect 27985 12795 28043 12801
rect 28074 12792 28080 12804
rect 28132 12792 28138 12844
rect 28166 12792 28172 12844
rect 28224 12832 28230 12844
rect 28718 12832 28724 12844
rect 28224 12804 28724 12832
rect 28224 12792 28230 12804
rect 28718 12792 28724 12804
rect 28776 12792 28782 12844
rect 28813 12835 28871 12841
rect 28813 12801 28825 12835
rect 28859 12832 28871 12835
rect 29012 12832 29040 12872
rect 29362 12860 29368 12872
rect 29420 12900 29426 12912
rect 29638 12900 29644 12912
rect 29420 12872 29644 12900
rect 29420 12860 29426 12872
rect 29638 12860 29644 12872
rect 29696 12860 29702 12912
rect 30374 12860 30380 12912
rect 30432 12860 30438 12912
rect 32585 12903 32643 12909
rect 32585 12869 32597 12903
rect 32631 12900 32643 12903
rect 34422 12900 34428 12912
rect 32631 12872 34428 12900
rect 32631 12869 32643 12872
rect 32585 12863 32643 12869
rect 34422 12860 34428 12872
rect 34480 12860 34486 12912
rect 37568 12900 37596 12940
rect 38562 12928 38568 12940
rect 38620 12928 38626 12980
rect 39390 12928 39396 12980
rect 39448 12968 39454 12980
rect 40865 12971 40923 12977
rect 40865 12968 40877 12971
rect 39448 12940 40877 12968
rect 39448 12928 39454 12940
rect 40865 12937 40877 12940
rect 40911 12937 40923 12971
rect 40865 12931 40923 12937
rect 38841 12903 38899 12909
rect 35636 12872 37674 12900
rect 28859 12804 29040 12832
rect 29089 12835 29147 12841
rect 28859 12801 28871 12804
rect 28813 12795 28871 12801
rect 29089 12801 29101 12835
rect 29135 12801 29147 12835
rect 29089 12795 29147 12801
rect 28445 12767 28503 12773
rect 28445 12764 28457 12767
rect 23716 12736 27476 12764
rect 27540 12736 28457 12764
rect 23716 12724 23722 12736
rect 19668 12668 22094 12696
rect 19668 12656 19674 12668
rect 2774 12628 2780 12640
rect 1504 12600 2780 12628
rect 2774 12588 2780 12600
rect 2832 12628 2838 12640
rect 3050 12628 3056 12640
rect 2832 12600 3056 12628
rect 2832 12588 2838 12600
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 3694 12588 3700 12640
rect 3752 12628 3758 12640
rect 4065 12631 4123 12637
rect 4065 12628 4077 12631
rect 3752 12600 4077 12628
rect 3752 12588 3758 12600
rect 4065 12597 4077 12600
rect 4111 12597 4123 12631
rect 4065 12591 4123 12597
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 5166 12628 5172 12640
rect 4764 12600 5172 12628
rect 4764 12588 4770 12600
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 6454 12588 6460 12640
rect 6512 12628 6518 12640
rect 6733 12631 6791 12637
rect 6733 12628 6745 12631
rect 6512 12600 6745 12628
rect 6512 12588 6518 12600
rect 6733 12597 6745 12600
rect 6779 12597 6791 12631
rect 6733 12591 6791 12597
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 9732 12600 10517 12628
rect 9732 12588 9738 12600
rect 10505 12597 10517 12600
rect 10551 12597 10563 12631
rect 10505 12591 10563 12597
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11974 12628 11980 12640
rect 11204 12600 11980 12628
rect 11204 12588 11210 12600
rect 11974 12588 11980 12600
rect 12032 12628 12038 12640
rect 13081 12631 13139 12637
rect 13081 12628 13093 12631
rect 12032 12600 13093 12628
rect 12032 12588 12038 12600
rect 13081 12597 13093 12600
rect 13127 12597 13139 12631
rect 13081 12591 13139 12597
rect 13265 12631 13323 12637
rect 13265 12597 13277 12631
rect 13311 12628 13323 12631
rect 13538 12628 13544 12640
rect 13311 12600 13544 12628
rect 13311 12597 13323 12600
rect 13265 12591 13323 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 18969 12631 19027 12637
rect 18969 12597 18981 12631
rect 19015 12628 19027 12631
rect 19334 12628 19340 12640
rect 19015 12600 19340 12628
rect 19015 12597 19027 12600
rect 18969 12591 19027 12597
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 24854 12588 24860 12640
rect 24912 12628 24918 12640
rect 25130 12628 25136 12640
rect 24912 12600 25136 12628
rect 24912 12588 24918 12600
rect 25130 12588 25136 12600
rect 25188 12628 25194 12640
rect 27540 12628 27568 12736
rect 28445 12733 28457 12736
rect 28491 12764 28503 12767
rect 28828 12764 28856 12795
rect 28491 12736 28856 12764
rect 28491 12733 28503 12736
rect 28445 12727 28503 12733
rect 27706 12656 27712 12708
rect 27764 12696 27770 12708
rect 27893 12699 27951 12705
rect 27893 12696 27905 12699
rect 27764 12668 27905 12696
rect 27764 12656 27770 12668
rect 27893 12665 27905 12668
rect 27939 12696 27951 12699
rect 27982 12696 27988 12708
rect 27939 12668 27988 12696
rect 27939 12665 27951 12668
rect 27893 12659 27951 12665
rect 27982 12656 27988 12668
rect 28040 12656 28046 12708
rect 28166 12656 28172 12708
rect 28224 12696 28230 12708
rect 29104 12696 29132 12795
rect 29270 12792 29276 12844
rect 29328 12792 29334 12844
rect 35636 12841 35664 12872
rect 38841 12869 38853 12903
rect 38887 12900 38899 12903
rect 40494 12900 40500 12912
rect 38887 12872 40500 12900
rect 38887 12869 38899 12872
rect 38841 12863 38899 12869
rect 40494 12860 40500 12872
rect 40552 12860 40558 12912
rect 33321 12835 33379 12841
rect 33321 12801 33333 12835
rect 33367 12832 33379 12835
rect 33781 12835 33839 12841
rect 33781 12832 33793 12835
rect 33367 12804 33793 12832
rect 33367 12801 33379 12804
rect 33321 12795 33379 12801
rect 33781 12801 33793 12804
rect 33827 12801 33839 12835
rect 33781 12795 33839 12801
rect 35621 12835 35679 12841
rect 35621 12801 35633 12835
rect 35667 12801 35679 12835
rect 35621 12795 35679 12801
rect 35710 12792 35716 12844
rect 35768 12792 35774 12844
rect 36633 12835 36691 12841
rect 36633 12801 36645 12835
rect 36679 12832 36691 12835
rect 37550 12832 37556 12844
rect 36679 12804 37556 12832
rect 36679 12801 36691 12804
rect 36633 12795 36691 12801
rect 37550 12792 37556 12804
rect 37608 12792 37614 12844
rect 39485 12835 39543 12841
rect 39485 12801 39497 12835
rect 39531 12832 39543 12835
rect 40402 12832 40408 12844
rect 39531 12804 40408 12832
rect 39531 12801 39543 12804
rect 39485 12795 39543 12801
rect 31110 12724 31116 12776
rect 31168 12724 31174 12776
rect 31389 12767 31447 12773
rect 31389 12733 31401 12767
rect 31435 12764 31447 12767
rect 31570 12764 31576 12776
rect 31435 12736 31576 12764
rect 31435 12733 31447 12736
rect 31389 12727 31447 12733
rect 31570 12724 31576 12736
rect 31628 12724 31634 12776
rect 31846 12724 31852 12776
rect 31904 12764 31910 12776
rect 32769 12767 32827 12773
rect 32769 12764 32781 12767
rect 31904 12736 32781 12764
rect 31904 12724 31910 12736
rect 32769 12733 32781 12736
rect 32815 12733 32827 12767
rect 32769 12727 32827 12733
rect 28224 12668 29132 12696
rect 32784 12696 32812 12727
rect 33134 12724 33140 12776
rect 33192 12764 33198 12776
rect 33502 12764 33508 12776
rect 33192 12736 33508 12764
rect 33192 12724 33198 12736
rect 33502 12724 33508 12736
rect 33560 12724 33566 12776
rect 33594 12724 33600 12776
rect 33652 12764 33658 12776
rect 34333 12767 34391 12773
rect 34333 12764 34345 12767
rect 33652 12736 34345 12764
rect 33652 12724 33658 12736
rect 34333 12733 34345 12736
rect 34379 12733 34391 12767
rect 34333 12727 34391 12733
rect 34514 12724 34520 12776
rect 34572 12764 34578 12776
rect 35069 12767 35127 12773
rect 35069 12764 35081 12767
rect 34572 12736 35081 12764
rect 34572 12724 34578 12736
rect 35069 12733 35081 12736
rect 35115 12733 35127 12767
rect 35069 12727 35127 12733
rect 36538 12724 36544 12776
rect 36596 12764 36602 12776
rect 36725 12767 36783 12773
rect 36725 12764 36737 12767
rect 36596 12736 36737 12764
rect 36596 12724 36602 12736
rect 36725 12733 36737 12736
rect 36771 12733 36783 12767
rect 36725 12727 36783 12733
rect 37369 12767 37427 12773
rect 37369 12733 37381 12767
rect 37415 12764 37427 12767
rect 38838 12764 38844 12776
rect 37415 12736 38844 12764
rect 37415 12733 37427 12736
rect 37369 12727 37427 12733
rect 38838 12724 38844 12736
rect 38896 12724 38902 12776
rect 39117 12767 39175 12773
rect 39117 12733 39129 12767
rect 39163 12733 39175 12767
rect 39117 12727 39175 12733
rect 36556 12696 36584 12724
rect 37642 12696 37648 12708
rect 32784 12668 36584 12696
rect 36648 12668 37648 12696
rect 28224 12656 28230 12668
rect 25188 12600 27568 12628
rect 25188 12588 25194 12600
rect 27614 12588 27620 12640
rect 27672 12628 27678 12640
rect 27801 12631 27859 12637
rect 27801 12628 27813 12631
rect 27672 12600 27813 12628
rect 27672 12588 27678 12600
rect 27801 12597 27813 12600
rect 27847 12597 27859 12631
rect 27801 12591 27859 12597
rect 28626 12588 28632 12640
rect 28684 12588 28690 12640
rect 28718 12588 28724 12640
rect 28776 12628 28782 12640
rect 29641 12631 29699 12637
rect 29641 12628 29653 12631
rect 28776 12600 29653 12628
rect 28776 12588 28782 12600
rect 29641 12597 29653 12600
rect 29687 12628 29699 12631
rect 31478 12628 31484 12640
rect 29687 12600 31484 12628
rect 29687 12597 29699 12600
rect 29641 12591 29699 12597
rect 31478 12588 31484 12600
rect 31536 12588 31542 12640
rect 32306 12588 32312 12640
rect 32364 12628 32370 12640
rect 32953 12631 33011 12637
rect 32953 12628 32965 12631
rect 32364 12600 32965 12628
rect 32364 12588 32370 12600
rect 32953 12597 32965 12600
rect 32999 12597 33011 12631
rect 32953 12591 33011 12597
rect 34517 12631 34575 12637
rect 34517 12597 34529 12631
rect 34563 12628 34575 12631
rect 34606 12628 34612 12640
rect 34563 12600 34612 12628
rect 34563 12597 34575 12600
rect 34517 12591 34575 12597
rect 34606 12588 34612 12600
rect 34664 12588 34670 12640
rect 35894 12588 35900 12640
rect 35952 12628 35958 12640
rect 36648 12628 36676 12668
rect 37642 12656 37648 12668
rect 37700 12656 37706 12708
rect 35952 12600 36676 12628
rect 35952 12588 35958 12600
rect 37458 12588 37464 12640
rect 37516 12628 37522 12640
rect 38470 12628 38476 12640
rect 37516 12600 38476 12628
rect 37516 12588 37522 12600
rect 38470 12588 38476 12600
rect 38528 12628 38534 12640
rect 39132 12628 39160 12727
rect 39206 12724 39212 12776
rect 39264 12724 39270 12776
rect 39500 12696 39528 12795
rect 40402 12792 40408 12804
rect 40460 12792 40466 12844
rect 41049 12835 41107 12841
rect 41049 12801 41061 12835
rect 41095 12832 41107 12835
rect 41506 12832 41512 12844
rect 41095 12804 41512 12832
rect 41095 12801 41107 12804
rect 41049 12795 41107 12801
rect 41506 12792 41512 12804
rect 41564 12832 41570 12844
rect 42150 12832 42156 12844
rect 41564 12804 42156 12832
rect 41564 12792 41570 12804
rect 42150 12792 42156 12804
rect 42208 12792 42214 12844
rect 40678 12724 40684 12776
rect 40736 12764 40742 12776
rect 41233 12767 41291 12773
rect 41233 12764 41245 12767
rect 40736 12736 41245 12764
rect 40736 12724 40742 12736
rect 41233 12733 41245 12736
rect 41279 12733 41291 12767
rect 41233 12727 41291 12733
rect 39224 12668 39528 12696
rect 39224 12640 39252 12668
rect 38528 12600 39160 12628
rect 38528 12588 38534 12600
rect 39206 12588 39212 12640
rect 39264 12588 39270 12640
rect 39298 12588 39304 12640
rect 39356 12628 39362 12640
rect 40129 12631 40187 12637
rect 40129 12628 40141 12631
rect 39356 12600 40141 12628
rect 39356 12588 39362 12600
rect 40129 12597 40141 12600
rect 40175 12597 40187 12631
rect 40129 12591 40187 12597
rect 1104 12538 42504 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 42504 12538
rect 1104 12464 42504 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 1762 12424 1768 12436
rect 1627 12396 1768 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 5169 12427 5227 12433
rect 5169 12393 5181 12427
rect 5215 12424 5227 12427
rect 5626 12424 5632 12436
rect 5215 12396 5632 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 5718 12384 5724 12436
rect 5776 12384 5782 12436
rect 6641 12427 6699 12433
rect 6641 12393 6653 12427
rect 6687 12393 6699 12427
rect 6641 12387 6699 12393
rect 2682 12356 2688 12368
rect 2056 12328 2688 12356
rect 2056 12297 2084 12328
rect 2682 12316 2688 12328
rect 2740 12356 2746 12368
rect 3789 12359 3847 12365
rect 3789 12356 3801 12359
rect 2740 12328 3801 12356
rect 2740 12316 2746 12328
rect 3789 12325 3801 12328
rect 3835 12325 3847 12359
rect 6273 12359 6331 12365
rect 6273 12356 6285 12359
rect 3789 12319 3847 12325
rect 5644 12328 6285 12356
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12288 5043 12291
rect 5442 12288 5448 12300
rect 5031 12260 5448 12288
rect 5031 12257 5043 12260
rect 4985 12251 5043 12257
rect 5442 12248 5448 12260
rect 5500 12288 5506 12300
rect 5644 12297 5672 12328
rect 6273 12325 6285 12328
rect 6319 12356 6331 12359
rect 6656 12356 6684 12387
rect 11238 12384 11244 12436
rect 11296 12384 11302 12436
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 12066 12424 12072 12436
rect 11992 12396 12072 12424
rect 11149 12359 11207 12365
rect 6319 12328 7880 12356
rect 6319 12325 6331 12328
rect 6273 12319 6331 12325
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 5500 12260 5641 12288
rect 5500 12248 5506 12260
rect 5629 12257 5641 12260
rect 5675 12257 5687 12291
rect 5629 12251 5687 12257
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 6181 12291 6239 12297
rect 6181 12288 6193 12291
rect 5776 12260 6193 12288
rect 5776 12248 5782 12260
rect 6181 12257 6193 12260
rect 6227 12257 6239 12291
rect 6181 12251 6239 12257
rect 6730 12248 6736 12300
rect 6788 12248 6794 12300
rect 6932 12260 7696 12288
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12220 2007 12223
rect 2866 12220 2872 12232
rect 1995 12192 2872 12220
rect 1995 12189 2007 12192
rect 1949 12183 2007 12189
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12220 3203 12223
rect 3418 12220 3424 12232
rect 3191 12192 3424 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12189 3571 12223
rect 3513 12183 3571 12189
rect 2409 12155 2467 12161
rect 2409 12121 2421 12155
rect 2455 12152 2467 12155
rect 2774 12152 2780 12164
rect 2455 12124 2780 12152
rect 2455 12121 2467 12124
rect 2409 12115 2467 12121
rect 2774 12112 2780 12124
rect 2832 12112 2838 12164
rect 3528 12152 3556 12183
rect 3602 12180 3608 12232
rect 3660 12220 3666 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3660 12192 3985 12220
rect 3660 12180 3666 12192
rect 3973 12189 3985 12192
rect 4019 12220 4031 12223
rect 4062 12220 4068 12232
rect 4019 12192 4068 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4614 12220 4620 12232
rect 4212 12192 4620 12220
rect 4212 12180 4218 12192
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 5166 12180 5172 12232
rect 5224 12220 5230 12232
rect 5261 12223 5319 12229
rect 5261 12220 5273 12223
rect 5224 12192 5273 12220
rect 5224 12180 5230 12192
rect 5261 12189 5273 12192
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 4522 12152 4528 12164
rect 3528 12124 4528 12152
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 5276 12152 5304 12183
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6932 12229 6960 12260
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 5960 12192 6101 12220
rect 5960 12180 5966 12192
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6365 12223 6423 12229
rect 6365 12210 6377 12223
rect 6089 12183 6147 12189
rect 6288 12189 6377 12210
rect 6411 12210 6423 12223
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 6564 12210 6929 12220
rect 6411 12192 6929 12210
rect 6411 12189 6592 12192
rect 6288 12182 6592 12189
rect 6917 12189 6929 12192
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 5537 12155 5595 12161
rect 5537 12152 5549 12155
rect 5276 12124 5549 12152
rect 5537 12121 5549 12124
rect 5583 12152 5595 12155
rect 6288 12152 6316 12182
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7064 12192 7389 12220
rect 7064 12180 7070 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 5583 12124 6316 12152
rect 5583 12121 5595 12124
rect 5537 12115 5595 12121
rect 6638 12112 6644 12164
rect 6696 12112 6702 12164
rect 7392 12152 7420 12183
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7668 12229 7696 12260
rect 7852 12229 7880 12328
rect 11149 12325 11161 12359
rect 11195 12356 11207 12359
rect 11992 12356 12020 12396
rect 12066 12384 12072 12396
rect 12124 12424 12130 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 12124 12396 12541 12424
rect 12124 12384 12130 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 12529 12387 12587 12393
rect 13446 12384 13452 12436
rect 13504 12384 13510 12436
rect 14093 12427 14151 12433
rect 14093 12393 14105 12427
rect 14139 12424 14151 12427
rect 15010 12424 15016 12436
rect 14139 12396 15016 12424
rect 14139 12393 14151 12396
rect 14093 12387 14151 12393
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 17773 12427 17831 12433
rect 17773 12393 17785 12427
rect 17819 12424 17831 12427
rect 17819 12396 22140 12424
rect 17819 12393 17831 12396
rect 17773 12387 17831 12393
rect 11195 12328 12020 12356
rect 11195 12325 11207 12328
rect 11149 12319 11207 12325
rect 9398 12248 9404 12300
rect 9456 12248 9462 12300
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 11330 12248 11336 12300
rect 11388 12248 11394 12300
rect 7561 12223 7619 12229
rect 7561 12220 7573 12223
rect 7524 12192 7573 12220
rect 7524 12180 7530 12192
rect 7561 12189 7573 12192
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 7653 12223 7711 12229
rect 7653 12189 7665 12223
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 10778 12180 10784 12232
rect 10836 12180 10842 12232
rect 11146 12180 11152 12232
rect 11204 12180 11210 12232
rect 11348 12220 11376 12248
rect 11992 12229 12020 12328
rect 12158 12316 12164 12368
rect 12216 12356 12222 12368
rect 12345 12359 12403 12365
rect 12345 12356 12357 12359
rect 12216 12328 12357 12356
rect 12216 12316 12222 12328
rect 12345 12325 12357 12328
rect 12391 12325 12403 12359
rect 12345 12319 12403 12325
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 13464 12356 13492 12384
rect 12492 12328 13492 12356
rect 13909 12359 13967 12365
rect 12492 12316 12498 12328
rect 13909 12325 13921 12359
rect 13955 12325 13967 12359
rect 13909 12319 13967 12325
rect 16546 12328 17724 12356
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 12452 12288 12480 12316
rect 12299 12260 12480 12288
rect 12544 12260 12756 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11348 12192 11897 12220
rect 7745 12155 7803 12161
rect 7745 12152 7757 12155
rect 7392 12124 7757 12152
rect 7745 12121 7757 12124
rect 7791 12121 7803 12155
rect 7745 12115 7803 12121
rect 3326 12044 3332 12096
rect 3384 12044 3390 12096
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 4798 12084 4804 12096
rect 4755 12056 4804 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 5810 12044 5816 12096
rect 5868 12044 5874 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 6730 12084 6736 12096
rect 6595 12056 6736 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7098 12044 7104 12096
rect 7156 12044 7162 12096
rect 7469 12087 7527 12093
rect 7469 12053 7481 12087
rect 7515 12084 7527 12087
rect 8846 12084 8852 12096
rect 7515 12056 8852 12084
rect 7515 12053 7527 12056
rect 7469 12047 7527 12053
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 10796 12084 10824 12180
rect 11164 12152 11192 12180
rect 11624 12161 11652 12192
rect 11885 12189 11897 12192
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12220 12127 12223
rect 12434 12220 12440 12232
rect 12115 12192 12440 12220
rect 12115 12189 12127 12192
rect 12069 12183 12127 12189
rect 11393 12155 11451 12161
rect 11393 12152 11405 12155
rect 11164 12124 11405 12152
rect 11393 12121 11405 12124
rect 11439 12121 11451 12155
rect 11393 12115 11451 12121
rect 11609 12155 11667 12161
rect 11609 12121 11621 12155
rect 11655 12121 11667 12155
rect 11900 12152 11928 12183
rect 12434 12180 12440 12192
rect 12492 12220 12498 12232
rect 12544 12229 12572 12260
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12492 12192 12541 12220
rect 12492 12180 12498 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12728 12220 12756 12260
rect 13354 12248 13360 12300
rect 13412 12288 13418 12300
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 13412 12260 13461 12288
rect 13412 12248 13418 12260
rect 13449 12257 13461 12260
rect 13495 12257 13507 12291
rect 13924 12288 13952 12319
rect 13924 12260 14412 12288
rect 13449 12251 13507 12257
rect 13538 12220 13544 12232
rect 12728 12192 13544 12220
rect 12621 12183 12679 12189
rect 11900 12124 12434 12152
rect 11609 12115 11667 12121
rect 8996 12056 10824 12084
rect 8996 12044 9002 12056
rect 11698 12044 11704 12096
rect 11756 12044 11762 12096
rect 12406 12084 12434 12124
rect 12636 12084 12664 12183
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 14384 12229 14412 12260
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13688 12192 14289 12220
rect 13688 12180 13694 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12189 14427 12223
rect 14737 12223 14795 12229
rect 14737 12220 14749 12223
rect 14369 12183 14427 12189
rect 14476 12192 14749 12220
rect 12802 12112 12808 12164
rect 12860 12112 12866 12164
rect 13556 12152 13584 12180
rect 14476 12152 14504 12192
rect 14737 12189 14749 12192
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 15896 12192 16405 12220
rect 15896 12180 15902 12192
rect 16393 12189 16405 12192
rect 16439 12220 16451 12223
rect 16546 12220 16574 12328
rect 16439 12192 16574 12220
rect 16669 12223 16727 12229
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 16669 12189 16681 12223
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12220 16911 12223
rect 16899 12192 17540 12220
rect 16899 12189 16911 12192
rect 16853 12183 16911 12189
rect 13556 12124 14504 12152
rect 14645 12155 14703 12161
rect 14645 12121 14657 12155
rect 14691 12121 14703 12155
rect 14645 12115 14703 12121
rect 12406 12056 12664 12084
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 14550 12084 14556 12096
rect 12952 12056 14556 12084
rect 12952 12044 12958 12056
rect 14550 12044 14556 12056
rect 14608 12084 14614 12096
rect 14660 12084 14688 12115
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 16684 12152 16712 12183
rect 16945 12155 17003 12161
rect 16945 12152 16957 12155
rect 16632 12124 16957 12152
rect 16632 12112 16638 12124
rect 16945 12121 16957 12124
rect 16991 12121 17003 12155
rect 17512 12152 17540 12192
rect 17586 12180 17592 12232
rect 17644 12180 17650 12232
rect 17696 12229 17724 12328
rect 20162 12316 20168 12368
rect 20220 12316 20226 12368
rect 22112 12356 22140 12396
rect 22186 12384 22192 12436
rect 22244 12384 22250 12436
rect 23198 12384 23204 12436
rect 23256 12424 23262 12436
rect 24121 12427 24179 12433
rect 24121 12424 24133 12427
rect 23256 12396 24133 12424
rect 23256 12384 23262 12396
rect 24121 12393 24133 12396
rect 24167 12424 24179 12427
rect 24302 12424 24308 12436
rect 24167 12396 24308 12424
rect 24167 12393 24179 12396
rect 24121 12387 24179 12393
rect 24302 12384 24308 12396
rect 24360 12424 24366 12436
rect 24360 12396 25176 12424
rect 24360 12384 24366 12396
rect 23658 12356 23664 12368
rect 22112 12328 23664 12356
rect 23658 12316 23664 12328
rect 23716 12316 23722 12368
rect 20349 12291 20407 12297
rect 20349 12257 20361 12291
rect 20395 12288 20407 12291
rect 21450 12288 21456 12300
rect 20395 12260 21456 12288
rect 20395 12257 20407 12260
rect 20349 12251 20407 12257
rect 21450 12248 21456 12260
rect 21508 12288 21514 12300
rect 21508 12260 22600 12288
rect 21508 12248 21514 12260
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 17862 12180 17868 12232
rect 17920 12180 17926 12232
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19337 12223 19395 12229
rect 19337 12220 19349 12223
rect 19208 12192 19349 12220
rect 19208 12180 19214 12192
rect 19337 12189 19349 12192
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 20254 12180 20260 12232
rect 20312 12180 20318 12232
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22370 12220 22376 12232
rect 22143 12192 22376 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22572 12220 22600 12260
rect 22646 12248 22652 12300
rect 22704 12248 22710 12300
rect 22833 12291 22891 12297
rect 22833 12257 22845 12291
rect 22879 12288 22891 12291
rect 22922 12288 22928 12300
rect 22879 12260 22928 12288
rect 22879 12257 22891 12260
rect 22833 12251 22891 12257
rect 22922 12248 22928 12260
rect 22980 12288 22986 12300
rect 22980 12260 23888 12288
rect 22980 12248 22986 12260
rect 23569 12223 23627 12229
rect 23569 12220 23581 12223
rect 22572 12192 23581 12220
rect 23569 12189 23581 12192
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 17880 12152 17908 12180
rect 17512 12124 17908 12152
rect 16945 12115 17003 12121
rect 19794 12112 19800 12164
rect 19852 12152 19858 12164
rect 20162 12152 20168 12164
rect 19852 12124 20168 12152
rect 19852 12112 19858 12124
rect 20162 12112 20168 12124
rect 20220 12152 20226 12164
rect 21821 12155 21879 12161
rect 20220 12124 20654 12152
rect 20220 12112 20226 12124
rect 21821 12121 21833 12155
rect 21867 12152 21879 12155
rect 22186 12152 22192 12164
rect 21867 12124 22192 12152
rect 21867 12121 21879 12124
rect 21821 12115 21879 12121
rect 22186 12112 22192 12124
rect 22244 12112 22250 12164
rect 22278 12112 22284 12164
rect 22336 12152 22342 12164
rect 22738 12152 22744 12164
rect 22336 12124 22744 12152
rect 22336 12112 22342 12124
rect 22738 12112 22744 12124
rect 22796 12112 22802 12164
rect 23860 12161 23888 12260
rect 24946 12248 24952 12300
rect 25004 12248 25010 12300
rect 25148 12297 25176 12396
rect 25222 12384 25228 12436
rect 25280 12424 25286 12436
rect 26418 12424 26424 12436
rect 25280 12396 26424 12424
rect 25280 12384 25286 12396
rect 26418 12384 26424 12396
rect 26476 12384 26482 12436
rect 26970 12384 26976 12436
rect 27028 12424 27034 12436
rect 29273 12427 29331 12433
rect 27028 12396 29224 12424
rect 27028 12384 27034 12396
rect 29196 12356 29224 12396
rect 29273 12393 29285 12427
rect 29319 12424 29331 12427
rect 29546 12424 29552 12436
rect 29319 12396 29552 12424
rect 29319 12393 29331 12396
rect 29273 12387 29331 12393
rect 29546 12384 29552 12396
rect 29604 12384 29610 12436
rect 30653 12427 30711 12433
rect 30653 12393 30665 12427
rect 30699 12424 30711 12427
rect 31110 12424 31116 12436
rect 30699 12396 31116 12424
rect 30699 12393 30711 12396
rect 30653 12387 30711 12393
rect 31110 12384 31116 12396
rect 31168 12384 31174 12436
rect 31312 12396 32536 12424
rect 31312 12356 31340 12396
rect 29196 12328 31340 12356
rect 32508 12356 32536 12396
rect 32950 12384 32956 12436
rect 33008 12384 33014 12436
rect 34333 12427 34391 12433
rect 34333 12393 34345 12427
rect 34379 12424 34391 12427
rect 34698 12424 34704 12436
rect 34379 12396 34704 12424
rect 34379 12393 34391 12396
rect 34333 12387 34391 12393
rect 34698 12384 34704 12396
rect 34756 12384 34762 12436
rect 38378 12384 38384 12436
rect 38436 12424 38442 12436
rect 39390 12424 39396 12436
rect 38436 12396 39396 12424
rect 38436 12384 38442 12396
rect 39390 12384 39396 12396
rect 39448 12384 39454 12436
rect 39482 12384 39488 12436
rect 39540 12424 39546 12436
rect 39540 12396 40540 12424
rect 39540 12384 39546 12396
rect 34517 12359 34575 12365
rect 34517 12356 34529 12359
rect 32508 12328 34529 12356
rect 34517 12325 34529 12328
rect 34563 12325 34575 12359
rect 35986 12356 35992 12368
rect 34517 12319 34575 12325
rect 35360 12328 35992 12356
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12288 25191 12291
rect 25866 12288 25872 12300
rect 25179 12260 25872 12288
rect 25179 12257 25191 12260
rect 25133 12251 25191 12257
rect 25866 12248 25872 12260
rect 25924 12248 25930 12300
rect 27341 12291 27399 12297
rect 27341 12257 27353 12291
rect 27387 12288 27399 12291
rect 27982 12288 27988 12300
rect 27387 12260 27988 12288
rect 27387 12257 27399 12260
rect 27341 12251 27399 12257
rect 24118 12180 24124 12232
rect 24176 12220 24182 12232
rect 24762 12220 24768 12232
rect 24176 12192 24768 12220
rect 24176 12180 24182 12192
rect 24762 12180 24768 12192
rect 24820 12220 24826 12232
rect 25774 12220 25780 12232
rect 24820 12192 25780 12220
rect 24820 12180 24826 12192
rect 25774 12180 25780 12192
rect 25832 12180 25838 12232
rect 26050 12180 26056 12232
rect 26108 12180 26114 12232
rect 26142 12180 26148 12232
rect 26200 12220 26206 12232
rect 26605 12223 26663 12229
rect 26605 12220 26617 12223
rect 26200 12192 26617 12220
rect 26200 12180 26206 12192
rect 26605 12189 26617 12192
rect 26651 12220 26663 12223
rect 27356 12220 27384 12251
rect 27982 12248 27988 12260
rect 28040 12248 28046 12300
rect 29089 12291 29147 12297
rect 29089 12288 29101 12291
rect 29012 12260 29101 12288
rect 26651 12192 27384 12220
rect 26651 12189 26663 12192
rect 26605 12183 26663 12189
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 26510 12152 26516 12164
rect 23891 12124 26516 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 26510 12112 26516 12124
rect 26568 12112 26574 12164
rect 27617 12155 27675 12161
rect 27617 12121 27629 12155
rect 27663 12121 27675 12155
rect 28902 12152 28908 12164
rect 28842 12124 28908 12152
rect 27617 12115 27675 12121
rect 14608 12056 14688 12084
rect 14608 12044 14614 12056
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 16209 12087 16267 12093
rect 16209 12084 16221 12087
rect 16172 12056 16221 12084
rect 16172 12044 16178 12056
rect 16209 12053 16221 12056
rect 16255 12053 16267 12087
rect 16209 12047 16267 12053
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 19576 12056 19993 12084
rect 19576 12044 19582 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 19981 12047 20039 12053
rect 20070 12044 20076 12096
rect 20128 12084 20134 12096
rect 22462 12084 22468 12096
rect 20128 12056 22468 12084
rect 20128 12044 20134 12056
rect 22462 12044 22468 12056
rect 22520 12044 22526 12096
rect 22557 12087 22615 12093
rect 22557 12053 22569 12087
rect 22603 12084 22615 12087
rect 23017 12087 23075 12093
rect 23017 12084 23029 12087
rect 22603 12056 23029 12084
rect 22603 12053 22615 12056
rect 22557 12047 22615 12053
rect 23017 12053 23029 12056
rect 23063 12053 23075 12087
rect 23017 12047 23075 12053
rect 24486 12044 24492 12096
rect 24544 12044 24550 12096
rect 24857 12087 24915 12093
rect 24857 12053 24869 12087
rect 24903 12084 24915 12087
rect 25501 12087 25559 12093
rect 25501 12084 25513 12087
rect 24903 12056 25513 12084
rect 24903 12053 24915 12056
rect 24857 12047 24915 12053
rect 25501 12053 25513 12056
rect 25547 12053 25559 12087
rect 27632 12084 27660 12115
rect 28902 12112 28908 12124
rect 28960 12112 28966 12164
rect 29012 12152 29040 12260
rect 29089 12257 29101 12260
rect 29135 12257 29147 12291
rect 29089 12251 29147 12257
rect 29454 12248 29460 12300
rect 29512 12288 29518 12300
rect 30285 12291 30343 12297
rect 30285 12288 30297 12291
rect 29512 12260 30297 12288
rect 29512 12248 29518 12260
rect 30285 12257 30297 12260
rect 30331 12257 30343 12291
rect 30285 12251 30343 12257
rect 31662 12248 31668 12300
rect 31720 12288 31726 12300
rect 32861 12291 32919 12297
rect 31720 12260 32628 12288
rect 31720 12248 31726 12260
rect 32600 12232 32628 12260
rect 32861 12257 32873 12291
rect 32907 12288 32919 12291
rect 33318 12288 33324 12300
rect 32907 12260 33324 12288
rect 32907 12257 32919 12260
rect 32861 12251 32919 12257
rect 33318 12248 33324 12260
rect 33376 12248 33382 12300
rect 33686 12248 33692 12300
rect 33744 12248 33750 12300
rect 33870 12248 33876 12300
rect 33928 12248 33934 12300
rect 33962 12248 33968 12300
rect 34020 12288 34026 12300
rect 34149 12291 34207 12297
rect 34149 12288 34161 12291
rect 34020 12260 34161 12288
rect 34020 12248 34026 12260
rect 34149 12257 34161 12260
rect 34195 12257 34207 12291
rect 34606 12288 34612 12300
rect 34149 12251 34207 12257
rect 34256 12260 34612 12288
rect 29178 12180 29184 12232
rect 29236 12180 29242 12232
rect 29270 12180 29276 12232
rect 29328 12220 29334 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29328 12192 29745 12220
rect 29328 12180 29334 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 30190 12180 30196 12232
rect 30248 12220 30254 12232
rect 30469 12223 30527 12229
rect 30469 12220 30481 12223
rect 30248 12192 30481 12220
rect 30248 12180 30254 12192
rect 30469 12189 30481 12192
rect 30515 12189 30527 12223
rect 30469 12183 30527 12189
rect 32582 12180 32588 12232
rect 32640 12180 32646 12232
rect 32950 12180 32956 12232
rect 33008 12180 33014 12232
rect 33597 12223 33655 12229
rect 33597 12189 33609 12223
rect 33643 12220 33655 12223
rect 34256 12220 34284 12260
rect 34606 12248 34612 12260
rect 34664 12248 34670 12300
rect 35360 12297 35388 12328
rect 35986 12316 35992 12328
rect 36044 12316 36050 12368
rect 38948 12328 39528 12356
rect 35345 12291 35403 12297
rect 35345 12257 35357 12291
rect 35391 12257 35403 12291
rect 35345 12251 35403 12257
rect 35529 12291 35587 12297
rect 35529 12257 35541 12291
rect 35575 12288 35587 12291
rect 35894 12288 35900 12300
rect 35575 12260 35900 12288
rect 35575 12257 35587 12260
rect 35529 12251 35587 12257
rect 35894 12248 35900 12260
rect 35952 12248 35958 12300
rect 36906 12288 36912 12300
rect 36280 12260 36912 12288
rect 33643 12192 34284 12220
rect 34333 12223 34391 12229
rect 33643 12189 33655 12192
rect 33597 12183 33655 12189
rect 34333 12189 34345 12223
rect 34379 12220 34391 12223
rect 36280 12220 36308 12260
rect 36906 12248 36912 12260
rect 36964 12248 36970 12300
rect 37458 12248 37464 12300
rect 37516 12288 37522 12300
rect 38105 12291 38163 12297
rect 38105 12288 38117 12291
rect 37516 12260 38117 12288
rect 37516 12248 37522 12260
rect 38105 12257 38117 12260
rect 38151 12257 38163 12291
rect 38105 12251 38163 12257
rect 38838 12248 38844 12300
rect 38896 12288 38902 12300
rect 38948 12297 38976 12328
rect 38933 12291 38991 12297
rect 38933 12288 38945 12291
rect 38896 12260 38945 12288
rect 38896 12248 38902 12260
rect 38933 12257 38945 12260
rect 38979 12257 38991 12291
rect 38933 12251 38991 12257
rect 39022 12248 39028 12300
rect 39080 12288 39086 12300
rect 39080 12260 39432 12288
rect 39080 12248 39086 12260
rect 34379 12192 36308 12220
rect 34379 12189 34391 12192
rect 34333 12183 34391 12189
rect 36354 12180 36360 12232
rect 36412 12180 36418 12232
rect 37182 12180 37188 12232
rect 37240 12180 37246 12232
rect 37550 12180 37556 12232
rect 37608 12220 37614 12232
rect 39206 12229 39212 12232
rect 38381 12223 38439 12229
rect 38381 12220 38393 12223
rect 37608 12192 38393 12220
rect 37608 12180 37614 12192
rect 38381 12189 38393 12192
rect 38427 12189 38439 12223
rect 38381 12183 38439 12189
rect 39163 12223 39212 12229
rect 39163 12189 39175 12223
rect 39209 12189 39212 12223
rect 39163 12183 39212 12189
rect 30101 12155 30159 12161
rect 30101 12152 30113 12155
rect 29012 12124 30113 12152
rect 30101 12121 30113 12124
rect 30147 12152 30159 12155
rect 31018 12152 31024 12164
rect 30147 12124 31024 12152
rect 30147 12121 30159 12124
rect 30101 12115 30159 12121
rect 31018 12112 31024 12124
rect 31076 12112 31082 12164
rect 31878 12124 32260 12152
rect 28626 12084 28632 12096
rect 27632 12056 28632 12084
rect 25501 12047 25559 12053
rect 28626 12044 28632 12056
rect 28684 12044 28690 12096
rect 28920 12084 28948 12112
rect 30374 12084 30380 12096
rect 28920 12056 30380 12084
rect 30374 12044 30380 12056
rect 30432 12044 30438 12096
rect 30834 12044 30840 12096
rect 30892 12044 30898 12096
rect 32232 12084 32260 12124
rect 32306 12112 32312 12164
rect 32364 12112 32370 12164
rect 32674 12112 32680 12164
rect 32732 12112 32738 12164
rect 34057 12155 34115 12161
rect 34057 12152 34069 12155
rect 33152 12124 34069 12152
rect 32858 12084 32864 12096
rect 32232 12056 32864 12084
rect 32858 12044 32864 12056
rect 32916 12084 32922 12096
rect 33042 12084 33048 12096
rect 32916 12056 33048 12084
rect 32916 12044 32922 12056
rect 33042 12044 33048 12056
rect 33100 12044 33106 12096
rect 33152 12093 33180 12124
rect 34057 12121 34069 12124
rect 34103 12121 34115 12155
rect 34057 12115 34115 12121
rect 35342 12112 35348 12164
rect 35400 12152 35406 12164
rect 35526 12152 35532 12164
rect 35400 12124 35532 12152
rect 35400 12112 35406 12124
rect 35526 12112 35532 12124
rect 35584 12112 35590 12164
rect 37366 12112 37372 12164
rect 37424 12152 37430 12164
rect 38194 12152 38200 12164
rect 37424 12124 38200 12152
rect 37424 12112 37430 12124
rect 38194 12112 38200 12124
rect 38252 12112 38258 12164
rect 38396 12152 38424 12183
rect 39206 12180 39212 12183
rect 39264 12180 39270 12232
rect 39404 12229 39432 12260
rect 39500 12229 39528 12328
rect 39574 12316 39580 12368
rect 39632 12316 39638 12368
rect 39669 12359 39727 12365
rect 39669 12325 39681 12359
rect 39715 12356 39727 12359
rect 40512 12356 40540 12396
rect 41509 12359 41567 12365
rect 41509 12356 41521 12359
rect 39715 12328 40448 12356
rect 40512 12328 41521 12356
rect 39715 12325 39727 12328
rect 39669 12319 39727 12325
rect 39592 12288 39620 12316
rect 39853 12291 39911 12297
rect 39853 12288 39865 12291
rect 39592 12260 39865 12288
rect 39853 12257 39865 12260
rect 39899 12257 39911 12291
rect 39853 12251 39911 12257
rect 39942 12248 39948 12300
rect 40000 12288 40006 12300
rect 40000 12260 40356 12288
rect 40000 12248 40006 12260
rect 39389 12223 39447 12229
rect 39389 12189 39401 12223
rect 39435 12189 39447 12223
rect 39389 12183 39447 12189
rect 39485 12223 39543 12229
rect 39485 12189 39497 12223
rect 39531 12189 39543 12223
rect 39485 12183 39543 12189
rect 39574 12180 39580 12232
rect 39632 12220 39638 12232
rect 40129 12223 40187 12229
rect 40129 12220 40141 12223
rect 39632 12192 40141 12220
rect 39632 12180 39638 12192
rect 40129 12189 40141 12192
rect 40175 12189 40187 12223
rect 40129 12183 40187 12189
rect 40218 12180 40224 12232
rect 40276 12180 40282 12232
rect 40328 12229 40356 12260
rect 40313 12223 40371 12229
rect 40313 12189 40325 12223
rect 40359 12189 40371 12223
rect 40420 12220 40448 12328
rect 41509 12325 41521 12328
rect 41555 12325 41567 12359
rect 41509 12319 41567 12325
rect 40494 12248 40500 12300
rect 40552 12248 40558 12300
rect 40678 12248 40684 12300
rect 40736 12288 40742 12300
rect 40736 12260 41368 12288
rect 40736 12248 40742 12260
rect 41340 12229 41368 12260
rect 41141 12223 41199 12229
rect 41141 12220 41153 12223
rect 40420 12192 41153 12220
rect 40313 12183 40371 12189
rect 41141 12189 41153 12192
rect 41187 12189 41199 12223
rect 41141 12183 41199 12189
rect 41325 12223 41383 12229
rect 41325 12189 41337 12223
rect 41371 12189 41383 12223
rect 41325 12183 41383 12189
rect 41506 12180 41512 12232
rect 41564 12180 41570 12232
rect 38930 12152 38936 12164
rect 38396 12124 38936 12152
rect 38930 12112 38936 12124
rect 38988 12112 38994 12164
rect 39298 12112 39304 12164
rect 39356 12112 39362 12164
rect 39758 12112 39764 12164
rect 39816 12152 39822 12164
rect 39991 12155 40049 12161
rect 39991 12152 40003 12155
rect 39816 12124 40003 12152
rect 39816 12112 39822 12124
rect 39991 12121 40003 12124
rect 40037 12121 40049 12155
rect 39991 12115 40049 12121
rect 33137 12087 33195 12093
rect 33137 12053 33149 12087
rect 33183 12053 33195 12087
rect 33137 12047 33195 12053
rect 33226 12044 33232 12096
rect 33284 12044 33290 12096
rect 33318 12044 33324 12096
rect 33376 12084 33382 12096
rect 34146 12084 34152 12096
rect 33376 12056 34152 12084
rect 33376 12044 33382 12056
rect 34146 12044 34152 12056
rect 34204 12044 34210 12096
rect 34790 12044 34796 12096
rect 34848 12084 34854 12096
rect 34885 12087 34943 12093
rect 34885 12084 34897 12087
rect 34848 12056 34897 12084
rect 34848 12044 34854 12056
rect 34885 12053 34897 12056
rect 34931 12053 34943 12087
rect 34885 12047 34943 12053
rect 35253 12087 35311 12093
rect 35253 12053 35265 12087
rect 35299 12084 35311 12087
rect 35805 12087 35863 12093
rect 35805 12084 35817 12087
rect 35299 12056 35817 12084
rect 35299 12053 35311 12056
rect 35253 12047 35311 12053
rect 35805 12053 35817 12056
rect 35851 12053 35863 12087
rect 35805 12047 35863 12053
rect 36541 12087 36599 12093
rect 36541 12053 36553 12087
rect 36587 12084 36599 12087
rect 36722 12084 36728 12096
rect 36587 12056 36728 12084
rect 36587 12053 36599 12056
rect 36541 12047 36599 12053
rect 36722 12044 36728 12056
rect 36780 12044 36786 12096
rect 37918 12044 37924 12096
rect 37976 12084 37982 12096
rect 39206 12084 39212 12096
rect 37976 12056 39212 12084
rect 37976 12044 37982 12056
rect 39206 12044 39212 12056
rect 39264 12044 39270 12096
rect 40586 12044 40592 12096
rect 40644 12044 40650 12096
rect 1104 11994 42504 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 42504 11994
rect 1104 11920 42504 11942
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11849 3295 11883
rect 3237 11843 3295 11849
rect 3252 11812 3280 11843
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4357 11883 4415 11889
rect 4357 11880 4369 11883
rect 4028 11852 4369 11880
rect 4028 11840 4034 11852
rect 4357 11849 4369 11852
rect 4403 11849 4415 11883
rect 4357 11843 4415 11849
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 4801 11883 4859 11889
rect 4801 11880 4813 11883
rect 4764 11852 4813 11880
rect 4764 11840 4770 11852
rect 4801 11849 4813 11852
rect 4847 11880 4859 11883
rect 5350 11880 5356 11892
rect 4847 11852 5356 11880
rect 4847 11849 4859 11852
rect 4801 11843 4859 11849
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5902 11840 5908 11892
rect 5960 11880 5966 11892
rect 6546 11880 6552 11892
rect 5960 11852 6552 11880
rect 5960 11840 5966 11852
rect 6546 11840 6552 11852
rect 6604 11880 6610 11892
rect 6917 11883 6975 11889
rect 6917 11880 6929 11883
rect 6604 11852 6929 11880
rect 6604 11840 6610 11852
rect 6917 11849 6929 11852
rect 6963 11849 6975 11883
rect 6917 11843 6975 11849
rect 7466 11840 7472 11892
rect 7524 11840 7530 11892
rect 8294 11880 8300 11892
rect 8128 11852 8300 11880
rect 4154 11812 4160 11824
rect 3252 11784 4160 11812
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 4617 11815 4675 11821
rect 4617 11781 4629 11815
rect 4663 11812 4675 11815
rect 5442 11812 5448 11824
rect 4663 11784 5448 11812
rect 4663 11781 4675 11784
rect 4617 11775 4675 11781
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 5810 11772 5816 11824
rect 5868 11812 5874 11824
rect 6641 11815 6699 11821
rect 6641 11812 6653 11815
rect 5868 11784 6653 11812
rect 5868 11772 5874 11784
rect 6641 11781 6653 11784
rect 6687 11812 6699 11815
rect 6730 11812 6736 11824
rect 6687 11784 6736 11812
rect 6687 11781 6699 11784
rect 6641 11775 6699 11781
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 7374 11772 7380 11824
rect 7432 11812 7438 11824
rect 7929 11815 7987 11821
rect 7929 11812 7941 11815
rect 7432 11784 7941 11812
rect 7432 11772 7438 11784
rect 7929 11781 7941 11784
rect 7975 11781 7987 11815
rect 7929 11775 7987 11781
rect 3234 11744 3240 11756
rect 2898 11716 3240 11744
rect 3234 11704 3240 11716
rect 3292 11704 3298 11756
rect 3510 11704 3516 11756
rect 3568 11704 3574 11756
rect 4798 11704 4804 11756
rect 4856 11744 4862 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4856 11716 4905 11744
rect 4856 11704 4862 11716
rect 4893 11713 4905 11716
rect 4939 11744 4951 11747
rect 5258 11744 5264 11756
rect 4939 11716 5264 11744
rect 4939 11713 4951 11716
rect 4893 11707 4951 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 6089 11747 6147 11753
rect 6089 11713 6101 11747
rect 6135 11713 6147 11747
rect 6089 11707 6147 11713
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11744 6515 11747
rect 6546 11744 6552 11756
rect 6503 11716 6552 11744
rect 6503 11713 6515 11716
rect 6457 11707 6515 11713
rect 1486 11636 1492 11688
rect 1544 11636 1550 11688
rect 1762 11636 1768 11688
rect 1820 11636 1826 11688
rect 4522 11636 4528 11688
rect 4580 11676 4586 11688
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 4580 11648 5733 11676
rect 4580 11636 4586 11648
rect 5721 11645 5733 11648
rect 5767 11645 5779 11679
rect 6104 11676 6132 11707
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 8128 11753 8156 11852
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 8444 11852 9996 11880
rect 8444 11840 8450 11852
rect 8404 11812 8432 11840
rect 8312 11784 8432 11812
rect 8312 11753 8340 11784
rect 8570 11772 8576 11824
rect 8628 11772 8634 11824
rect 8665 11815 8723 11821
rect 8665 11781 8677 11815
rect 8711 11812 8723 11815
rect 9033 11815 9091 11821
rect 9033 11812 9045 11815
rect 8711 11784 9045 11812
rect 8711 11781 8723 11784
rect 8665 11775 8723 11781
rect 9033 11781 9045 11784
rect 9079 11781 9091 11815
rect 9033 11775 9091 11781
rect 9490 11772 9496 11824
rect 9548 11812 9554 11824
rect 9968 11812 9996 11852
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 12066 11880 12072 11892
rect 10100 11852 12072 11880
rect 10100 11840 10106 11852
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12434 11880 12440 11892
rect 12207 11852 12440 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12802 11840 12808 11892
rect 12860 11840 12866 11892
rect 12897 11883 12955 11889
rect 12897 11849 12909 11883
rect 12943 11880 12955 11883
rect 13354 11880 13360 11892
rect 12943 11852 13360 11880
rect 12943 11849 12955 11852
rect 12897 11843 12955 11849
rect 12526 11812 12532 11824
rect 9548 11784 9904 11812
rect 9968 11784 12204 11812
rect 9548 11772 9554 11784
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 6880 11716 7113 11744
rect 6880 11704 6886 11716
rect 7101 11713 7113 11716
rect 7147 11744 7159 11747
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 7147 11716 7665 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 7653 11713 7665 11716
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11713 8447 11747
rect 8389 11707 8447 11713
rect 7006 11676 7012 11688
rect 6104 11648 7012 11676
rect 5721 11639 5779 11645
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7340 11648 7757 11676
rect 7340 11636 7346 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 8404 11676 8432 11707
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 8904 11716 9781 11744
rect 8904 11704 8910 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9876 11744 9904 11784
rect 12176 11756 12204 11784
rect 12268 11784 12532 11812
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9876 11716 9965 11744
rect 9769 11707 9827 11713
rect 9953 11713 9965 11716
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 7745 11639 7803 11645
rect 8312 11648 8432 11676
rect 8772 11676 8800 11704
rect 9490 11676 9496 11688
rect 8772 11648 9496 11676
rect 3418 11568 3424 11620
rect 3476 11608 3482 11620
rect 8312 11617 8340 11648
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 10428 11676 10456 11707
rect 10686 11676 10692 11688
rect 9732 11648 10692 11676
rect 9732 11636 9738 11648
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 11882 11636 11888 11688
rect 11940 11636 11946 11688
rect 11992 11676 12020 11707
rect 12158 11704 12164 11756
rect 12216 11704 12222 11756
rect 12268 11753 12296 11784
rect 12526 11772 12532 11784
rect 12584 11812 12590 11824
rect 12912 11812 12940 11843
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 15160 11852 17356 11880
rect 15160 11840 15166 11852
rect 13170 11812 13176 11824
rect 12584 11784 12940 11812
rect 13004 11784 13176 11812
rect 12584 11772 12590 11784
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12618 11704 12624 11756
rect 12676 11704 12682 11756
rect 12360 11676 12388 11704
rect 11992 11648 12388 11676
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 13004 11676 13032 11784
rect 13170 11772 13176 11784
rect 13228 11812 13234 11824
rect 13817 11815 13875 11821
rect 13817 11812 13829 11815
rect 13228 11784 13829 11812
rect 13228 11772 13234 11784
rect 13817 11781 13829 11784
rect 13863 11812 13875 11815
rect 13998 11812 14004 11824
rect 13863 11784 14004 11812
rect 13863 11781 13875 11784
rect 13817 11775 13875 11781
rect 13998 11772 14004 11784
rect 14056 11772 14062 11824
rect 16485 11815 16543 11821
rect 16485 11781 16497 11815
rect 16531 11812 16543 11815
rect 16945 11815 17003 11821
rect 16945 11812 16957 11815
rect 16531 11784 16957 11812
rect 16531 11781 16543 11784
rect 16485 11775 16543 11781
rect 16945 11781 16957 11784
rect 16991 11781 17003 11815
rect 17328 11812 17356 11852
rect 19150 11840 19156 11892
rect 19208 11840 19214 11892
rect 19613 11883 19671 11889
rect 19613 11849 19625 11883
rect 19659 11880 19671 11883
rect 19978 11880 19984 11892
rect 19659 11852 19984 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 22370 11840 22376 11892
rect 22428 11880 22434 11892
rect 26142 11880 26148 11892
rect 22428 11852 26148 11880
rect 22428 11840 22434 11852
rect 17328 11784 17434 11812
rect 16945 11775 17003 11781
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 21085 11815 21143 11821
rect 21085 11812 21097 11815
rect 20772 11784 21097 11812
rect 20772 11772 20778 11784
rect 21085 11781 21097 11784
rect 21131 11781 21143 11815
rect 22922 11812 22928 11824
rect 21085 11775 21143 11781
rect 21284 11784 22928 11812
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13446 11744 13452 11756
rect 13127 11716 13452 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 12483 11648 13032 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 4617 11611 4675 11617
rect 4617 11608 4629 11611
rect 3476 11580 4629 11608
rect 3476 11568 3482 11580
rect 4617 11577 4629 11580
rect 4663 11577 4675 11611
rect 4617 11571 4675 11577
rect 8297 11611 8355 11617
rect 8297 11577 8309 11611
rect 8343 11577 8355 11611
rect 10321 11611 10379 11617
rect 10321 11608 10333 11611
rect 8297 11571 8355 11577
rect 9876 11580 10333 11608
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4120 11512 4353 11540
rect 4120 11500 4126 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 4525 11543 4583 11549
rect 4525 11509 4537 11543
rect 4571 11540 4583 11543
rect 5626 11540 5632 11552
rect 4571 11512 5632 11540
rect 4571 11509 4583 11512
rect 4525 11503 4583 11509
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 6871 11512 7389 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 7377 11509 7389 11512
rect 7423 11540 7435 11543
rect 7466 11540 7472 11552
rect 7423 11512 7472 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 7466 11500 7472 11512
rect 7524 11540 7530 11552
rect 7653 11543 7711 11549
rect 7653 11540 7665 11543
rect 7524 11512 7665 11540
rect 7524 11500 7530 11512
rect 7653 11509 7665 11512
rect 7699 11509 7711 11543
rect 7653 11503 7711 11509
rect 8938 11500 8944 11552
rect 8996 11500 9002 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9876 11540 9904 11580
rect 10321 11577 10333 11580
rect 10367 11577 10379 11611
rect 11900 11608 11928 11636
rect 10321 11571 10379 11577
rect 11808 11580 11928 11608
rect 11977 11611 12035 11617
rect 9088 11512 9904 11540
rect 9088 11500 9094 11512
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 11808 11540 11836 11580
rect 11977 11577 11989 11611
rect 12023 11608 12035 11611
rect 12250 11608 12256 11620
rect 12023 11580 12256 11608
rect 12023 11577 12035 11580
rect 11977 11571 12035 11577
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 10192 11512 11836 11540
rect 10192 11500 10198 11512
rect 11882 11500 11888 11552
rect 11940 11540 11946 11552
rect 12452 11540 12480 11639
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 13228 11648 13277 11676
rect 13228 11636 13234 11648
rect 13265 11645 13277 11648
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 13354 11636 13360 11688
rect 13412 11676 13418 11688
rect 13556 11676 13584 11707
rect 13412 11648 13584 11676
rect 13412 11636 13418 11648
rect 12802 11568 12808 11620
rect 12860 11608 12866 11620
rect 13648 11608 13676 11707
rect 14550 11704 14556 11756
rect 14608 11704 14614 11756
rect 15838 11704 15844 11756
rect 15896 11744 15902 11756
rect 16117 11747 16175 11753
rect 16117 11744 16129 11747
rect 15896 11716 16129 11744
rect 15896 11704 15902 11716
rect 16117 11713 16129 11716
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16574 11744 16580 11756
rect 16347 11716 16580 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11744 19579 11747
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 19567 11716 20361 11744
rect 19567 11713 19579 11716
rect 19521 11707 19579 11713
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 21284 11744 21312 11784
rect 22922 11772 22928 11784
rect 22980 11772 22986 11824
rect 24118 11812 24124 11824
rect 23874 11784 24124 11812
rect 24118 11772 24124 11784
rect 24176 11772 24182 11824
rect 20349 11707 20407 11713
rect 20456 11716 21312 11744
rect 13906 11636 13912 11688
rect 13964 11676 13970 11688
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 13964 11648 14105 11676
rect 13964 11636 13970 11648
rect 14093 11645 14105 11648
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 14458 11636 14464 11688
rect 14516 11636 14522 11688
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 16540 11648 16681 11676
rect 16540 11636 16546 11648
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 19610 11676 19616 11688
rect 19484 11648 19616 11676
rect 19484 11636 19490 11648
rect 19610 11636 19616 11648
rect 19668 11676 19674 11688
rect 19705 11679 19763 11685
rect 19705 11676 19717 11679
rect 19668 11648 19717 11676
rect 19668 11636 19674 11648
rect 19705 11645 19717 11648
rect 19751 11676 19763 11679
rect 20456 11676 20484 11716
rect 21358 11704 21364 11756
rect 21416 11704 21422 11756
rect 22370 11704 22376 11756
rect 22428 11704 22434 11756
rect 24228 11753 24256 11852
rect 26142 11840 26148 11852
rect 26200 11840 26206 11892
rect 26789 11883 26847 11889
rect 26789 11849 26801 11883
rect 26835 11880 26847 11883
rect 27522 11880 27528 11892
rect 26835 11852 27528 11880
rect 26835 11849 26847 11852
rect 26789 11843 26847 11849
rect 27522 11840 27528 11852
rect 27580 11840 27586 11892
rect 27614 11840 27620 11892
rect 27672 11880 27678 11892
rect 27672 11852 28212 11880
rect 27672 11840 27678 11852
rect 24486 11772 24492 11824
rect 24544 11772 24550 11824
rect 25774 11812 25780 11824
rect 25714 11784 25780 11812
rect 25774 11772 25780 11784
rect 25832 11812 25838 11824
rect 26326 11812 26332 11824
rect 25832 11784 26332 11812
rect 25832 11772 25838 11784
rect 26326 11772 26332 11784
rect 26384 11812 26390 11824
rect 27433 11815 27491 11821
rect 26384 11784 27292 11812
rect 26384 11772 26390 11784
rect 24213 11747 24271 11753
rect 24213 11713 24225 11747
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 26421 11747 26479 11753
rect 26421 11713 26433 11747
rect 26467 11744 26479 11747
rect 26970 11744 26976 11756
rect 26467 11716 26976 11744
rect 26467 11713 26479 11716
rect 26421 11707 26479 11713
rect 26970 11704 26976 11716
rect 27028 11704 27034 11756
rect 27062 11704 27068 11756
rect 27120 11744 27126 11756
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 27120 11716 27169 11744
rect 27120 11704 27126 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27264 11744 27292 11784
rect 27433 11781 27445 11815
rect 27479 11812 27491 11815
rect 27798 11812 27804 11824
rect 27479 11784 27804 11812
rect 27479 11781 27491 11784
rect 27433 11775 27491 11781
rect 27798 11772 27804 11784
rect 27856 11772 27862 11824
rect 28184 11821 28212 11852
rect 28994 11840 29000 11892
rect 29052 11880 29058 11892
rect 29641 11883 29699 11889
rect 29641 11880 29653 11883
rect 29052 11852 29653 11880
rect 29052 11840 29058 11852
rect 29641 11849 29653 11852
rect 29687 11849 29699 11883
rect 29641 11843 29699 11849
rect 30469 11883 30527 11889
rect 30469 11849 30481 11883
rect 30515 11880 30527 11883
rect 30926 11880 30932 11892
rect 30515 11852 30932 11880
rect 30515 11849 30527 11852
rect 30469 11843 30527 11849
rect 30926 11840 30932 11852
rect 30984 11840 30990 11892
rect 32582 11840 32588 11892
rect 32640 11880 32646 11892
rect 32640 11852 34560 11880
rect 32640 11840 32646 11852
rect 28169 11815 28227 11821
rect 28169 11781 28181 11815
rect 28215 11781 28227 11815
rect 28169 11775 28227 11781
rect 28902 11772 28908 11824
rect 28960 11772 28966 11824
rect 30558 11772 30564 11824
rect 30616 11812 30622 11824
rect 31665 11815 31723 11821
rect 31665 11812 31677 11815
rect 30616 11784 31677 11812
rect 30616 11772 30622 11784
rect 31665 11781 31677 11784
rect 31711 11781 31723 11815
rect 31665 11775 31723 11781
rect 31846 11772 31852 11824
rect 31904 11772 31910 11824
rect 27525 11747 27583 11753
rect 27525 11744 27537 11747
rect 27264 11716 27537 11744
rect 27157 11707 27215 11713
rect 27525 11713 27537 11716
rect 27571 11713 27583 11747
rect 27525 11707 27583 11713
rect 27709 11747 27767 11753
rect 27709 11713 27721 11747
rect 27755 11713 27767 11747
rect 27709 11707 27767 11713
rect 19751 11648 20484 11676
rect 19751 11645 19763 11648
rect 19705 11639 19763 11645
rect 20530 11636 20536 11688
rect 20588 11676 20594 11688
rect 20901 11679 20959 11685
rect 20901 11676 20913 11679
rect 20588 11648 20913 11676
rect 20588 11636 20594 11648
rect 20901 11645 20913 11648
rect 20947 11645 20959 11679
rect 20901 11639 20959 11645
rect 21269 11679 21327 11685
rect 21269 11645 21281 11679
rect 21315 11676 21327 11679
rect 22278 11676 22284 11688
rect 21315 11648 22284 11676
rect 21315 11645 21327 11648
rect 21269 11639 21327 11645
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 22646 11636 22652 11688
rect 22704 11636 22710 11688
rect 26513 11679 26571 11685
rect 24044 11648 26464 11676
rect 12860 11580 13676 11608
rect 18417 11611 18475 11617
rect 12860 11568 12866 11580
rect 18417 11577 18429 11611
rect 18463 11608 18475 11611
rect 20070 11608 20076 11620
rect 18463 11580 20076 11608
rect 18463 11577 18475 11580
rect 18417 11571 18475 11577
rect 20070 11568 20076 11580
rect 20128 11568 20134 11620
rect 11940 11512 12480 11540
rect 12621 11543 12679 11549
rect 11940 11500 11946 11512
rect 12621 11509 12633 11543
rect 12667 11540 12679 11543
rect 13170 11540 13176 11552
rect 12667 11512 13176 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 13780 11512 13829 11540
rect 13780 11500 13786 11512
rect 13817 11509 13829 11512
rect 13863 11509 13875 11543
rect 13817 11503 13875 11509
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11540 14795 11543
rect 15470 11540 15476 11552
rect 14783 11512 15476 11540
rect 14783 11509 14795 11512
rect 14737 11503 14795 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 19978 11500 19984 11552
rect 20036 11540 20042 11552
rect 21085 11543 21143 11549
rect 21085 11540 21097 11543
rect 20036 11512 21097 11540
rect 20036 11500 20042 11512
rect 21085 11509 21097 11512
rect 21131 11509 21143 11543
rect 21085 11503 21143 11509
rect 21545 11543 21603 11549
rect 21545 11509 21557 11543
rect 21591 11540 21603 11543
rect 24044 11540 24072 11648
rect 21591 11512 24072 11540
rect 21591 11509 21603 11512
rect 21545 11503 21603 11509
rect 24118 11500 24124 11552
rect 24176 11500 24182 11552
rect 24854 11500 24860 11552
rect 24912 11540 24918 11552
rect 25222 11540 25228 11552
rect 24912 11512 25228 11540
rect 24912 11500 24918 11512
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 25961 11543 26019 11549
rect 25961 11540 25973 11543
rect 25556 11512 25973 11540
rect 25556 11500 25562 11512
rect 25961 11509 25973 11512
rect 26007 11540 26019 11543
rect 26050 11540 26056 11552
rect 26007 11512 26056 11540
rect 26007 11509 26019 11512
rect 25961 11503 26019 11509
rect 26050 11500 26056 11512
rect 26108 11500 26114 11552
rect 26436 11549 26464 11648
rect 26513 11645 26525 11679
rect 26559 11645 26571 11679
rect 26513 11639 26571 11645
rect 26528 11608 26556 11639
rect 26602 11636 26608 11688
rect 26660 11676 26666 11688
rect 26660 11648 27200 11676
rect 26660 11636 26666 11648
rect 26973 11611 27031 11617
rect 26973 11608 26985 11611
rect 26528 11580 26985 11608
rect 26973 11577 26985 11580
rect 27019 11577 27031 11611
rect 26973 11571 27031 11577
rect 27172 11549 27200 11648
rect 27246 11636 27252 11688
rect 27304 11636 27310 11688
rect 27722 11676 27750 11707
rect 27890 11704 27896 11756
rect 27948 11704 27954 11756
rect 30377 11747 30435 11753
rect 30377 11713 30389 11747
rect 30423 11744 30435 11747
rect 30929 11747 30987 11753
rect 30929 11744 30941 11747
rect 30423 11716 30941 11744
rect 30423 11713 30435 11716
rect 30377 11707 30435 11713
rect 30929 11713 30941 11716
rect 30975 11713 30987 11747
rect 30929 11707 30987 11713
rect 31018 11704 31024 11756
rect 31076 11744 31082 11756
rect 32692 11753 32720 11852
rect 32953 11815 33011 11821
rect 32953 11781 32965 11815
rect 32999 11812 33011 11815
rect 33226 11812 33232 11824
rect 32999 11784 33232 11812
rect 32999 11781 33011 11784
rect 32953 11775 33011 11781
rect 33226 11772 33232 11784
rect 33284 11772 33290 11824
rect 33410 11772 33416 11824
rect 33468 11772 33474 11824
rect 34532 11753 34560 11852
rect 36170 11840 36176 11892
rect 36228 11880 36234 11892
rect 36265 11883 36323 11889
rect 36265 11880 36277 11883
rect 36228 11852 36277 11880
rect 36228 11840 36234 11852
rect 36265 11849 36277 11852
rect 36311 11880 36323 11883
rect 36354 11880 36360 11892
rect 36311 11852 36360 11880
rect 36311 11849 36323 11852
rect 36265 11843 36323 11849
rect 36354 11840 36360 11852
rect 36412 11840 36418 11892
rect 36722 11840 36728 11892
rect 36780 11840 36786 11892
rect 36814 11840 36820 11892
rect 36872 11840 36878 11892
rect 40586 11880 40592 11892
rect 39224 11852 40592 11880
rect 34790 11772 34796 11824
rect 34848 11772 34854 11824
rect 35342 11772 35348 11824
rect 35400 11772 35406 11824
rect 39224 11821 39252 11852
rect 40586 11840 40592 11852
rect 40644 11840 40650 11892
rect 40678 11840 40684 11892
rect 40736 11840 40742 11892
rect 39209 11815 39267 11821
rect 39209 11781 39221 11815
rect 39255 11781 39267 11815
rect 39209 11775 39267 11781
rect 32677 11747 32735 11753
rect 31076 11716 31708 11744
rect 31076 11704 31082 11716
rect 30558 11676 30564 11688
rect 27722 11648 30564 11676
rect 30558 11636 30564 11648
rect 30616 11636 30622 11688
rect 30653 11679 30711 11685
rect 30653 11645 30665 11679
rect 30699 11676 30711 11679
rect 31386 11676 31392 11688
rect 30699 11648 31392 11676
rect 30699 11645 30711 11648
rect 30653 11639 30711 11645
rect 31386 11636 31392 11648
rect 31444 11636 31450 11688
rect 31570 11636 31576 11688
rect 31628 11636 31634 11688
rect 31680 11676 31708 11716
rect 32677 11713 32689 11747
rect 32723 11713 32735 11747
rect 32677 11707 32735 11713
rect 34517 11747 34575 11753
rect 34517 11713 34529 11747
rect 34563 11713 34575 11747
rect 41138 11744 41144 11756
rect 40342 11730 41144 11744
rect 34517 11707 34575 11713
rect 40328 11716 41144 11730
rect 37001 11679 37059 11685
rect 31680 11648 36492 11676
rect 26421 11543 26479 11549
rect 26421 11509 26433 11543
rect 26467 11509 26479 11543
rect 26421 11503 26479 11509
rect 27157 11543 27215 11549
rect 27157 11509 27169 11543
rect 27203 11509 27215 11543
rect 27264 11540 27292 11636
rect 29178 11568 29184 11620
rect 29236 11608 29242 11620
rect 32030 11608 32036 11620
rect 29236 11580 32036 11608
rect 29236 11568 29242 11580
rect 32030 11568 32036 11580
rect 32088 11608 32094 11620
rect 32490 11608 32496 11620
rect 32088 11580 32496 11608
rect 32088 11568 32094 11580
rect 32490 11568 32496 11580
rect 32548 11568 32554 11620
rect 34425 11611 34483 11617
rect 34425 11577 34437 11611
rect 34471 11608 34483 11611
rect 34514 11608 34520 11620
rect 34471 11580 34520 11608
rect 34471 11577 34483 11580
rect 34425 11571 34483 11577
rect 34514 11568 34520 11580
rect 34572 11568 34578 11620
rect 36078 11568 36084 11620
rect 36136 11608 36142 11620
rect 36357 11611 36415 11617
rect 36357 11608 36369 11611
rect 36136 11580 36369 11608
rect 36136 11568 36142 11580
rect 36357 11577 36369 11580
rect 36403 11577 36415 11611
rect 36464 11608 36492 11648
rect 37001 11645 37013 11679
rect 37047 11676 37059 11679
rect 37642 11676 37648 11688
rect 37047 11648 37648 11676
rect 37047 11645 37059 11648
rect 37001 11639 37059 11645
rect 37642 11636 37648 11648
rect 37700 11636 37706 11688
rect 37918 11636 37924 11688
rect 37976 11676 37982 11688
rect 38470 11676 38476 11688
rect 37976 11648 38476 11676
rect 37976 11636 37982 11648
rect 38470 11636 38476 11648
rect 38528 11676 38534 11688
rect 38933 11679 38991 11685
rect 38933 11676 38945 11679
rect 38528 11648 38945 11676
rect 38528 11636 38534 11648
rect 38933 11645 38945 11648
rect 38979 11645 38991 11679
rect 40328 11676 40356 11716
rect 41138 11704 41144 11716
rect 41196 11704 41202 11756
rect 38933 11639 38991 11645
rect 39040 11648 40356 11676
rect 37550 11608 37556 11620
rect 36464 11580 37556 11608
rect 36357 11571 36415 11577
rect 37550 11568 37556 11580
rect 37608 11568 37614 11620
rect 38378 11568 38384 11620
rect 38436 11608 38442 11620
rect 38562 11608 38568 11620
rect 38436 11580 38568 11608
rect 38436 11568 38442 11580
rect 38562 11568 38568 11580
rect 38620 11608 38626 11620
rect 39040 11608 39068 11648
rect 38620 11580 39068 11608
rect 38620 11568 38626 11580
rect 28718 11540 28724 11552
rect 27264 11512 28724 11540
rect 27157 11503 27215 11509
rect 28718 11500 28724 11512
rect 28776 11500 28782 11552
rect 29822 11500 29828 11552
rect 29880 11540 29886 11552
rect 30009 11543 30067 11549
rect 30009 11540 30021 11543
rect 29880 11512 30021 11540
rect 29880 11500 29886 11512
rect 30009 11509 30021 11512
rect 30055 11509 30067 11543
rect 30009 11503 30067 11509
rect 30190 11500 30196 11552
rect 30248 11540 30254 11552
rect 35526 11540 35532 11552
rect 30248 11512 35532 11540
rect 30248 11500 30254 11512
rect 35526 11500 35532 11512
rect 35584 11500 35590 11552
rect 1104 11450 42504 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 42504 11450
rect 1104 11376 42504 11398
rect 3329 11339 3387 11345
rect 3329 11305 3341 11339
rect 3375 11336 3387 11339
rect 4062 11336 4068 11348
rect 3375 11308 4068 11336
rect 3375 11305 3387 11308
rect 3329 11299 3387 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9198 11339 9256 11345
rect 9198 11336 9210 11339
rect 8996 11308 9210 11336
rect 8996 11296 9002 11308
rect 9198 11305 9210 11308
rect 9244 11305 9256 11339
rect 9198 11299 9256 11305
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 11701 11339 11759 11345
rect 11701 11336 11713 11339
rect 9364 11308 11713 11336
rect 9364 11296 9370 11308
rect 11701 11305 11713 11308
rect 11747 11305 11759 11339
rect 11701 11299 11759 11305
rect 12526 11296 12532 11348
rect 12584 11296 12590 11348
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13136 11308 13277 11336
rect 13136 11296 13142 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 13446 11296 13452 11348
rect 13504 11296 13510 11348
rect 13722 11296 13728 11348
rect 13780 11296 13786 11348
rect 13906 11296 13912 11348
rect 13964 11296 13970 11348
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 17586 11345 17592 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14516 11308 14933 11336
rect 14516 11296 14522 11308
rect 14921 11305 14933 11308
rect 14967 11305 14979 11339
rect 14921 11299 14979 11305
rect 17543 11339 17592 11345
rect 17543 11305 17555 11339
rect 17589 11305 17592 11339
rect 17543 11299 17592 11305
rect 17586 11296 17592 11299
rect 17644 11296 17650 11348
rect 19610 11336 19616 11348
rect 19352 11308 19616 11336
rect 3234 11228 3240 11280
rect 3292 11268 3298 11280
rect 3292 11240 3924 11268
rect 3292 11228 3298 11240
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 1581 11203 1639 11209
rect 1581 11200 1593 11203
rect 1544 11172 1593 11200
rect 1544 11160 1550 11172
rect 1581 11169 1593 11172
rect 1627 11200 1639 11203
rect 2866 11200 2872 11212
rect 1627 11172 2872 11200
rect 1627 11169 1639 11172
rect 1581 11163 1639 11169
rect 2866 11160 2872 11172
rect 2924 11200 2930 11212
rect 3510 11200 3516 11212
rect 2924 11172 3516 11200
rect 2924 11160 2930 11172
rect 3510 11160 3516 11172
rect 3568 11200 3574 11212
rect 3789 11203 3847 11209
rect 3789 11200 3801 11203
rect 3568 11172 3801 11200
rect 3568 11160 3574 11172
rect 3789 11169 3801 11172
rect 3835 11169 3847 11203
rect 3896 11200 3924 11240
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 7432 11240 8217 11268
rect 7432 11228 7438 11240
rect 8205 11237 8217 11240
rect 8251 11237 8263 11271
rect 8205 11231 8263 11237
rect 10686 11228 10692 11280
rect 10744 11228 10750 11280
rect 12897 11271 12955 11277
rect 12897 11268 12909 11271
rect 12360 11240 12909 11268
rect 8846 11200 8852 11212
rect 3896 11172 8852 11200
rect 3789 11163 3847 11169
rect 3418 11092 3424 11144
rect 3476 11092 3482 11144
rect 3602 11092 3608 11144
rect 3660 11092 3666 11144
rect 5184 11118 5212 11172
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11200 8999 11203
rect 11514 11200 11520 11212
rect 8987 11172 11520 11200
rect 8987 11169 8999 11172
rect 8941 11163 8999 11169
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 12360 11209 12388 11240
rect 12897 11237 12909 11240
rect 12943 11237 12955 11271
rect 12897 11231 12955 11237
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 12345 11203 12403 11209
rect 11655 11172 12112 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 6730 11092 6736 11144
rect 6788 11092 6794 11144
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 1857 11067 1915 11073
rect 1857 11033 1869 11067
rect 1903 11064 1915 11067
rect 3234 11064 3240 11076
rect 1903 11036 2268 11064
rect 3082 11036 3240 11064
rect 1903 11033 1915 11036
rect 1857 11027 1915 11033
rect 2240 10996 2268 11036
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 3513 11067 3571 11073
rect 3513 11033 3525 11067
rect 3559 11064 3571 11067
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 3559 11036 4077 11064
rect 3559 11033 3571 11036
rect 3513 11027 3571 11033
rect 4065 11033 4077 11036
rect 4111 11033 4123 11067
rect 4065 11027 4123 11033
rect 2774 10996 2780 11008
rect 2240 10968 2780 10996
rect 2774 10956 2780 10968
rect 2832 10956 2838 11008
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 4890 10996 4896 11008
rect 4304 10968 4896 10996
rect 4304 10956 4310 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5442 10956 5448 11008
rect 5500 10996 5506 11008
rect 5537 10999 5595 11005
rect 5537 10996 5549 10999
rect 5500 10968 5549 10996
rect 5500 10956 5506 10968
rect 5537 10965 5549 10968
rect 5583 10965 5595 10999
rect 5537 10959 5595 10965
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 6549 10999 6607 11005
rect 6549 10996 6561 10999
rect 5960 10968 6561 10996
rect 5960 10956 5966 10968
rect 6549 10965 6561 10968
rect 6595 10965 6607 10999
rect 8404 10996 8432 11095
rect 8478 11092 8484 11144
rect 8536 11092 8542 11144
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 8588 11064 8616 11095
rect 8662 11092 8668 11144
rect 8720 11092 8726 11144
rect 10318 11092 10324 11144
rect 10376 11092 10382 11144
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 11977 11135 12035 11141
rect 11977 11132 11989 11135
rect 11756 11104 11989 11132
rect 11756 11092 11762 11104
rect 11977 11101 11989 11104
rect 12023 11101 12035 11135
rect 12084 11132 12112 11172
rect 12345 11169 12357 11203
rect 12391 11169 12403 11203
rect 12986 11200 12992 11212
rect 12345 11163 12403 11169
rect 12636 11172 12992 11200
rect 12526 11132 12532 11144
rect 12084 11104 12532 11132
rect 11977 11095 12035 11101
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 12636 11141 12664 11172
rect 12986 11160 12992 11172
rect 13044 11160 13050 11212
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 12719 11135 12777 11141
rect 12719 11101 12731 11135
rect 12765 11101 12777 11135
rect 12719 11095 12777 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11132 12955 11135
rect 13464 11132 13492 11296
rect 18966 11268 18972 11280
rect 18800 11240 18972 11268
rect 13630 11160 13636 11212
rect 13688 11160 13694 11212
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14277 11203 14335 11209
rect 14277 11200 14289 11203
rect 14056 11172 14289 11200
rect 14056 11160 14062 11172
rect 14277 11169 14289 11172
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 15746 11160 15752 11212
rect 15804 11200 15810 11212
rect 16482 11200 16488 11212
rect 15804 11172 16488 11200
rect 15804 11160 15810 11172
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 18800 11209 18828 11240
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11169 18843 11203
rect 18785 11163 18843 11169
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 19352 11200 19380 11308
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 22557 11339 22615 11345
rect 22557 11305 22569 11339
rect 22603 11336 22615 11339
rect 22646 11336 22652 11348
rect 22603 11308 22652 11336
rect 22603 11305 22615 11308
rect 22557 11299 22615 11305
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 29178 11336 29184 11348
rect 22756 11308 29184 11336
rect 22462 11228 22468 11280
rect 22520 11268 22526 11280
rect 22756 11268 22784 11308
rect 29178 11296 29184 11308
rect 29236 11296 29242 11348
rect 30374 11296 30380 11348
rect 30432 11336 30438 11348
rect 30432 11308 31340 11336
rect 30432 11296 30438 11308
rect 24854 11268 24860 11280
rect 22520 11240 22784 11268
rect 23124 11240 24860 11268
rect 22520 11228 22526 11240
rect 18923 11172 19380 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 19518 11160 19524 11212
rect 19576 11160 19582 11212
rect 19886 11160 19892 11212
rect 19944 11200 19950 11212
rect 20530 11200 20536 11212
rect 19944 11172 20536 11200
rect 19944 11160 19950 11172
rect 20530 11160 20536 11172
rect 20588 11200 20594 11212
rect 20993 11203 21051 11209
rect 20993 11200 21005 11203
rect 20588 11172 21005 11200
rect 20588 11160 20594 11172
rect 20993 11169 21005 11172
rect 21039 11169 21051 11203
rect 23124 11200 23152 11240
rect 24854 11228 24860 11240
rect 24912 11228 24918 11280
rect 26510 11228 26516 11280
rect 26568 11268 26574 11280
rect 29270 11268 29276 11280
rect 26568 11240 29276 11268
rect 26568 11228 26574 11240
rect 29270 11228 29276 11240
rect 29328 11228 29334 11280
rect 31312 11277 31340 11308
rect 31386 11296 31392 11348
rect 31444 11336 31450 11348
rect 31481 11339 31539 11345
rect 31481 11336 31493 11339
rect 31444 11308 31493 11336
rect 31444 11296 31450 11308
rect 31481 11305 31493 11308
rect 31527 11336 31539 11339
rect 32766 11336 32772 11348
rect 31527 11308 32772 11336
rect 31527 11305 31539 11308
rect 31481 11299 31539 11305
rect 32766 11296 32772 11308
rect 32824 11296 32830 11348
rect 34146 11296 34152 11348
rect 34204 11336 34210 11348
rect 34606 11336 34612 11348
rect 34204 11308 34612 11336
rect 34204 11296 34210 11308
rect 34606 11296 34612 11308
rect 34664 11296 34670 11348
rect 35526 11296 35532 11348
rect 35584 11296 35590 11348
rect 37182 11296 37188 11348
rect 37240 11336 37246 11348
rect 37553 11339 37611 11345
rect 37553 11336 37565 11339
rect 37240 11308 37565 11336
rect 37240 11296 37246 11308
rect 37553 11305 37565 11308
rect 37599 11305 37611 11339
rect 37553 11299 37611 11305
rect 31297 11271 31355 11277
rect 31297 11237 31309 11271
rect 31343 11268 31355 11271
rect 31570 11268 31576 11280
rect 31343 11240 31576 11268
rect 31343 11237 31355 11240
rect 31297 11231 31355 11237
rect 31570 11228 31576 11240
rect 31628 11228 31634 11280
rect 33042 11228 33048 11280
rect 33100 11268 33106 11280
rect 35342 11268 35348 11280
rect 33100 11240 35348 11268
rect 33100 11228 33106 11240
rect 35342 11228 35348 11240
rect 35400 11228 35406 11280
rect 35434 11228 35440 11280
rect 35492 11268 35498 11280
rect 35492 11240 35848 11268
rect 35492 11228 35498 11240
rect 20993 11163 21051 11169
rect 22112 11172 23152 11200
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 12943 11104 13553 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 9306 11064 9312 11076
rect 8588 11036 9312 11064
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 11808 11036 12480 11064
rect 9030 10996 9036 11008
rect 8404 10968 9036 10996
rect 6549 10959 6607 10965
rect 9030 10956 9036 10968
rect 9088 10956 9094 11008
rect 11808 11005 11836 11036
rect 11793 10999 11851 11005
rect 11793 10965 11805 10999
rect 11839 10965 11851 10999
rect 11793 10959 11851 10965
rect 11882 10956 11888 11008
rect 11940 10956 11946 11008
rect 12066 10956 12072 11008
rect 12124 10956 12130 11008
rect 12452 10996 12480 11036
rect 12728 10996 12756 11095
rect 16114 11092 16120 11144
rect 16172 11092 16178 11144
rect 18322 11092 18328 11144
rect 18380 11132 18386 11144
rect 22112 11141 22140 11172
rect 23198 11160 23204 11212
rect 23256 11160 23262 11212
rect 24118 11160 24124 11212
rect 24176 11160 24182 11212
rect 24949 11203 25007 11209
rect 24949 11169 24961 11203
rect 24995 11200 25007 11203
rect 26418 11200 26424 11212
rect 24995 11172 26424 11200
rect 24995 11169 25007 11172
rect 24949 11163 25007 11169
rect 26418 11160 26424 11172
rect 26476 11160 26482 11212
rect 26602 11160 26608 11212
rect 26660 11200 26666 11212
rect 26697 11203 26755 11209
rect 26697 11200 26709 11203
rect 26660 11172 26709 11200
rect 26660 11160 26666 11172
rect 26697 11169 26709 11172
rect 26743 11200 26755 11203
rect 27341 11203 27399 11209
rect 27341 11200 27353 11203
rect 26743 11172 27353 11200
rect 26743 11169 26755 11172
rect 26697 11163 26755 11169
rect 27341 11169 27353 11172
rect 27387 11169 27399 11203
rect 27341 11163 27399 11169
rect 29549 11203 29607 11209
rect 29549 11169 29561 11203
rect 29595 11200 29607 11203
rect 31662 11200 31668 11212
rect 29595 11172 31668 11200
rect 29595 11169 29607 11172
rect 29549 11163 29607 11169
rect 31662 11160 31668 11172
rect 31720 11160 31726 11212
rect 33502 11160 33508 11212
rect 33560 11160 33566 11212
rect 35250 11160 35256 11212
rect 35308 11200 35314 11212
rect 35820 11209 35848 11240
rect 35621 11203 35679 11209
rect 35621 11200 35633 11203
rect 35308 11172 35633 11200
rect 35308 11160 35314 11172
rect 35621 11169 35633 11172
rect 35667 11169 35679 11203
rect 35621 11163 35679 11169
rect 35805 11203 35863 11209
rect 35805 11169 35817 11203
rect 35851 11169 35863 11203
rect 35805 11163 35863 11169
rect 36078 11160 36084 11212
rect 36136 11160 36142 11212
rect 38378 11200 38384 11212
rect 37200 11172 38384 11200
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18380 11104 19257 11132
rect 18380 11092 18386 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 22005 11135 22063 11141
rect 22005 11101 22017 11135
rect 22051 11101 22063 11135
rect 22005 11095 22063 11101
rect 22097 11135 22155 11141
rect 22097 11101 22109 11135
rect 22143 11101 22155 11135
rect 22097 11095 22155 11101
rect 12802 11024 12808 11076
rect 12860 11064 12866 11076
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 12860 11036 13093 11064
rect 12860 11024 12866 11036
rect 13081 11033 13093 11036
rect 13127 11033 13139 11067
rect 13081 11027 13139 11033
rect 14550 11024 14556 11076
rect 14608 11064 14614 11076
rect 15102 11064 15108 11076
rect 14608 11036 15108 11064
rect 14608 11024 14614 11036
rect 15102 11024 15108 11036
rect 15160 11064 15166 11076
rect 18693 11067 18751 11073
rect 15160 11036 15884 11064
rect 15160 11024 15166 11036
rect 13170 10996 13176 11008
rect 12452 10968 13176 10996
rect 13170 10956 13176 10968
rect 13228 10956 13234 11008
rect 13262 10956 13268 11008
rect 13320 11005 13326 11008
rect 13320 10999 13339 11005
rect 13327 10965 13339 10999
rect 15856 10996 15884 11036
rect 16408 11036 16514 11064
rect 16408 10996 16436 11036
rect 18693 11033 18705 11067
rect 18739 11064 18751 11067
rect 19426 11064 19432 11076
rect 18739 11036 19432 11064
rect 18739 11033 18751 11036
rect 18693 11027 18751 11033
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 20162 11024 20168 11076
rect 20220 11024 20226 11076
rect 22020 11064 22048 11095
rect 22370 11092 22376 11144
rect 22428 11092 22434 11144
rect 23017 11135 23075 11141
rect 23017 11101 23029 11135
rect 23063 11132 23075 11135
rect 23290 11132 23296 11144
rect 23063 11104 23296 11132
rect 23063 11101 23075 11104
rect 23017 11095 23075 11101
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 26326 11092 26332 11144
rect 26384 11092 26390 11144
rect 27982 11092 27988 11144
rect 28040 11132 28046 11144
rect 28261 11135 28319 11141
rect 28261 11132 28273 11135
rect 28040 11104 28273 11132
rect 28040 11092 28046 11104
rect 28261 11101 28273 11104
rect 28307 11101 28319 11135
rect 31846 11132 31852 11144
rect 28261 11095 28319 11101
rect 31128 11104 31852 11132
rect 22189 11067 22247 11073
rect 22020 11036 22094 11064
rect 15856 10968 16436 10996
rect 18325 10999 18383 11005
rect 13320 10959 13339 10965
rect 18325 10965 18337 10999
rect 18371 10996 18383 10999
rect 18598 10996 18604 11008
rect 18371 10968 18604 10996
rect 18371 10965 18383 10968
rect 18325 10959 18383 10965
rect 13320 10956 13326 10959
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 21082 10956 21088 11008
rect 21140 10996 21146 11008
rect 21821 10999 21879 11005
rect 21821 10996 21833 10999
rect 21140 10968 21833 10996
rect 21140 10956 21146 10968
rect 21821 10965 21833 10968
rect 21867 10965 21879 10999
rect 22066 10996 22094 11036
rect 22189 11033 22201 11067
rect 22235 11064 22247 11067
rect 22830 11064 22836 11076
rect 22235 11036 22836 11064
rect 22235 11033 22247 11036
rect 22189 11027 22247 11033
rect 22830 11024 22836 11036
rect 22888 11024 22894 11076
rect 22925 11067 22983 11073
rect 22925 11033 22937 11067
rect 22971 11064 22983 11067
rect 23569 11067 23627 11073
rect 23569 11064 23581 11067
rect 22971 11036 23581 11064
rect 22971 11033 22983 11036
rect 22925 11027 22983 11033
rect 23569 11033 23581 11036
rect 23615 11033 23627 11067
rect 23569 11027 23627 11033
rect 25222 11024 25228 11076
rect 25280 11024 25286 11076
rect 29822 11024 29828 11076
rect 29880 11024 29886 11076
rect 30466 11024 30472 11076
rect 30524 11024 30530 11076
rect 23290 10996 23296 11008
rect 22066 10968 23296 10996
rect 21821 10959 21879 10965
rect 23290 10956 23296 10968
rect 23348 10956 23354 11008
rect 26786 10956 26792 11008
rect 26844 10956 26850 11008
rect 27706 10956 27712 11008
rect 27764 10956 27770 11008
rect 30558 10956 30564 11008
rect 30616 10996 30622 11008
rect 31128 10996 31156 11104
rect 31846 11092 31852 11104
rect 31904 11092 31910 11144
rect 32490 11092 32496 11144
rect 32548 11092 32554 11144
rect 31757 11067 31815 11073
rect 31757 11033 31769 11067
rect 31803 11064 31815 11067
rect 32030 11064 32036 11076
rect 31803 11036 32036 11064
rect 31803 11033 31815 11036
rect 31757 11027 31815 11033
rect 32030 11024 32036 11036
rect 32088 11024 32094 11076
rect 32766 11024 32772 11076
rect 32824 11064 32830 11076
rect 33520 11064 33548 11160
rect 34514 11092 34520 11144
rect 34572 11132 34578 11144
rect 34793 11135 34851 11141
rect 34793 11132 34805 11135
rect 34572 11104 34805 11132
rect 34572 11092 34578 11104
rect 34793 11101 34805 11104
rect 34839 11101 34851 11135
rect 34793 11095 34851 11101
rect 34885 11135 34943 11141
rect 34885 11101 34897 11135
rect 34931 11132 34943 11135
rect 35342 11132 35348 11144
rect 34931 11104 35348 11132
rect 34931 11101 34943 11104
rect 34885 11095 34943 11101
rect 35342 11092 35348 11104
rect 35400 11092 35406 11144
rect 35434 11092 35440 11144
rect 35492 11092 35498 11144
rect 37200 11118 37228 11172
rect 38378 11160 38384 11172
rect 38436 11160 38442 11212
rect 37645 11135 37703 11141
rect 37645 11101 37657 11135
rect 37691 11101 37703 11135
rect 37645 11095 37703 11101
rect 33870 11064 33876 11076
rect 32824 11036 33876 11064
rect 32824 11024 32830 11036
rect 33870 11024 33876 11036
rect 33928 11064 33934 11076
rect 35158 11064 35164 11076
rect 33928 11036 35164 11064
rect 33928 11024 33934 11036
rect 35158 11024 35164 11036
rect 35216 11064 35222 11076
rect 37660 11064 37688 11095
rect 37826 11092 37832 11144
rect 37884 11092 37890 11144
rect 38013 11135 38071 11141
rect 38013 11101 38025 11135
rect 38059 11101 38071 11135
rect 38013 11095 38071 11101
rect 35216 11036 36492 11064
rect 35216 11024 35222 11036
rect 30616 10968 31156 10996
rect 30616 10956 30622 10968
rect 31938 10956 31944 11008
rect 31996 10956 32002 11008
rect 32306 10956 32312 11008
rect 32364 10996 32370 11008
rect 36354 10996 36360 11008
rect 32364 10968 36360 10996
rect 32364 10956 32370 10968
rect 36354 10956 36360 10968
rect 36412 10956 36418 11008
rect 36464 10996 36492 11036
rect 37384 11036 37688 11064
rect 37737 11067 37795 11073
rect 37384 10996 37412 11036
rect 37737 11033 37749 11067
rect 37783 11064 37795 11067
rect 38028 11064 38056 11095
rect 37783 11036 38056 11064
rect 37783 11033 37795 11036
rect 37737 11027 37795 11033
rect 36464 10968 37412 10996
rect 37826 10956 37832 11008
rect 37884 10996 37890 11008
rect 38197 10999 38255 11005
rect 38197 10996 38209 10999
rect 37884 10968 38209 10996
rect 37884 10956 37890 10968
rect 38197 10965 38209 10968
rect 38243 10996 38255 10999
rect 38286 10996 38292 11008
rect 38243 10968 38292 10996
rect 38243 10965 38255 10968
rect 38197 10959 38255 10965
rect 38286 10956 38292 10968
rect 38344 10956 38350 11008
rect 1104 10906 42504 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 42504 10906
rect 1104 10832 42504 10854
rect 1210 10752 1216 10804
rect 1268 10792 1274 10804
rect 1489 10795 1547 10801
rect 1489 10792 1501 10795
rect 1268 10764 1501 10792
rect 1268 10752 1274 10764
rect 1489 10761 1501 10764
rect 1535 10761 1547 10795
rect 1489 10755 1547 10761
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 1820 10764 2513 10792
rect 1820 10752 1826 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 2501 10755 2559 10761
rect 3602 10752 3608 10804
rect 3660 10792 3666 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 3660 10764 4537 10792
rect 3660 10752 3666 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 4693 10795 4751 10801
rect 4693 10761 4705 10795
rect 4739 10792 4751 10795
rect 4798 10792 4804 10804
rect 4739 10764 4804 10792
rect 4739 10761 4751 10764
rect 4693 10755 4751 10761
rect 4798 10752 4804 10764
rect 4856 10792 4862 10804
rect 4856 10764 6408 10792
rect 4856 10752 4862 10764
rect 3694 10724 3700 10736
rect 2608 10696 3700 10724
rect 2608 10665 2636 10696
rect 3694 10684 3700 10696
rect 3752 10684 3758 10736
rect 4893 10727 4951 10733
rect 4893 10693 4905 10727
rect 4939 10693 4951 10727
rect 4893 10687 4951 10693
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 2409 10659 2467 10665
rect 2409 10625 2421 10659
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10625 2651 10659
rect 2593 10619 2651 10625
rect 1688 10520 1716 10619
rect 2424 10588 2452 10619
rect 2682 10616 2688 10668
rect 2740 10656 2746 10668
rect 2777 10659 2835 10665
rect 2777 10656 2789 10659
rect 2740 10628 2789 10656
rect 2740 10616 2746 10628
rect 2777 10625 2789 10628
rect 2823 10625 2835 10659
rect 2777 10619 2835 10625
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 3099 10628 3249 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 3970 10656 3976 10668
rect 3237 10619 3295 10625
rect 3804 10628 3976 10656
rect 2700 10588 2728 10616
rect 2424 10560 2728 10588
rect 2884 10588 2912 10619
rect 3804 10588 3832 10628
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4522 10656 4528 10668
rect 4295 10628 4528 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 2884 10560 3832 10588
rect 3881 10591 3939 10597
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 4172 10588 4200 10616
rect 4798 10588 4804 10600
rect 3927 10560 4200 10588
rect 4356 10560 4804 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 4246 10520 4252 10532
rect 1688 10492 4252 10520
rect 4246 10480 4252 10492
rect 4304 10480 4310 10532
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 3142 10452 3148 10464
rect 3099 10424 3148 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 4356 10452 4384 10560
rect 4798 10548 4804 10560
rect 4856 10588 4862 10600
rect 4908 10588 4936 10687
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5684 10628 5733 10656
rect 5684 10616 5690 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6380 10665 6408 10764
rect 8294 10752 8300 10804
rect 8352 10752 8358 10804
rect 8386 10752 8392 10804
rect 8444 10792 8450 10804
rect 8481 10795 8539 10801
rect 8481 10792 8493 10795
rect 8444 10764 8493 10792
rect 8444 10752 8450 10764
rect 8481 10761 8493 10764
rect 8527 10761 8539 10795
rect 8481 10755 8539 10761
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 9125 10795 9183 10801
rect 9125 10792 9137 10795
rect 8720 10764 9137 10792
rect 8720 10752 8726 10764
rect 9125 10761 9137 10764
rect 9171 10761 9183 10795
rect 9125 10755 9183 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13722 10792 13728 10804
rect 12860 10764 13728 10792
rect 12860 10752 12866 10764
rect 7098 10724 7104 10736
rect 6472 10696 7104 10724
rect 6365 10659 6423 10665
rect 5868 10628 6316 10656
rect 5868 10616 5874 10628
rect 5442 10588 5448 10600
rect 4856 10560 5448 10588
rect 4856 10548 4862 10560
rect 5442 10548 5448 10560
rect 5500 10588 5506 10600
rect 5905 10591 5963 10597
rect 5905 10588 5917 10591
rect 5500 10560 5917 10588
rect 5500 10548 5506 10560
rect 5905 10557 5917 10560
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 5994 10548 6000 10600
rect 6052 10548 6058 10600
rect 6288 10588 6316 10628
rect 6365 10625 6377 10659
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6472 10588 6500 10696
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 7300 10696 7972 10724
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 7300 10656 7328 10696
rect 6549 10619 6607 10625
rect 7024 10628 7328 10656
rect 6288 10560 6500 10588
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 6564 10520 6592 10619
rect 5592 10492 6592 10520
rect 5592 10480 5598 10492
rect 4203 10424 4384 10452
rect 4433 10455 4491 10461
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4614 10452 4620 10464
rect 4479 10424 4620 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4706 10412 4712 10464
rect 4764 10412 4770 10464
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 5316 10424 6469 10452
rect 5316 10412 5322 10424
rect 6457 10421 6469 10424
rect 6503 10452 6515 10455
rect 7024 10452 7052 10628
rect 7374 10616 7380 10668
rect 7432 10616 7438 10668
rect 7944 10665 7972 10696
rect 8128 10696 9076 10724
rect 8128 10665 8156 10696
rect 9048 10668 9076 10696
rect 10318 10684 10324 10736
rect 10376 10724 10382 10736
rect 10376 10696 12282 10724
rect 10376 10684 10382 10696
rect 13078 10684 13084 10736
rect 13136 10724 13142 10736
rect 13648 10733 13676 10764
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 13998 10752 14004 10804
rect 14056 10752 14062 10804
rect 19426 10752 19432 10804
rect 19484 10792 19490 10804
rect 20165 10795 20223 10801
rect 20165 10792 20177 10795
rect 19484 10764 20177 10792
rect 19484 10752 19490 10764
rect 20165 10761 20177 10764
rect 20211 10761 20223 10795
rect 20165 10755 20223 10761
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 22925 10795 22983 10801
rect 22925 10792 22937 10795
rect 22428 10764 22937 10792
rect 22428 10752 22434 10764
rect 22925 10761 22937 10764
rect 22971 10761 22983 10795
rect 22925 10755 22983 10761
rect 13541 10727 13599 10733
rect 13541 10724 13553 10727
rect 13136 10696 13553 10724
rect 13136 10684 13142 10696
rect 13541 10693 13553 10696
rect 13587 10693 13599 10727
rect 13541 10687 13599 10693
rect 13633 10727 13691 10733
rect 13633 10693 13645 10727
rect 13679 10693 13691 10727
rect 13633 10687 13691 10693
rect 14458 10684 14464 10736
rect 14516 10684 14522 10736
rect 15470 10684 15476 10736
rect 15528 10684 15534 10736
rect 18598 10684 18604 10736
rect 18656 10684 18662 10736
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8113 10659 8171 10665
rect 7975 10628 8064 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 7156 10560 7481 10588
rect 7156 10548 7162 10560
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10557 7895 10591
rect 8036 10588 8064 10628
rect 8113 10625 8125 10659
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8260 10628 8677 10656
rect 8260 10616 8266 10628
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 9140 10628 9689 10656
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8036 10560 8585 10588
rect 7837 10551 7895 10557
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 7852 10520 7880 10551
rect 7926 10520 7932 10532
rect 7392 10492 7932 10520
rect 7392 10464 7420 10492
rect 7926 10480 7932 10492
rect 7984 10480 7990 10532
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 9140 10520 9168 10628
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 13354 10616 13360 10668
rect 13412 10616 13418 10668
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10588 9459 10591
rect 9766 10588 9772 10600
rect 9447 10560 9772 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 13262 10588 13268 10600
rect 12492 10560 13268 10588
rect 12492 10548 12498 10560
rect 13262 10548 13268 10560
rect 13320 10588 13326 10600
rect 13630 10588 13636 10600
rect 13320 10560 13636 10588
rect 13320 10548 13326 10560
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 11422 10520 11428 10532
rect 8536 10492 9168 10520
rect 9508 10492 11428 10520
rect 8536 10480 8542 10492
rect 7282 10452 7288 10464
rect 6503 10424 7288 10452
rect 6503 10421 6515 10424
rect 6457 10415 6515 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7374 10412 7380 10464
rect 7432 10412 7438 10464
rect 7745 10455 7803 10461
rect 7745 10421 7757 10455
rect 7791 10452 7803 10455
rect 9508 10452 9536 10492
rect 11422 10480 11428 10492
rect 11480 10480 11486 10532
rect 12894 10480 12900 10532
rect 12952 10520 12958 10532
rect 13740 10520 13768 10619
rect 15746 10616 15752 10668
rect 15804 10616 15810 10668
rect 20162 10656 20168 10668
rect 19734 10628 20168 10656
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 22940 10656 22968 10755
rect 25222 10752 25228 10804
rect 25280 10792 25286 10804
rect 25501 10795 25559 10801
rect 25501 10792 25513 10795
rect 25280 10764 25513 10792
rect 25280 10752 25286 10764
rect 25501 10761 25513 10764
rect 25547 10761 25559 10795
rect 25501 10755 25559 10761
rect 25958 10752 25964 10804
rect 26016 10752 26022 10804
rect 27341 10795 27399 10801
rect 27341 10761 27353 10795
rect 27387 10792 27399 10795
rect 27706 10792 27712 10804
rect 27387 10764 27712 10792
rect 27387 10761 27399 10764
rect 27341 10755 27399 10761
rect 27706 10752 27712 10764
rect 27764 10752 27770 10804
rect 28718 10752 28724 10804
rect 28776 10752 28782 10804
rect 32125 10795 32183 10801
rect 32125 10761 32137 10795
rect 32171 10792 32183 10795
rect 32490 10792 32496 10804
rect 32171 10764 32496 10792
rect 32171 10761 32183 10764
rect 32125 10755 32183 10761
rect 32490 10752 32496 10764
rect 32548 10752 32554 10804
rect 32585 10795 32643 10801
rect 32585 10761 32597 10795
rect 32631 10792 32643 10795
rect 32674 10792 32680 10804
rect 32631 10764 32680 10792
rect 32631 10761 32643 10764
rect 32585 10755 32643 10761
rect 32674 10752 32680 10764
rect 32732 10752 32738 10804
rect 35250 10752 35256 10804
rect 35308 10792 35314 10804
rect 35345 10795 35403 10801
rect 35345 10792 35357 10795
rect 35308 10764 35357 10792
rect 35308 10752 35314 10764
rect 35345 10761 35357 10764
rect 35391 10761 35403 10795
rect 35345 10755 35403 10761
rect 36354 10752 36360 10804
rect 36412 10792 36418 10804
rect 39114 10792 39120 10804
rect 36412 10764 39120 10792
rect 36412 10752 36418 10764
rect 39114 10752 39120 10764
rect 39172 10792 39178 10804
rect 39942 10792 39948 10804
rect 39172 10764 39948 10792
rect 39172 10752 39178 10764
rect 39942 10752 39948 10764
rect 40000 10792 40006 10804
rect 40589 10795 40647 10801
rect 40589 10792 40601 10795
rect 40000 10764 40601 10792
rect 40000 10752 40006 10764
rect 40589 10761 40601 10764
rect 40635 10761 40647 10795
rect 40589 10755 40647 10761
rect 23661 10727 23719 10733
rect 23661 10693 23673 10727
rect 23707 10724 23719 10727
rect 25869 10727 25927 10733
rect 23707 10696 24348 10724
rect 23707 10693 23719 10696
rect 23661 10687 23719 10693
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 22940 10628 23949 10656
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 24029 10659 24087 10665
rect 24029 10625 24041 10659
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10656 24179 10659
rect 24210 10656 24216 10668
rect 24167 10628 24216 10656
rect 24167 10625 24179 10628
rect 24121 10619 24179 10625
rect 18322 10548 18328 10600
rect 18380 10548 18386 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 20088 10560 20729 10588
rect 12952 10492 13768 10520
rect 12952 10480 12958 10492
rect 20088 10464 20116 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22244 10560 22293 10588
rect 22244 10548 22250 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 23014 10548 23020 10600
rect 23072 10548 23078 10600
rect 24044 10588 24072 10619
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 24320 10665 24348 10696
rect 25869 10693 25881 10727
rect 25915 10724 25927 10727
rect 26786 10724 26792 10736
rect 25915 10696 26792 10724
rect 25915 10693 25927 10696
rect 25869 10687 25927 10693
rect 26786 10684 26792 10696
rect 26844 10684 26850 10736
rect 26878 10684 26884 10736
rect 26936 10724 26942 10736
rect 27433 10727 27491 10733
rect 27433 10724 27445 10727
rect 26936 10696 27445 10724
rect 26936 10684 26942 10696
rect 27433 10693 27445 10696
rect 27479 10693 27491 10727
rect 27433 10687 27491 10693
rect 28552 10696 29500 10724
rect 24305 10659 24363 10665
rect 24305 10625 24317 10659
rect 24351 10625 24363 10659
rect 24305 10619 24363 10625
rect 26697 10659 26755 10665
rect 26697 10625 26709 10659
rect 26743 10656 26755 10659
rect 27338 10656 27344 10668
rect 26743 10628 27344 10656
rect 26743 10625 26755 10628
rect 26697 10619 26755 10625
rect 27338 10616 27344 10628
rect 27396 10656 27402 10668
rect 28552 10656 28580 10696
rect 27396 10628 28580 10656
rect 28813 10659 28871 10665
rect 27396 10616 27402 10628
rect 28813 10625 28825 10659
rect 28859 10656 28871 10659
rect 29365 10659 29423 10665
rect 29365 10656 29377 10659
rect 28859 10628 29377 10656
rect 28859 10625 28871 10628
rect 28813 10619 28871 10625
rect 29365 10625 29377 10628
rect 29411 10625 29423 10659
rect 29472 10656 29500 10696
rect 30834 10684 30840 10736
rect 30892 10724 30898 10736
rect 33502 10724 33508 10736
rect 30892 10696 33508 10724
rect 30892 10684 30898 10696
rect 33502 10684 33508 10696
rect 33560 10684 33566 10736
rect 34517 10727 34575 10733
rect 34517 10693 34529 10727
rect 34563 10724 34575 10727
rect 35713 10727 35771 10733
rect 35713 10724 35725 10727
rect 34563 10696 35725 10724
rect 34563 10693 34575 10696
rect 34517 10687 34575 10693
rect 35713 10693 35725 10696
rect 35759 10693 35771 10727
rect 36173 10727 36231 10733
rect 36173 10724 36185 10727
rect 35713 10687 35771 10693
rect 36004 10696 36185 10724
rect 32306 10656 32312 10668
rect 29472 10628 32312 10656
rect 29365 10619 29423 10625
rect 32306 10616 32312 10628
rect 32364 10616 32370 10668
rect 32493 10659 32551 10665
rect 32493 10625 32505 10659
rect 32539 10656 32551 10659
rect 32953 10659 33011 10665
rect 32953 10656 32965 10659
rect 32539 10628 32965 10656
rect 32539 10625 32551 10628
rect 32493 10619 32551 10625
rect 32953 10625 32965 10628
rect 32999 10625 33011 10659
rect 32953 10619 33011 10625
rect 34241 10659 34299 10665
rect 34241 10625 34253 10659
rect 34287 10656 34299 10659
rect 34790 10656 34796 10668
rect 34287 10628 34796 10656
rect 34287 10625 34299 10628
rect 34241 10619 34299 10625
rect 34790 10616 34796 10628
rect 34848 10616 34854 10668
rect 35526 10665 35532 10668
rect 35524 10656 35532 10665
rect 35487 10628 35532 10656
rect 35524 10619 35532 10628
rect 35526 10616 35532 10619
rect 35584 10616 35590 10668
rect 36004 10665 36032 10696
rect 36173 10693 36185 10696
rect 36219 10693 36231 10727
rect 36173 10687 36231 10693
rect 38470 10684 38476 10736
rect 38528 10724 38534 10736
rect 38528 10696 38686 10724
rect 38528 10684 38534 10696
rect 35621 10659 35679 10665
rect 35621 10625 35633 10659
rect 35667 10625 35679 10659
rect 35621 10619 35679 10625
rect 35896 10659 35954 10665
rect 35896 10625 35908 10659
rect 35942 10625 35954 10659
rect 35896 10619 35954 10625
rect 35989 10659 36047 10665
rect 35989 10625 36001 10659
rect 36035 10625 36047 10659
rect 35989 10619 36047 10625
rect 25130 10588 25136 10600
rect 24044 10560 25136 10588
rect 25130 10548 25136 10560
rect 25188 10548 25194 10600
rect 25866 10548 25872 10600
rect 25924 10588 25930 10600
rect 26053 10591 26111 10597
rect 26053 10588 26065 10591
rect 25924 10560 26065 10588
rect 25924 10548 25930 10560
rect 26053 10557 26065 10560
rect 26099 10588 26111 10591
rect 27525 10591 27583 10597
rect 27525 10588 27537 10591
rect 26099 10560 27537 10588
rect 26099 10557 26111 10560
rect 26053 10551 26111 10557
rect 27525 10557 27537 10560
rect 27571 10588 27583 10591
rect 28537 10591 28595 10597
rect 28537 10588 28549 10591
rect 27571 10560 28549 10588
rect 27571 10557 27583 10560
rect 27525 10551 27583 10557
rect 28537 10557 28549 10560
rect 28583 10588 28595 10591
rect 28902 10588 28908 10600
rect 28583 10560 28908 10588
rect 28583 10557 28595 10560
rect 28537 10551 28595 10557
rect 28902 10548 28908 10560
rect 28960 10548 28966 10600
rect 29086 10548 29092 10600
rect 29144 10588 29150 10600
rect 29917 10591 29975 10597
rect 29917 10588 29929 10591
rect 29144 10560 29929 10588
rect 29144 10548 29150 10560
rect 29917 10557 29929 10560
rect 29963 10588 29975 10591
rect 30190 10588 30196 10600
rect 29963 10560 30196 10588
rect 29963 10557 29975 10560
rect 29917 10551 29975 10557
rect 30190 10548 30196 10560
rect 30248 10548 30254 10600
rect 32766 10548 32772 10600
rect 32824 10548 32830 10600
rect 33134 10548 33140 10600
rect 33192 10588 33198 10600
rect 33505 10591 33563 10597
rect 33505 10588 33517 10591
rect 33192 10560 33517 10588
rect 33192 10548 33198 10560
rect 33505 10557 33517 10560
rect 33551 10557 33563 10591
rect 33505 10551 33563 10557
rect 34514 10548 34520 10600
rect 34572 10548 34578 10600
rect 35342 10548 35348 10600
rect 35400 10588 35406 10600
rect 35636 10588 35664 10619
rect 35400 10560 35664 10588
rect 35912 10588 35940 10619
rect 36078 10616 36084 10668
rect 36136 10616 36142 10668
rect 36265 10659 36323 10665
rect 36265 10625 36277 10659
rect 36311 10656 36323 10659
rect 36354 10656 36360 10668
rect 36311 10628 36360 10656
rect 36311 10625 36323 10628
rect 36265 10619 36323 10625
rect 36354 10616 36360 10628
rect 36412 10616 36418 10668
rect 37645 10659 37703 10665
rect 37645 10625 37657 10659
rect 37691 10656 37703 10659
rect 37691 10628 37725 10656
rect 37691 10625 37703 10628
rect 37645 10619 37703 10625
rect 36170 10588 36176 10600
rect 35912 10560 36176 10588
rect 35400 10548 35406 10560
rect 36170 10548 36176 10560
rect 36228 10548 36234 10600
rect 37366 10548 37372 10600
rect 37424 10588 37430 10600
rect 37660 10588 37688 10619
rect 37918 10616 37924 10668
rect 37976 10616 37982 10668
rect 40497 10659 40555 10665
rect 40497 10656 40509 10659
rect 39408 10628 40509 10656
rect 37737 10591 37795 10597
rect 37737 10588 37749 10591
rect 37424 10560 37749 10588
rect 37424 10548 37430 10560
rect 37737 10557 37749 10560
rect 37783 10588 37795 10591
rect 37826 10588 37832 10600
rect 37783 10560 37832 10588
rect 37783 10557 37795 10560
rect 37737 10551 37795 10557
rect 37826 10548 37832 10560
rect 37884 10548 37890 10600
rect 38197 10591 38255 10597
rect 38197 10557 38209 10591
rect 38243 10588 38255 10591
rect 38562 10588 38568 10600
rect 38243 10560 38568 10588
rect 38243 10557 38255 10560
rect 38197 10551 38255 10557
rect 38562 10548 38568 10560
rect 38620 10548 38626 10600
rect 38930 10548 38936 10600
rect 38988 10588 38994 10600
rect 39408 10588 39436 10628
rect 40497 10625 40509 10628
rect 40543 10625 40555 10659
rect 40497 10619 40555 10625
rect 40770 10616 40776 10668
rect 40828 10616 40834 10668
rect 38988 10560 39436 10588
rect 39669 10591 39727 10597
rect 38988 10548 38994 10560
rect 39669 10557 39681 10591
rect 39715 10588 39727 10591
rect 40313 10591 40371 10597
rect 40313 10588 40325 10591
rect 39715 10560 40325 10588
rect 39715 10557 39727 10560
rect 39669 10551 39727 10557
rect 40313 10557 40325 10560
rect 40359 10557 40371 10591
rect 40313 10551 40371 10557
rect 21266 10480 21272 10532
rect 21324 10520 21330 10532
rect 26694 10520 26700 10532
rect 21324 10492 26700 10520
rect 21324 10480 21330 10492
rect 26694 10480 26700 10492
rect 26752 10520 26758 10532
rect 26752 10492 35480 10520
rect 26752 10480 26758 10492
rect 7791 10424 9536 10452
rect 9585 10455 9643 10461
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 10042 10452 10048 10464
rect 9631 10424 10048 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 13262 10412 13268 10464
rect 13320 10412 13326 10464
rect 13906 10412 13912 10464
rect 13964 10412 13970 10464
rect 20070 10412 20076 10464
rect 20128 10412 20134 10464
rect 23750 10412 23756 10464
rect 23808 10412 23814 10464
rect 26326 10412 26332 10464
rect 26384 10452 26390 10464
rect 26421 10455 26479 10461
rect 26421 10452 26433 10455
rect 26384 10424 26433 10452
rect 26384 10412 26390 10424
rect 26421 10421 26433 10424
rect 26467 10421 26479 10455
rect 26421 10415 26479 10421
rect 26510 10412 26516 10464
rect 26568 10452 26574 10464
rect 26973 10455 27031 10461
rect 26973 10452 26985 10455
rect 26568 10424 26985 10452
rect 26568 10412 26574 10424
rect 26973 10421 26985 10424
rect 27019 10421 27031 10455
rect 26973 10415 27031 10421
rect 29181 10455 29239 10461
rect 29181 10421 29193 10455
rect 29227 10452 29239 10455
rect 30098 10452 30104 10464
rect 29227 10424 30104 10452
rect 29227 10421 29239 10424
rect 29181 10415 29239 10421
rect 30098 10412 30104 10424
rect 30156 10412 30162 10464
rect 34330 10412 34336 10464
rect 34388 10412 34394 10464
rect 35452 10452 35480 10492
rect 35526 10480 35532 10532
rect 35584 10520 35590 10532
rect 37642 10520 37648 10532
rect 35584 10492 37648 10520
rect 35584 10480 35590 10492
rect 37642 10480 37648 10492
rect 37700 10480 37706 10532
rect 37366 10452 37372 10464
rect 35452 10424 37372 10452
rect 37366 10412 37372 10424
rect 37424 10412 37430 10464
rect 37458 10412 37464 10464
rect 37516 10412 37522 10464
rect 38838 10412 38844 10464
rect 38896 10452 38902 10464
rect 39761 10455 39819 10461
rect 39761 10452 39773 10455
rect 38896 10424 39773 10452
rect 38896 10412 38902 10424
rect 39761 10421 39773 10424
rect 39807 10421 39819 10455
rect 39761 10415 39819 10421
rect 1104 10362 42504 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 42504 10362
rect 1104 10288 42504 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 3329 10251 3387 10257
rect 3329 10248 3341 10251
rect 2832 10220 3341 10248
rect 2832 10208 2838 10220
rect 3329 10217 3341 10220
rect 3375 10217 3387 10251
rect 3329 10211 3387 10217
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10248 5595 10251
rect 5994 10248 6000 10260
rect 5583 10220 6000 10248
rect 5583 10217 5595 10220
rect 5537 10211 5595 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7374 10248 7380 10260
rect 7055 10220 7380 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11790 10248 11796 10260
rect 11655 10220 11796 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 13354 10208 13360 10260
rect 13412 10208 13418 10260
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13780 10220 14105 10248
rect 13780 10208 13786 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 22186 10208 22192 10260
rect 22244 10208 22250 10260
rect 23290 10208 23296 10260
rect 23348 10208 23354 10260
rect 25685 10251 25743 10257
rect 23860 10220 25084 10248
rect 6546 10180 6552 10192
rect 5552 10152 6552 10180
rect 3142 10004 3148 10056
rect 3200 10004 3206 10056
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10044 3387 10047
rect 3418 10044 3424 10056
rect 3375 10016 3424 10044
rect 3375 10013 3387 10016
rect 3329 10007 3387 10013
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 4672 10016 5365 10044
rect 4672 10004 4678 10016
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 5368 9976 5396 10007
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 5552 10053 5580 10152
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 5644 10084 6316 10112
rect 5644 10053 5672 10084
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5500 10016 5549 10044
rect 5500 10004 5506 10016
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 5644 9976 5672 10007
rect 5810 10004 5816 10056
rect 5868 10004 5874 10056
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5960 10016 6009 10044
rect 5960 10004 5966 10016
rect 5997 10013 6009 10016
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6086 10004 6092 10056
rect 6144 10004 6150 10056
rect 6288 10053 6316 10084
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 11793 10115 11851 10121
rect 11793 10112 11805 10115
rect 11756 10084 11805 10112
rect 11756 10072 11762 10084
rect 11793 10081 11805 10084
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 12066 10072 12072 10124
rect 12124 10112 12130 10124
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 12124 10084 12265 10112
rect 12124 10072 12130 10084
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12253 10075 12311 10081
rect 13262 10072 13268 10124
rect 13320 10072 13326 10124
rect 13630 10072 13636 10124
rect 13688 10072 13694 10124
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 15565 10115 15623 10121
rect 15565 10112 15577 10115
rect 13964 10084 15577 10112
rect 13964 10072 13970 10084
rect 15565 10081 15577 10084
rect 15611 10081 15623 10115
rect 15565 10075 15623 10081
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10112 20775 10115
rect 21082 10112 21088 10124
rect 20763 10084 21088 10112
rect 20763 10081 20775 10084
rect 20717 10075 20775 10081
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 21358 10072 21364 10124
rect 21416 10112 21422 10124
rect 22741 10115 22799 10121
rect 22741 10112 22753 10115
rect 21416 10084 22753 10112
rect 21416 10072 21422 10084
rect 22741 10081 22753 10084
rect 22787 10081 22799 10115
rect 22741 10075 22799 10081
rect 23032 10084 23796 10112
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 5368 9948 5672 9976
rect 5718 9936 5724 9988
rect 5776 9936 5782 9988
rect 6196 9976 6224 10007
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 6730 10004 6736 10056
rect 6788 10044 6794 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6788 10016 6837 10044
rect 6788 10004 6794 10016
rect 6825 10013 6837 10016
rect 6871 10044 6883 10047
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 6871 10016 7113 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 7282 10004 7288 10056
rect 7340 10004 7346 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 12621 10047 12679 10053
rect 12621 10044 12633 10047
rect 11931 10016 12633 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 12621 10013 12633 10016
rect 12667 10013 12679 10047
rect 12621 10007 12679 10013
rect 13722 10004 13728 10056
rect 13780 10004 13786 10056
rect 15838 10004 15844 10056
rect 15896 10004 15902 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 20441 10047 20499 10053
rect 20441 10044 20453 10047
rect 18380 10016 20453 10044
rect 18380 10004 18386 10016
rect 20441 10013 20453 10016
rect 20487 10013 20499 10047
rect 20441 10007 20499 10013
rect 22278 10004 22284 10056
rect 22336 10044 22342 10056
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 22336 10016 22477 10044
rect 22336 10004 22342 10016
rect 22465 10013 22477 10016
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 22646 10004 22652 10056
rect 22704 10004 22710 10056
rect 22830 10004 22836 10056
rect 22888 10004 22894 10056
rect 23032 10053 23060 10084
rect 23017 10047 23075 10053
rect 23017 10013 23029 10047
rect 23063 10013 23075 10047
rect 23017 10007 23075 10013
rect 23290 10004 23296 10056
rect 23348 10004 23354 10056
rect 23382 10004 23388 10056
rect 23440 10044 23446 10056
rect 23477 10047 23535 10053
rect 23477 10044 23489 10047
rect 23440 10016 23489 10044
rect 23440 10004 23446 10016
rect 23477 10013 23489 10016
rect 23523 10013 23535 10047
rect 23477 10007 23535 10013
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 6104 9948 6224 9976
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 6104 9908 6132 9948
rect 14550 9936 14556 9988
rect 14608 9936 14614 9988
rect 20162 9936 20168 9988
rect 20220 9976 20226 9988
rect 21174 9976 21180 9988
rect 20220 9948 21180 9976
rect 20220 9936 20226 9948
rect 21174 9936 21180 9948
rect 21232 9936 21238 9988
rect 23201 9979 23259 9985
rect 23201 9945 23213 9979
rect 23247 9976 23259 9979
rect 23584 9976 23612 10007
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 23247 9948 23612 9976
rect 23768 9976 23796 10084
rect 23860 10053 23888 10220
rect 25056 10124 25084 10220
rect 25685 10217 25697 10251
rect 25731 10248 25743 10251
rect 25731 10220 28396 10248
rect 25731 10217 25743 10220
rect 25685 10211 25743 10217
rect 27982 10140 27988 10192
rect 28040 10180 28046 10192
rect 28258 10180 28264 10192
rect 28040 10152 28264 10180
rect 28040 10140 28046 10152
rect 28258 10140 28264 10152
rect 28316 10140 28322 10192
rect 24118 10112 24124 10124
rect 23952 10084 24124 10112
rect 23952 10053 23980 10084
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 25038 10072 25044 10124
rect 25096 10112 25102 10124
rect 25317 10115 25375 10121
rect 25317 10112 25329 10115
rect 25096 10084 25329 10112
rect 25096 10072 25102 10084
rect 25317 10081 25329 10084
rect 25363 10081 25375 10115
rect 25317 10075 25375 10081
rect 26142 10072 26148 10124
rect 26200 10112 26206 10124
rect 26237 10115 26295 10121
rect 26237 10112 26249 10115
rect 26200 10084 26249 10112
rect 26200 10072 26206 10084
rect 26237 10081 26249 10084
rect 26283 10081 26295 10115
rect 26237 10075 26295 10081
rect 26510 10072 26516 10124
rect 26568 10072 26574 10124
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10013 23903 10047
rect 23845 10007 23903 10013
rect 23937 10047 23995 10053
rect 23937 10013 23949 10047
rect 23983 10013 23995 10047
rect 23937 10007 23995 10013
rect 24034 10047 24092 10053
rect 24034 10013 24046 10047
rect 24080 10013 24092 10047
rect 24949 10047 25007 10053
rect 24949 10044 24961 10047
rect 24034 10007 24092 10013
rect 24228 10016 24961 10044
rect 23952 9976 23980 10007
rect 23768 9948 23980 9976
rect 23247 9945 23259 9948
rect 23201 9939 23259 9945
rect 5408 9880 6132 9908
rect 5408 9868 5414 9880
rect 6454 9868 6460 9920
rect 6512 9868 6518 9920
rect 6638 9868 6644 9920
rect 6696 9868 6702 9920
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9908 7251 9911
rect 8570 9908 8576 9920
rect 7239 9880 8576 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 22830 9868 22836 9920
rect 22888 9908 22894 9920
rect 24044 9908 24072 10007
rect 24228 9917 24256 10016
rect 24949 10013 24961 10016
rect 24995 10013 25007 10047
rect 25133 10047 25191 10053
rect 25133 10044 25145 10047
rect 24949 10007 25007 10013
rect 25056 10016 25145 10044
rect 25056 9988 25084 10016
rect 25133 10013 25145 10016
rect 25179 10013 25191 10047
rect 25133 10007 25191 10013
rect 25225 10047 25283 10053
rect 25225 10013 25237 10047
rect 25271 10013 25283 10047
rect 25225 10007 25283 10013
rect 25038 9936 25044 9988
rect 25096 9936 25102 9988
rect 25240 9976 25268 10007
rect 25498 10004 25504 10056
rect 25556 10004 25562 10056
rect 28074 10004 28080 10056
rect 28132 10046 28138 10056
rect 28132 10018 28175 10046
rect 28132 10004 28138 10018
rect 28258 10004 28264 10056
rect 28316 10004 28322 10056
rect 28368 10053 28396 10220
rect 28442 10208 28448 10260
rect 28500 10248 28506 10260
rect 28905 10251 28963 10257
rect 28905 10248 28917 10251
rect 28500 10220 28917 10248
rect 28500 10208 28506 10220
rect 28905 10217 28917 10220
rect 28951 10217 28963 10251
rect 28905 10211 28963 10217
rect 33134 10208 33140 10260
rect 33192 10208 33198 10260
rect 34514 10208 34520 10260
rect 34572 10248 34578 10260
rect 36817 10251 36875 10257
rect 36817 10248 36829 10251
rect 34572 10220 36829 10248
rect 34572 10208 34578 10220
rect 36817 10217 36829 10220
rect 36863 10217 36875 10251
rect 36817 10211 36875 10217
rect 38562 10208 38568 10260
rect 38620 10208 38626 10260
rect 28813 10183 28871 10189
rect 28813 10149 28825 10183
rect 28859 10180 28871 10183
rect 30837 10183 30895 10189
rect 28859 10152 30788 10180
rect 28859 10149 28871 10152
rect 28813 10143 28871 10149
rect 30098 10072 30104 10124
rect 30156 10072 30162 10124
rect 30190 10072 30196 10124
rect 30248 10112 30254 10124
rect 30248 10084 30604 10112
rect 30248 10072 30254 10084
rect 28353 10047 28411 10053
rect 28353 10013 28365 10047
rect 28399 10013 28411 10047
rect 28353 10007 28411 10013
rect 28445 10047 28503 10053
rect 28445 10013 28457 10047
rect 28491 10013 28503 10047
rect 28445 10007 28503 10013
rect 26602 9976 26608 9988
rect 25240 9948 26608 9976
rect 26602 9936 26608 9948
rect 26660 9936 26666 9988
rect 28166 9976 28172 9988
rect 27738 9948 28172 9976
rect 28166 9936 28172 9948
rect 28224 9936 28230 9988
rect 22888 9880 24072 9908
rect 24213 9911 24271 9917
rect 22888 9868 22894 9880
rect 24213 9877 24225 9911
rect 24259 9877 24271 9911
rect 24213 9871 24271 9877
rect 27338 9868 27344 9920
rect 27396 9908 27402 9920
rect 28460 9908 28488 10007
rect 28534 10004 28540 10056
rect 28592 10044 28598 10056
rect 28629 10047 28687 10053
rect 28629 10044 28641 10047
rect 28592 10016 28641 10044
rect 28592 10004 28598 10016
rect 28629 10013 28641 10016
rect 28675 10013 28687 10047
rect 28629 10007 28687 10013
rect 30285 10047 30343 10053
rect 30285 10013 30297 10047
rect 30331 10044 30343 10047
rect 30374 10044 30380 10056
rect 30331 10016 30380 10044
rect 30331 10013 30343 10016
rect 30285 10007 30343 10013
rect 30374 10004 30380 10016
rect 30432 10004 30438 10056
rect 30576 10053 30604 10084
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10013 30619 10047
rect 30561 10007 30619 10013
rect 30653 10047 30711 10053
rect 30653 10013 30665 10047
rect 30699 10013 30711 10047
rect 30760 10044 30788 10152
rect 30837 10149 30849 10183
rect 30883 10180 30895 10183
rect 31021 10183 31079 10189
rect 31021 10180 31033 10183
rect 30883 10152 31033 10180
rect 30883 10149 30895 10152
rect 30837 10143 30895 10149
rect 31021 10149 31033 10152
rect 31067 10149 31079 10183
rect 31021 10143 31079 10149
rect 32674 10140 32680 10192
rect 32732 10180 32738 10192
rect 34701 10183 34759 10189
rect 34701 10180 34713 10183
rect 32732 10152 33640 10180
rect 32732 10140 32738 10152
rect 31202 10072 31208 10124
rect 31260 10072 31266 10124
rect 31389 10115 31447 10121
rect 31389 10081 31401 10115
rect 31435 10112 31447 10115
rect 31754 10112 31760 10124
rect 31435 10084 31760 10112
rect 31435 10081 31447 10084
rect 31389 10075 31447 10081
rect 31754 10072 31760 10084
rect 31812 10072 31818 10124
rect 32214 10072 32220 10124
rect 32272 10112 32278 10124
rect 32272 10084 32904 10112
rect 32272 10072 32278 10084
rect 30929 10047 30987 10053
rect 30929 10044 30941 10047
rect 30760 10016 30941 10044
rect 30653 10007 30711 10013
rect 30929 10013 30941 10016
rect 30975 10013 30987 10047
rect 32876 10044 32904 10084
rect 33134 10072 33140 10124
rect 33192 10112 33198 10124
rect 33229 10115 33287 10121
rect 33229 10112 33241 10115
rect 33192 10084 33241 10112
rect 33192 10072 33198 10084
rect 33229 10081 33241 10084
rect 33275 10081 33287 10115
rect 33229 10075 33287 10081
rect 33612 10063 33640 10152
rect 34532 10152 34713 10180
rect 34532 10121 34560 10152
rect 34701 10149 34713 10152
rect 34747 10149 34759 10183
rect 34701 10143 34759 10149
rect 37829 10183 37887 10189
rect 37829 10149 37841 10183
rect 37875 10180 37887 10183
rect 37875 10152 37964 10180
rect 37875 10149 37887 10152
rect 37829 10143 37887 10149
rect 34517 10115 34575 10121
rect 34517 10081 34529 10115
rect 34563 10081 34575 10115
rect 34517 10075 34575 10081
rect 34606 10072 34612 10124
rect 34664 10112 34670 10124
rect 35161 10115 35219 10121
rect 35161 10112 35173 10115
rect 34664 10084 35173 10112
rect 34664 10072 34670 10084
rect 35161 10081 35173 10084
rect 35207 10081 35219 10115
rect 35161 10075 35219 10081
rect 35342 10072 35348 10124
rect 35400 10072 35406 10124
rect 35434 10072 35440 10124
rect 35492 10112 35498 10124
rect 36357 10115 36415 10121
rect 36357 10112 36369 10115
rect 35492 10084 36369 10112
rect 35492 10072 35498 10084
rect 36357 10081 36369 10084
rect 36403 10081 36415 10115
rect 37182 10112 37188 10124
rect 36357 10075 36415 10081
rect 36556 10084 37188 10112
rect 33602 10057 33660 10063
rect 33413 10047 33471 10053
rect 33413 10044 33425 10047
rect 32876 10016 33425 10044
rect 30929 10007 30987 10013
rect 33413 10013 33425 10016
rect 33459 10013 33471 10047
rect 33413 10007 33471 10013
rect 29086 9936 29092 9988
rect 29144 9936 29150 9988
rect 29273 9979 29331 9985
rect 29273 9945 29285 9979
rect 29319 9976 29331 9979
rect 29319 9948 29868 9976
rect 29319 9945 29331 9948
rect 29273 9939 29331 9945
rect 27396 9880 28488 9908
rect 27396 9868 27402 9880
rect 29546 9868 29552 9920
rect 29604 9868 29610 9920
rect 29840 9908 29868 9948
rect 30466 9936 30472 9988
rect 30524 9936 30530 9988
rect 30190 9908 30196 9920
rect 29840 9880 30196 9908
rect 30190 9868 30196 9880
rect 30248 9908 30254 9920
rect 30668 9908 30696 10007
rect 33502 10004 33508 10056
rect 33560 10004 33566 10056
rect 33602 10023 33614 10057
rect 33648 10023 33660 10057
rect 33602 10017 33660 10023
rect 36078 10004 36084 10056
rect 36136 10044 36142 10056
rect 36265 10047 36323 10053
rect 36265 10044 36277 10047
rect 36136 10016 36277 10044
rect 36136 10004 36142 10016
rect 36265 10013 36277 10016
rect 36311 10013 36323 10047
rect 36265 10007 36323 10013
rect 36446 10004 36452 10056
rect 36504 10044 36510 10056
rect 36556 10053 36584 10084
rect 37182 10072 37188 10084
rect 37240 10072 37246 10124
rect 37936 10121 37964 10152
rect 37921 10115 37979 10121
rect 37292 10084 37780 10112
rect 36541 10047 36599 10053
rect 36541 10044 36553 10047
rect 36504 10016 36553 10044
rect 36504 10004 36510 10016
rect 36541 10013 36553 10016
rect 36587 10013 36599 10047
rect 36541 10007 36599 10013
rect 36630 10004 36636 10056
rect 36688 10004 36694 10056
rect 37292 10053 37320 10084
rect 37277 10047 37335 10053
rect 37277 10013 37289 10047
rect 37323 10013 37335 10047
rect 37277 10007 37335 10013
rect 37550 10004 37556 10056
rect 37608 10004 37614 10056
rect 37642 10004 37648 10056
rect 37700 10004 37706 10056
rect 37752 10044 37780 10084
rect 37921 10081 37933 10115
rect 37967 10081 37979 10115
rect 37921 10075 37979 10081
rect 38838 10044 38844 10056
rect 37752 10016 38844 10044
rect 38838 10004 38844 10016
rect 38896 10004 38902 10056
rect 38930 10004 38936 10056
rect 38988 10004 38994 10056
rect 39209 10047 39267 10053
rect 39209 10013 39221 10047
rect 39255 10044 39267 10047
rect 39853 10047 39911 10053
rect 39853 10044 39865 10047
rect 39255 10016 39865 10044
rect 39255 10013 39267 10016
rect 39209 10007 39267 10013
rect 39853 10013 39865 10016
rect 39899 10013 39911 10047
rect 39853 10007 39911 10013
rect 40402 10004 40408 10056
rect 40460 10004 40466 10056
rect 31665 9979 31723 9985
rect 31665 9945 31677 9979
rect 31711 9976 31723 9979
rect 31938 9976 31944 9988
rect 31711 9948 31944 9976
rect 31711 9945 31723 9948
rect 31665 9939 31723 9945
rect 31938 9936 31944 9948
rect 31996 9936 32002 9988
rect 33042 9976 33048 9988
rect 32890 9948 33048 9976
rect 33042 9936 33048 9948
rect 33100 9936 33106 9988
rect 33226 9936 33232 9988
rect 33284 9985 33290 9988
rect 33284 9979 33333 9985
rect 33284 9945 33287 9979
rect 33321 9945 33333 9979
rect 33284 9939 33333 9945
rect 35069 9979 35127 9985
rect 35069 9945 35081 9979
rect 35115 9976 35127 9979
rect 35529 9979 35587 9985
rect 35529 9976 35541 9979
rect 35115 9948 35541 9976
rect 35115 9945 35127 9948
rect 35069 9939 35127 9945
rect 35529 9945 35541 9948
rect 35575 9945 35587 9979
rect 35529 9939 35587 9945
rect 33284 9936 33290 9939
rect 36998 9936 37004 9988
rect 37056 9976 37062 9988
rect 37458 9976 37464 9988
rect 37056 9948 37464 9976
rect 37056 9936 37062 9948
rect 37458 9936 37464 9948
rect 37516 9936 37522 9988
rect 39025 9979 39083 9985
rect 39025 9976 39037 9979
rect 37568 9948 39037 9976
rect 30248 9880 30696 9908
rect 31205 9911 31263 9917
rect 30248 9868 30254 9880
rect 31205 9877 31217 9911
rect 31251 9908 31263 9911
rect 32582 9908 32588 9920
rect 31251 9880 32588 9908
rect 31251 9877 31263 9880
rect 31205 9871 31263 9877
rect 32582 9868 32588 9880
rect 32640 9868 32646 9920
rect 33870 9868 33876 9920
rect 33928 9868 33934 9920
rect 37274 9868 37280 9920
rect 37332 9908 37338 9920
rect 37568 9908 37596 9948
rect 39025 9945 39037 9948
rect 39071 9945 39083 9979
rect 39025 9939 39083 9945
rect 37332 9880 37596 9908
rect 37332 9868 37338 9880
rect 38654 9868 38660 9920
rect 38712 9868 38718 9920
rect 39040 9908 39068 9939
rect 39942 9936 39948 9988
rect 40000 9976 40006 9988
rect 40681 9979 40739 9985
rect 40681 9976 40693 9979
rect 40000 9948 40693 9976
rect 40000 9936 40006 9948
rect 40681 9945 40693 9948
rect 40727 9945 40739 9979
rect 40681 9939 40739 9945
rect 40773 9911 40831 9917
rect 40773 9908 40785 9911
rect 39040 9880 40785 9908
rect 40773 9877 40785 9880
rect 40819 9877 40831 9911
rect 40773 9871 40831 9877
rect 1104 9818 42504 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 42504 9818
rect 1104 9744 42504 9766
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 6641 9707 6699 9713
rect 6641 9704 6653 9707
rect 5776 9676 6653 9704
rect 5776 9664 5782 9676
rect 6641 9673 6653 9676
rect 6687 9704 6699 9707
rect 6822 9704 6828 9716
rect 6687 9676 6828 9704
rect 6687 9673 6699 9676
rect 6641 9667 6699 9673
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 8205 9707 8263 9713
rect 8205 9673 8217 9707
rect 8251 9704 8263 9707
rect 8251 9676 8524 9704
rect 8251 9673 8263 9676
rect 8205 9667 8263 9673
rect 3053 9639 3111 9645
rect 3053 9636 3065 9639
rect 2700 9608 3065 9636
rect 2498 9528 2504 9580
rect 2556 9528 2562 9580
rect 2700 9577 2728 9608
rect 3053 9605 3065 9608
rect 3099 9605 3111 9639
rect 6178 9636 6184 9648
rect 3053 9599 3111 9605
rect 5460 9608 5764 9636
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 2976 9500 3004 9531
rect 3142 9528 3148 9580
rect 3200 9528 3206 9580
rect 5258 9528 5264 9580
rect 5316 9528 5322 9580
rect 5460 9577 5488 9608
rect 5736 9580 5764 9608
rect 6012 9608 6184 9636
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9568 5595 9571
rect 5626 9568 5632 9580
rect 5583 9540 5632 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5718 9528 5724 9580
rect 5776 9528 5782 9580
rect 6012 9577 6040 9608
rect 6178 9596 6184 9608
rect 6236 9636 6242 9648
rect 6236 9608 7328 9636
rect 6236 9596 6242 9608
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6638 9571 6696 9577
rect 6638 9537 6650 9571
rect 6684 9568 6696 9571
rect 6914 9568 6920 9580
rect 6684 9540 6920 9568
rect 6684 9537 6696 9540
rect 6638 9531 6696 9537
rect 6914 9528 6920 9540
rect 6972 9568 6978 9580
rect 7300 9577 7328 9608
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 8389 9639 8447 9645
rect 8389 9636 8401 9639
rect 7432 9608 8401 9636
rect 7432 9596 7438 9608
rect 8389 9605 8401 9608
rect 8435 9605 8447 9639
rect 8496 9636 8524 9676
rect 23658 9664 23664 9716
rect 23716 9704 23722 9716
rect 25498 9704 25504 9716
rect 23716 9676 25504 9704
rect 23716 9664 23722 9676
rect 25498 9664 25504 9676
rect 25556 9664 25562 9716
rect 28166 9664 28172 9716
rect 28224 9704 28230 9716
rect 28718 9704 28724 9716
rect 28224 9676 28724 9704
rect 28224 9664 28230 9676
rect 28718 9664 28724 9676
rect 28776 9664 28782 9716
rect 31202 9664 31208 9716
rect 31260 9664 31266 9716
rect 34790 9664 34796 9716
rect 34848 9704 34854 9716
rect 34848 9676 35480 9704
rect 34848 9664 34854 9676
rect 11330 9636 11336 9648
rect 8496 9608 11336 9636
rect 8389 9599 8447 9605
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 20070 9636 20076 9648
rect 19444 9608 20076 9636
rect 7285 9571 7343 9577
rect 6972 9540 7236 9568
rect 6972 9528 6978 9540
rect 3418 9500 3424 9512
rect 2976 9472 3424 9500
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 4672 9472 5825 9500
rect 4672 9460 4678 9472
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9469 7159 9503
rect 7208 9500 7236 9540
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 8294 9528 8300 9580
rect 8352 9528 8358 9580
rect 10045 9571 10103 9577
rect 10045 9537 10057 9571
rect 10091 9568 10103 9571
rect 10134 9568 10140 9580
rect 10091 9540 10140 9568
rect 10091 9537 10103 9540
rect 10045 9531 10103 9537
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 7208 9472 7389 9500
rect 7101 9463 7159 9469
rect 7377 9469 7389 9472
rect 7423 9469 7435 9503
rect 7377 9463 7435 9469
rect 5994 9432 6000 9444
rect 5828 9404 6000 9432
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2501 9367 2559 9373
rect 2501 9364 2513 9367
rect 1728 9336 2513 9364
rect 1728 9324 1734 9336
rect 2501 9333 2513 9336
rect 2547 9333 2559 9367
rect 2501 9327 2559 9333
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 5828 9373 5856 9404
rect 5994 9392 6000 9404
rect 6052 9392 6058 9444
rect 6270 9392 6276 9444
rect 6328 9432 6334 9444
rect 7009 9435 7067 9441
rect 7009 9432 7021 9435
rect 6328 9404 7021 9432
rect 6328 9392 6334 9404
rect 7009 9401 7021 9404
rect 7055 9401 7067 9435
rect 7116 9432 7144 9463
rect 7466 9460 7472 9512
rect 7524 9460 7530 9512
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 8478 9500 8484 9512
rect 7791 9472 8484 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 7282 9432 7288 9444
rect 7116 9404 7288 9432
rect 7009 9395 7067 9401
rect 7282 9392 7288 9404
rect 7340 9392 7346 9444
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 3476 9336 5273 9364
rect 3476 9324 3482 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 5261 9327 5319 9333
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9333 5871 9367
rect 5813 9327 5871 9333
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 5960 9336 6193 9364
rect 5960 9324 5966 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6181 9327 6239 9333
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6420 9336 6469 9364
rect 6420 9324 6426 9336
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 7576 9364 7604 9463
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 8386 9392 8392 9444
rect 8444 9432 8450 9444
rect 8573 9435 8631 9441
rect 8573 9432 8585 9435
rect 8444 9404 8585 9432
rect 8444 9392 8450 9404
rect 8573 9401 8585 9404
rect 8619 9401 8631 9435
rect 10060 9432 10088 9531
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10410 9528 10416 9580
rect 10468 9528 10474 9580
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 11514 9568 11520 9580
rect 11287 9540 11520 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 11514 9528 11520 9540
rect 11572 9568 11578 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11572 9540 11621 9568
rect 11572 9528 11578 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 18414 9528 18420 9580
rect 18472 9528 18478 9580
rect 19444 9577 19472 9608
rect 20070 9596 20076 9608
rect 20128 9636 20134 9648
rect 20533 9639 20591 9645
rect 20533 9636 20545 9639
rect 20128 9608 20545 9636
rect 20128 9596 20134 9608
rect 20533 9605 20545 9608
rect 20579 9605 20591 9639
rect 22002 9636 22008 9648
rect 20533 9599 20591 9605
rect 21468 9608 22008 9636
rect 21468 9580 21496 9608
rect 22002 9596 22008 9608
rect 22060 9596 22066 9648
rect 23198 9636 23204 9648
rect 22862 9608 23204 9636
rect 23198 9596 23204 9608
rect 23256 9596 23262 9648
rect 23293 9639 23351 9645
rect 23293 9605 23305 9639
rect 23339 9636 23351 9639
rect 23750 9636 23756 9648
rect 23339 9608 23756 9636
rect 23339 9605 23351 9608
rect 23293 9599 23351 9605
rect 23750 9596 23756 9608
rect 23808 9596 23814 9648
rect 25682 9636 25688 9648
rect 25346 9608 25688 9636
rect 25682 9596 25688 9608
rect 25740 9596 25746 9648
rect 26602 9596 26608 9648
rect 26660 9636 26666 9648
rect 27249 9639 27307 9645
rect 27249 9636 27261 9639
rect 26660 9608 27261 9636
rect 26660 9596 26666 9608
rect 27249 9605 27261 9608
rect 27295 9605 27307 9639
rect 27249 9599 27307 9605
rect 27338 9596 27344 9648
rect 27396 9596 27402 9648
rect 28810 9596 28816 9648
rect 28868 9596 28874 9648
rect 29457 9639 29515 9645
rect 29457 9605 29469 9639
rect 29503 9636 29515 9639
rect 29546 9636 29552 9648
rect 29503 9608 29552 9636
rect 29503 9605 29515 9608
rect 29457 9599 29515 9605
rect 29546 9596 29552 9608
rect 29604 9596 29610 9648
rect 31754 9636 31760 9648
rect 29748 9608 31248 9636
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 19518 9528 19524 9580
rect 19576 9577 19582 9580
rect 19576 9571 19625 9577
rect 19576 9537 19579 9571
rect 19613 9537 19625 9571
rect 19576 9531 19625 9537
rect 19576 9528 19582 9531
rect 19702 9528 19708 9580
rect 19760 9528 19766 9580
rect 19794 9528 19800 9580
rect 19852 9528 19858 9580
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20165 9571 20223 9577
rect 20165 9568 20177 9571
rect 19935 9540 20177 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 20165 9537 20177 9540
rect 20211 9537 20223 9571
rect 20165 9531 20223 9537
rect 20346 9528 20352 9580
rect 20404 9528 20410 9580
rect 21450 9528 21456 9580
rect 21508 9528 21514 9580
rect 21637 9571 21695 9577
rect 21637 9537 21649 9571
rect 21683 9537 21695 9571
rect 21637 9531 21695 9537
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9500 10379 9503
rect 12158 9500 12164 9512
rect 10367 9472 12164 9500
rect 10367 9469 10379 9472
rect 10321 9463 10379 9469
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9500 20131 9503
rect 21358 9500 21364 9512
rect 20119 9472 21364 9500
rect 20119 9469 20131 9472
rect 20073 9463 20131 9469
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 21652 9500 21680 9531
rect 26694 9528 26700 9580
rect 26752 9528 26758 9580
rect 27154 9528 27160 9580
rect 27212 9528 27218 9580
rect 27525 9571 27583 9577
rect 27525 9537 27537 9571
rect 27571 9568 27583 9571
rect 27982 9568 27988 9580
rect 27571 9540 27988 9568
rect 27571 9537 27583 9540
rect 27525 9531 27583 9537
rect 27982 9528 27988 9540
rect 28040 9528 28046 9580
rect 29748 9577 29776 9608
rect 29733 9571 29791 9577
rect 29733 9537 29745 9571
rect 29779 9537 29791 9571
rect 29733 9531 29791 9537
rect 30374 9528 30380 9580
rect 30432 9568 30438 9580
rect 30653 9571 30711 9577
rect 30653 9568 30665 9571
rect 30432 9540 30665 9568
rect 30432 9528 30438 9540
rect 30653 9537 30665 9540
rect 30699 9537 30711 9571
rect 30653 9531 30711 9537
rect 30834 9528 30840 9580
rect 30892 9568 30898 9580
rect 30929 9571 30987 9577
rect 30929 9568 30941 9571
rect 30892 9540 30941 9568
rect 30892 9528 30898 9540
rect 30929 9537 30941 9540
rect 30975 9537 30987 9571
rect 30929 9531 30987 9537
rect 31021 9571 31079 9577
rect 31021 9537 31033 9571
rect 31067 9537 31079 9571
rect 31220 9568 31248 9608
rect 31680 9608 31760 9636
rect 31680 9568 31708 9608
rect 31754 9596 31760 9608
rect 31812 9596 31818 9648
rect 32125 9639 32183 9645
rect 32125 9605 32137 9639
rect 32171 9636 32183 9639
rect 32398 9636 32404 9648
rect 32171 9608 32404 9636
rect 32171 9605 32183 9608
rect 32125 9599 32183 9605
rect 32398 9596 32404 9608
rect 32456 9596 32462 9648
rect 33870 9596 33876 9648
rect 33928 9596 33934 9648
rect 35452 9645 35480 9676
rect 37642 9664 37648 9716
rect 37700 9704 37706 9716
rect 38289 9707 38347 9713
rect 38289 9704 38301 9707
rect 37700 9676 38301 9704
rect 37700 9664 37706 9676
rect 38289 9673 38301 9676
rect 38335 9673 38347 9707
rect 38289 9667 38347 9673
rect 38378 9664 38384 9716
rect 38436 9704 38442 9716
rect 38436 9676 39068 9704
rect 38436 9664 38442 9676
rect 35437 9639 35495 9645
rect 35437 9605 35449 9639
rect 35483 9605 35495 9639
rect 35437 9599 35495 9605
rect 35986 9596 35992 9648
rect 36044 9636 36050 9648
rect 36173 9639 36231 9645
rect 36173 9636 36185 9639
rect 36044 9608 36185 9636
rect 36044 9596 36050 9608
rect 36173 9605 36185 9608
rect 36219 9605 36231 9639
rect 36173 9599 36231 9605
rect 36446 9596 36452 9648
rect 36504 9596 36510 9648
rect 38654 9596 38660 9648
rect 38712 9636 38718 9648
rect 38933 9639 38991 9645
rect 38933 9636 38945 9639
rect 38712 9608 38945 9636
rect 38712 9596 38718 9608
rect 38933 9605 38945 9608
rect 38979 9605 38991 9639
rect 39040 9636 39068 9676
rect 39040 9608 39422 9636
rect 38933 9599 38991 9605
rect 31849 9571 31907 9577
rect 31849 9568 31861 9571
rect 31220 9540 31861 9568
rect 31021 9531 31079 9537
rect 31849 9537 31861 9540
rect 31895 9537 31907 9571
rect 31849 9531 31907 9537
rect 21726 9500 21732 9512
rect 21652 9472 21732 9500
rect 21726 9460 21732 9472
rect 21784 9500 21790 9512
rect 23290 9500 23296 9512
rect 21784 9472 23296 9500
rect 21784 9460 21790 9472
rect 23290 9460 23296 9472
rect 23348 9460 23354 9512
rect 23566 9460 23572 9512
rect 23624 9500 23630 9512
rect 23845 9503 23903 9509
rect 23845 9500 23857 9503
rect 23624 9472 23857 9500
rect 23624 9460 23630 9472
rect 23845 9469 23857 9472
rect 23891 9469 23903 9503
rect 23845 9463 23903 9469
rect 24121 9503 24179 9509
rect 24121 9469 24133 9503
rect 24167 9500 24179 9503
rect 24578 9500 24584 9512
rect 24167 9472 24584 9500
rect 24167 9469 24179 9472
rect 24121 9463 24179 9469
rect 24578 9460 24584 9472
rect 24636 9460 24642 9512
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9500 25651 9503
rect 26237 9503 26295 9509
rect 26237 9500 26249 9503
rect 25639 9472 26249 9500
rect 25639 9469 25651 9472
rect 25593 9463 25651 9469
rect 26237 9469 26249 9472
rect 26283 9469 26295 9503
rect 26237 9463 26295 9469
rect 12250 9432 12256 9444
rect 10060 9404 12256 9432
rect 8573 9395 8631 9401
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 21269 9435 21327 9441
rect 21269 9401 21281 9435
rect 21315 9432 21327 9435
rect 22278 9432 22284 9444
rect 21315 9404 22284 9432
rect 21315 9401 21327 9404
rect 21269 9395 21327 9401
rect 22278 9392 22284 9404
rect 22336 9392 22342 9444
rect 25406 9392 25412 9444
rect 25464 9432 25470 9444
rect 26513 9435 26571 9441
rect 26513 9432 26525 9435
rect 25464 9404 26525 9432
rect 25464 9392 25470 9404
rect 26513 9401 26525 9404
rect 26559 9401 26571 9435
rect 26513 9395 26571 9401
rect 26973 9435 27031 9441
rect 26973 9401 26985 9435
rect 27019 9432 27031 9435
rect 28258 9432 28264 9444
rect 27019 9404 28264 9432
rect 27019 9401 27031 9404
rect 26973 9395 27031 9401
rect 6880 9336 7604 9364
rect 6880 9324 6886 9336
rect 8018 9324 8024 9376
rect 8076 9324 8082 9376
rect 10134 9324 10140 9376
rect 10192 9324 10198 9376
rect 10226 9324 10232 9376
rect 10284 9324 10290 9376
rect 21634 9324 21640 9376
rect 21692 9324 21698 9376
rect 21821 9367 21879 9373
rect 21821 9333 21833 9367
rect 21867 9364 21879 9367
rect 22094 9364 22100 9376
rect 21867 9336 22100 9364
rect 21867 9333 21879 9336
rect 21821 9327 21879 9333
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 25130 9324 25136 9376
rect 25188 9364 25194 9376
rect 25685 9367 25743 9373
rect 25685 9364 25697 9367
rect 25188 9336 25697 9364
rect 25188 9324 25194 9336
rect 25685 9333 25697 9336
rect 25731 9333 25743 9367
rect 26528 9364 26556 9395
rect 28258 9392 28264 9404
rect 28316 9392 28322 9444
rect 31036 9432 31064 9531
rect 31864 9500 31892 9531
rect 32953 9503 33011 9509
rect 32953 9500 32965 9503
rect 31864 9472 32965 9500
rect 32953 9469 32965 9472
rect 32999 9500 33011 9503
rect 33042 9500 33048 9512
rect 32999 9472 33048 9500
rect 32999 9469 33011 9472
rect 32953 9463 33011 9469
rect 33042 9460 33048 9472
rect 33100 9500 33106 9512
rect 33597 9503 33655 9509
rect 33597 9500 33609 9503
rect 33100 9472 33609 9500
rect 33100 9460 33106 9472
rect 33597 9469 33609 9472
rect 33643 9469 33655 9503
rect 33597 9463 33655 9469
rect 32674 9432 32680 9444
rect 31036 9404 32680 9432
rect 32674 9392 32680 9404
rect 32732 9392 32738 9444
rect 27614 9364 27620 9376
rect 26528 9336 27620 9364
rect 25685 9327 25743 9333
rect 27614 9324 27620 9336
rect 27672 9324 27678 9376
rect 27985 9367 28043 9373
rect 27985 9333 27997 9367
rect 28031 9364 28043 9367
rect 29086 9364 29092 9376
rect 28031 9336 29092 9364
rect 28031 9333 28043 9336
rect 27985 9327 28043 9333
rect 29086 9324 29092 9336
rect 29144 9324 29150 9376
rect 29822 9324 29828 9376
rect 29880 9364 29886 9376
rect 30466 9364 30472 9376
rect 29880 9336 30472 9364
rect 29880 9324 29886 9336
rect 30466 9324 30472 9336
rect 30524 9364 30530 9376
rect 30745 9367 30803 9373
rect 30745 9364 30757 9367
rect 30524 9336 30757 9364
rect 30524 9324 30530 9336
rect 30745 9333 30757 9336
rect 30791 9333 30803 9367
rect 30745 9327 30803 9333
rect 30834 9324 30840 9376
rect 30892 9364 30898 9376
rect 33318 9364 33324 9376
rect 30892 9336 33324 9364
rect 30892 9324 30898 9336
rect 33318 9324 33324 9336
rect 33376 9324 33382 9376
rect 34992 9364 35020 9554
rect 35526 9528 35532 9580
rect 35584 9568 35590 9580
rect 35621 9571 35679 9577
rect 35621 9568 35633 9571
rect 35584 9540 35633 9568
rect 35584 9528 35590 9540
rect 35621 9537 35633 9540
rect 35667 9537 35679 9571
rect 35621 9531 35679 9537
rect 36354 9528 36360 9580
rect 36412 9528 36418 9580
rect 36538 9568 36544 9580
rect 36596 9577 36602 9580
rect 36504 9540 36544 9568
rect 36538 9528 36544 9540
rect 36596 9531 36604 9577
rect 37737 9571 37795 9577
rect 37737 9537 37749 9571
rect 37783 9537 37795 9571
rect 38197 9571 38255 9577
rect 38197 9568 38209 9571
rect 37737 9531 37795 9537
rect 38120 9540 38209 9568
rect 36596 9528 36602 9531
rect 35345 9503 35403 9509
rect 35345 9469 35357 9503
rect 35391 9500 35403 9503
rect 35805 9503 35863 9509
rect 35805 9500 35817 9503
rect 35391 9472 35817 9500
rect 35391 9469 35403 9472
rect 35345 9463 35403 9469
rect 35805 9469 35817 9472
rect 35851 9500 35863 9503
rect 36078 9500 36084 9512
rect 35851 9472 36084 9500
rect 35851 9469 35863 9472
rect 35805 9463 35863 9469
rect 36078 9460 36084 9472
rect 36136 9460 36142 9512
rect 36170 9392 36176 9444
rect 36228 9392 36234 9444
rect 36262 9364 36268 9376
rect 34992 9336 36268 9364
rect 36262 9324 36268 9336
rect 36320 9324 36326 9376
rect 37752 9364 37780 9531
rect 38120 9509 38148 9540
rect 38197 9537 38209 9540
rect 38243 9537 38255 9571
rect 38197 9531 38255 9537
rect 37829 9503 37887 9509
rect 37829 9469 37841 9503
rect 37875 9469 37887 9503
rect 37829 9463 37887 9469
rect 38105 9503 38163 9509
rect 38105 9469 38117 9503
rect 38151 9469 38163 9503
rect 38105 9463 38163 9469
rect 37844 9432 37872 9463
rect 38654 9460 38660 9512
rect 38712 9460 38718 9512
rect 40402 9500 40408 9512
rect 38764 9472 40408 9500
rect 38562 9432 38568 9444
rect 37844 9404 38568 9432
rect 38562 9392 38568 9404
rect 38620 9392 38626 9444
rect 38764 9432 38792 9472
rect 40402 9460 40408 9472
rect 40460 9460 40466 9512
rect 38679 9404 38792 9432
rect 38679 9364 38707 9404
rect 37752 9336 38707 9364
rect 1104 9274 42504 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 42504 9274
rect 1104 9200 42504 9222
rect 3970 9160 3976 9172
rect 3620 9132 3976 9160
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2958 9024 2964 9036
rect 1443 8996 2964 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 3620 9033 3648 9132
rect 3970 9120 3976 9132
rect 4028 9160 4034 9172
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 4028 9132 4537 9160
rect 4028 9120 4034 9132
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 4525 9123 4583 9129
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 6236 9132 6469 9160
rect 6236 9120 6242 9132
rect 6457 9129 6469 9132
rect 6503 9129 6515 9163
rect 6457 9123 6515 9129
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 6641 9163 6699 9169
rect 6641 9160 6653 9163
rect 6604 9132 6653 9160
rect 6604 9120 6610 9132
rect 6641 9129 6653 9132
rect 6687 9129 6699 9163
rect 6641 9123 6699 9129
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 7524 9132 9045 9160
rect 7524 9120 7530 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9756 9163 9814 9169
rect 9756 9129 9768 9163
rect 9802 9160 9814 9163
rect 10226 9160 10232 9172
rect 9802 9132 10232 9160
rect 9802 9129 9814 9132
rect 9756 9123 9814 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 12158 9120 12164 9172
rect 12216 9120 12222 9172
rect 17576 9163 17634 9169
rect 17576 9129 17588 9163
rect 17622 9160 17634 9163
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 17622 9132 19257 9160
rect 17622 9129 17634 9132
rect 17576 9123 17634 9129
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 21726 9120 21732 9172
rect 21784 9160 21790 9172
rect 21913 9163 21971 9169
rect 21913 9160 21925 9163
rect 21784 9132 21925 9160
rect 21784 9120 21790 9132
rect 21913 9129 21925 9132
rect 21959 9129 21971 9163
rect 22370 9160 22376 9172
rect 21913 9123 21971 9129
rect 22066 9132 22376 9160
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 5261 9095 5319 9101
rect 3844 9064 4660 9092
rect 3844 9052 3850 9064
rect 4632 9033 4660 9064
rect 5261 9061 5273 9095
rect 5307 9092 5319 9095
rect 5307 9064 6776 9092
rect 5307 9061 5319 9064
rect 5261 9055 5319 9061
rect 3605 9027 3663 9033
rect 3605 9024 3617 9027
rect 3200 8996 3617 9024
rect 3200 8984 3206 8996
rect 3605 8993 3617 8996
rect 3651 8993 3663 9027
rect 3605 8987 3663 8993
rect 4617 9027 4675 9033
rect 4617 8993 4629 9027
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 5534 8984 5540 9036
rect 5592 8984 5598 9036
rect 5902 8984 5908 9036
rect 5960 8984 5966 9036
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 9024 6055 9027
rect 6362 9024 6368 9036
rect 6043 8996 6368 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 2806 8928 3372 8956
rect 1670 8848 1676 8900
rect 1728 8848 1734 8900
rect 3237 8891 3295 8897
rect 3237 8888 3249 8891
rect 2976 8860 3249 8888
rect 1946 8780 1952 8832
rect 2004 8820 2010 8832
rect 2498 8820 2504 8832
rect 2004 8792 2504 8820
rect 2004 8780 2010 8792
rect 2498 8780 2504 8792
rect 2556 8820 2562 8832
rect 2976 8820 3004 8860
rect 3237 8857 3249 8860
rect 3283 8857 3295 8891
rect 3344 8888 3372 8928
rect 3418 8916 3424 8968
rect 3476 8916 3482 8968
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8956 4491 8959
rect 4706 8956 4712 8968
rect 4479 8928 4712 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 4706 8916 4712 8928
rect 4764 8956 4770 8968
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 4764 8928 4813 8956
rect 4764 8916 4770 8928
rect 4801 8925 4813 8928
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 3694 8888 3700 8900
rect 3344 8860 3700 8888
rect 3237 8851 3295 8857
rect 3694 8848 3700 8860
rect 3752 8848 3758 8900
rect 3878 8848 3884 8900
rect 3936 8888 3942 8900
rect 4525 8891 4583 8897
rect 4525 8888 4537 8891
rect 3936 8860 4537 8888
rect 3936 8848 3942 8860
rect 4525 8857 4537 8860
rect 4571 8857 4583 8891
rect 5276 8888 5304 8919
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5408 8928 5457 8956
rect 5408 8916 5414 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 5810 8916 5816 8968
rect 5868 8956 5874 8968
rect 6273 8959 6331 8965
rect 6273 8956 6285 8959
rect 5868 8928 6285 8956
rect 5868 8916 5874 8928
rect 6273 8925 6285 8928
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6546 8956 6552 8968
rect 6503 8928 6552 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6748 8956 6776 9064
rect 19518 9052 19524 9104
rect 19576 9092 19582 9104
rect 19981 9095 20039 9101
rect 19981 9092 19993 9095
rect 19576 9064 19993 9092
rect 19576 9052 19582 9064
rect 19981 9061 19993 9064
rect 20027 9061 20039 9095
rect 22066 9092 22094 9132
rect 22370 9120 22376 9132
rect 22428 9160 22434 9172
rect 22557 9163 22615 9169
rect 22557 9160 22569 9163
rect 22428 9132 22569 9160
rect 22428 9120 22434 9132
rect 22557 9129 22569 9132
rect 22603 9129 22615 9163
rect 22557 9123 22615 9129
rect 22738 9120 22744 9172
rect 22796 9160 22802 9172
rect 23382 9160 23388 9172
rect 22796 9132 23388 9160
rect 22796 9120 22802 9132
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 24578 9120 24584 9172
rect 24636 9120 24642 9172
rect 32214 9120 32220 9172
rect 32272 9120 32278 9172
rect 32769 9163 32827 9169
rect 32769 9129 32781 9163
rect 32815 9160 32827 9163
rect 34330 9160 34336 9172
rect 32815 9132 34336 9160
rect 32815 9129 32827 9132
rect 32769 9123 32827 9129
rect 34330 9120 34336 9132
rect 34388 9120 34394 9172
rect 36354 9120 36360 9172
rect 36412 9160 36418 9172
rect 38565 9163 38623 9169
rect 38565 9160 38577 9163
rect 36412 9132 38577 9160
rect 36412 9120 36418 9132
rect 38565 9129 38577 9132
rect 38611 9129 38623 9163
rect 38565 9123 38623 9129
rect 19981 9055 20039 9061
rect 21468 9064 22094 9092
rect 22281 9095 22339 9101
rect 6822 8984 6828 9036
rect 6880 8984 6886 9036
rect 7285 9027 7343 9033
rect 7285 8993 7297 9027
rect 7331 9024 7343 9027
rect 8018 9024 8024 9036
rect 7331 8996 8024 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 9364 8996 9505 9024
rect 9364 8984 9370 8996
rect 9493 8993 9505 8996
rect 9539 9024 9551 9027
rect 11054 9024 11060 9036
rect 9539 8996 11060 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 11054 8984 11060 8996
rect 11112 9024 11118 9036
rect 11514 9024 11520 9036
rect 11112 8996 11520 9024
rect 11112 8984 11118 8996
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 12713 9027 12771 9033
rect 11756 8996 12296 9024
rect 11756 8984 11762 8996
rect 6914 8956 6920 8968
rect 6748 8928 6920 8956
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8386 8956 8392 8968
rect 8251 8928 8392 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9398 8956 9404 8968
rect 9263 8928 9404 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 6086 8888 6092 8900
rect 4525 8851 4583 8857
rect 5000 8860 6092 8888
rect 2556 8792 3004 8820
rect 2556 8780 2562 8792
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 5000 8829 5028 8860
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 6181 8891 6239 8897
rect 6181 8857 6193 8891
rect 6227 8888 6239 8891
rect 6730 8888 6736 8900
rect 6227 8860 6736 8888
rect 6227 8857 6239 8860
rect 6181 8851 6239 8857
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 9048 8888 9076 8919
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 12268 8965 12296 8996
rect 12713 8993 12725 9027
rect 12759 9024 12771 9027
rect 12802 9024 12808 9036
rect 12759 8996 12808 9024
rect 12759 8993 12771 8996
rect 12713 8987 12771 8993
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 11256 8928 11345 8956
rect 10042 8888 10048 8900
rect 9048 8860 10048 8888
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 10318 8848 10324 8900
rect 10376 8848 10382 8900
rect 11256 8832 11284 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 12023 8928 12081 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 12253 8959 12311 8965
rect 12253 8925 12265 8959
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 12268 8888 12296 8919
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 13004 8956 13032 8987
rect 15286 8984 15292 9036
rect 15344 9024 15350 9036
rect 15838 9024 15844 9036
rect 15344 8996 15844 9024
rect 15344 8984 15350 8996
rect 15838 8984 15844 8996
rect 15896 9024 15902 9036
rect 17313 9027 17371 9033
rect 17313 9024 17325 9027
rect 15896 8996 17325 9024
rect 15896 8984 15902 8996
rect 17313 8993 17325 8996
rect 17359 9024 17371 9027
rect 18322 9024 18328 9036
rect 17359 8996 18328 9024
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 19392 8996 19441 9024
rect 19392 8984 19398 8996
rect 19429 8993 19441 8996
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 19702 8984 19708 9036
rect 19760 9024 19766 9036
rect 20441 9027 20499 9033
rect 20441 9024 20453 9027
rect 19760 8996 20453 9024
rect 19760 8984 19766 8996
rect 20441 8993 20453 8996
rect 20487 9024 20499 9027
rect 21468 9024 21496 9064
rect 22281 9061 22293 9095
rect 22327 9092 22339 9095
rect 22646 9092 22652 9104
rect 22327 9064 22652 9092
rect 22327 9061 22339 9064
rect 22281 9055 22339 9061
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 22922 9052 22928 9104
rect 22980 9092 22986 9104
rect 24210 9092 24216 9104
rect 22980 9064 24216 9092
rect 22980 9052 22986 9064
rect 24210 9052 24216 9064
rect 24268 9092 24274 9104
rect 33226 9092 33232 9104
rect 24268 9064 25268 9092
rect 24268 9052 24274 9064
rect 20487 8996 21496 9024
rect 20487 8993 20499 8996
rect 20441 8987 20499 8993
rect 12400 8928 13032 8956
rect 12400 8916 12406 8928
rect 13078 8916 13084 8968
rect 13136 8916 13142 8968
rect 19518 8916 19524 8968
rect 19576 8916 19582 8968
rect 20162 8956 20168 8968
rect 19720 8928 20168 8956
rect 13170 8888 13176 8900
rect 12268 8860 13176 8888
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 19720 8888 19748 8928
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 20346 8916 20352 8968
rect 20404 8916 20410 8968
rect 21468 8965 21496 8996
rect 21634 8984 21640 9036
rect 21692 9024 21698 9036
rect 21821 9027 21879 9033
rect 21821 9024 21833 9027
rect 21692 8996 21833 9024
rect 21692 8984 21698 8996
rect 21821 8993 21833 8996
rect 21867 9024 21879 9027
rect 22738 9024 22744 9036
rect 21867 8996 22744 9024
rect 21867 8993 21879 8996
rect 21821 8987 21879 8993
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 21560 8928 21864 8956
rect 18814 8860 19748 8888
rect 19794 8848 19800 8900
rect 19852 8848 19858 8900
rect 19889 8891 19947 8897
rect 19889 8857 19901 8891
rect 19935 8888 19947 8891
rect 19978 8888 19984 8900
rect 19935 8860 19984 8888
rect 19935 8857 19947 8860
rect 19889 8851 19947 8857
rect 19978 8848 19984 8860
rect 20036 8848 20042 8900
rect 20364 8888 20392 8916
rect 21560 8897 21588 8928
rect 21545 8891 21603 8897
rect 21545 8888 21557 8891
rect 20364 8860 21557 8888
rect 21545 8857 21557 8860
rect 21591 8857 21603 8891
rect 21545 8851 21603 8857
rect 21729 8891 21787 8897
rect 21729 8857 21741 8891
rect 21775 8857 21787 8891
rect 21836 8888 21864 8928
rect 22002 8916 22008 8968
rect 22060 8956 22066 8968
rect 22097 8959 22155 8965
rect 22097 8956 22109 8959
rect 22060 8928 22109 8956
rect 22060 8916 22066 8928
rect 22097 8925 22109 8928
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22278 8916 22284 8968
rect 22336 8956 22342 8968
rect 22940 8956 22968 9052
rect 25130 8984 25136 9036
rect 25188 8984 25194 9036
rect 25240 9033 25268 9064
rect 32140 9064 33232 9092
rect 25225 9027 25283 9033
rect 25225 8993 25237 9027
rect 25271 9024 25283 9027
rect 25406 9024 25412 9036
rect 25271 8996 25412 9024
rect 25271 8993 25283 8996
rect 25225 8987 25283 8993
rect 25406 8984 25412 8996
rect 25464 8984 25470 9036
rect 26418 8984 26424 9036
rect 26476 9024 26482 9036
rect 27065 9027 27123 9033
rect 27065 9024 27077 9027
rect 26476 8996 27077 9024
rect 26476 8984 26482 8996
rect 27065 8993 27077 8996
rect 27111 8993 27123 9027
rect 27065 8987 27123 8993
rect 29733 9027 29791 9033
rect 29733 8993 29745 9027
rect 29779 9024 29791 9027
rect 30006 9024 30012 9036
rect 29779 8996 30012 9024
rect 29779 8993 29791 8996
rect 29733 8987 29791 8993
rect 30006 8984 30012 8996
rect 30064 8984 30070 9036
rect 32140 9033 32168 9064
rect 33226 9052 33232 9064
rect 33284 9052 33290 9104
rect 33318 9052 33324 9104
rect 33376 9092 33382 9104
rect 36722 9092 36728 9104
rect 33376 9064 36728 9092
rect 33376 9052 33382 9064
rect 36722 9052 36728 9064
rect 36780 9092 36786 9104
rect 37645 9095 37703 9101
rect 36780 9064 37504 9092
rect 36780 9052 36786 9064
rect 32125 9027 32183 9033
rect 32125 8993 32137 9027
rect 32171 8993 32183 9027
rect 32950 9024 32956 9036
rect 32125 8987 32183 8993
rect 32784 8996 32956 9024
rect 22336 8928 22968 8956
rect 22336 8916 22342 8928
rect 24762 8916 24768 8968
rect 24820 8916 24826 8968
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8956 24915 8959
rect 25038 8956 25044 8968
rect 24903 8928 25044 8956
rect 24903 8925 24915 8928
rect 24857 8919 24915 8925
rect 25038 8916 25044 8928
rect 25096 8956 25102 8968
rect 25096 8928 25544 8956
rect 25096 8916 25102 8928
rect 22373 8891 22431 8897
rect 22373 8888 22385 8891
rect 21836 8860 22385 8888
rect 21729 8851 21787 8857
rect 22373 8857 22385 8860
rect 22419 8857 22431 8891
rect 22373 8851 22431 8857
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3384 8792 3801 8820
rect 3384 8780 3390 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8789 5043 8823
rect 4985 8783 5043 8789
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 6546 8820 6552 8832
rect 5592 8792 6552 8820
rect 5592 8780 5598 8792
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 8757 8823 8815 8829
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 9030 8820 9036 8832
rect 8803 8792 9036 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 11238 8780 11244 8832
rect 11296 8780 11302 8832
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 12986 8820 12992 8832
rect 11756 8792 12992 8820
rect 11756 8780 11762 8792
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 19058 8780 19064 8832
rect 19116 8780 19122 8832
rect 21744 8820 21772 8851
rect 22462 8848 22468 8900
rect 22520 8888 22526 8900
rect 22589 8891 22647 8897
rect 22589 8888 22601 8891
rect 22520 8860 22601 8888
rect 22520 8848 22526 8860
rect 22589 8857 22601 8860
rect 22635 8888 22647 8891
rect 23014 8888 23020 8900
rect 22635 8860 23020 8888
rect 22635 8857 22647 8860
rect 22589 8851 22647 8857
rect 23014 8848 23020 8860
rect 23072 8848 23078 8900
rect 22094 8820 22100 8832
rect 21744 8792 22100 8820
rect 22094 8780 22100 8792
rect 22152 8820 22158 8832
rect 22480 8820 22508 8848
rect 22152 8792 22508 8820
rect 22152 8780 22158 8792
rect 25038 8780 25044 8832
rect 25096 8820 25102 8832
rect 25317 8823 25375 8829
rect 25317 8820 25329 8823
rect 25096 8792 25329 8820
rect 25096 8780 25102 8792
rect 25317 8789 25329 8792
rect 25363 8789 25375 8823
rect 25516 8820 25544 8928
rect 25682 8916 25688 8968
rect 25740 8916 25746 8968
rect 29822 8916 29828 8968
rect 29880 8916 29886 8968
rect 32644 8959 32702 8965
rect 32644 8925 32656 8959
rect 32690 8956 32702 8959
rect 32784 8956 32812 8996
rect 32950 8984 32956 8996
rect 33008 8984 33014 9036
rect 33336 9024 33364 9052
rect 36354 9024 36360 9036
rect 33152 8996 33364 9024
rect 36280 8996 36360 9024
rect 32690 8928 32812 8956
rect 32690 8925 32702 8928
rect 32644 8919 32702 8925
rect 32858 8916 32864 8968
rect 32916 8916 32922 8968
rect 26786 8848 26792 8900
rect 26844 8848 26850 8900
rect 26878 8848 26884 8900
rect 26936 8888 26942 8900
rect 29914 8888 29920 8900
rect 26936 8860 29920 8888
rect 26936 8848 26942 8860
rect 29914 8848 29920 8860
rect 29972 8848 29978 8900
rect 30098 8848 30104 8900
rect 30156 8848 30162 8900
rect 30193 8891 30251 8897
rect 30193 8857 30205 8891
rect 30239 8888 30251 8891
rect 30282 8888 30288 8900
rect 30239 8860 30288 8888
rect 30239 8857 30251 8860
rect 30193 8851 30251 8857
rect 30282 8848 30288 8860
rect 30340 8848 30346 8900
rect 31846 8848 31852 8900
rect 31904 8888 31910 8900
rect 33152 8897 33180 8996
rect 33226 8916 33232 8968
rect 33284 8965 33290 8968
rect 33284 8959 33311 8965
rect 33299 8925 33311 8959
rect 33284 8919 33311 8925
rect 33284 8916 33290 8919
rect 36170 8916 36176 8968
rect 36228 8916 36234 8968
rect 36280 8965 36308 8996
rect 36354 8984 36360 8996
rect 36412 8984 36418 9036
rect 36446 8984 36452 9036
rect 36504 9024 36510 9036
rect 36633 9027 36691 9033
rect 36633 9024 36645 9027
rect 36504 8996 36645 9024
rect 36504 8984 36510 8996
rect 36633 8993 36645 8996
rect 36679 9024 36691 9027
rect 36998 9024 37004 9036
rect 36679 8996 37004 9024
rect 36679 8993 36691 8996
rect 36633 8987 36691 8993
rect 36998 8984 37004 8996
rect 37056 8984 37062 9036
rect 37476 9024 37504 9064
rect 37645 9061 37657 9095
rect 37691 9092 37703 9095
rect 37691 9064 37780 9092
rect 37691 9061 37703 9064
rect 37645 9055 37703 9061
rect 37752 9033 37780 9064
rect 37737 9027 37795 9033
rect 37476 8996 37688 9024
rect 36265 8959 36323 8965
rect 36265 8925 36277 8959
rect 36311 8925 36323 8959
rect 36265 8919 36323 8925
rect 36372 8928 36676 8956
rect 33045 8891 33103 8897
rect 33045 8888 33057 8891
rect 31904 8860 33057 8888
rect 31904 8848 31910 8860
rect 33045 8857 33057 8860
rect 33091 8857 33103 8891
rect 33045 8851 33103 8857
rect 33137 8891 33195 8897
rect 33137 8857 33149 8891
rect 33183 8857 33195 8891
rect 36372 8888 36400 8928
rect 33137 8851 33195 8857
rect 33244 8860 36400 8888
rect 36541 8891 36599 8897
rect 27154 8820 27160 8832
rect 25516 8792 27160 8820
rect 25317 8783 25375 8789
rect 27154 8780 27160 8792
rect 27212 8780 27218 8832
rect 29549 8823 29607 8829
rect 29549 8789 29561 8823
rect 29595 8820 29607 8823
rect 29730 8820 29736 8832
rect 29595 8792 29736 8820
rect 29595 8789 29607 8792
rect 29549 8783 29607 8789
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 32582 8780 32588 8832
rect 32640 8780 32646 8832
rect 33060 8820 33088 8851
rect 33244 8820 33272 8860
rect 36541 8857 36553 8891
rect 36587 8857 36599 8891
rect 36648 8888 36676 8928
rect 37090 8916 37096 8968
rect 37148 8916 37154 8968
rect 37274 8956 37280 8968
rect 37200 8928 37280 8956
rect 37200 8888 37228 8928
rect 37274 8916 37280 8928
rect 37332 8916 37338 8968
rect 37458 8916 37464 8968
rect 37516 8916 37522 8968
rect 36648 8860 37228 8888
rect 37369 8891 37427 8897
rect 36541 8851 36599 8857
rect 37369 8857 37381 8891
rect 37415 8888 37427 8891
rect 37660 8888 37688 8996
rect 37737 8993 37749 9027
rect 37783 8993 37795 9027
rect 37737 8987 37795 8993
rect 38010 8916 38016 8968
rect 38068 8956 38074 8968
rect 38473 8959 38531 8965
rect 38473 8956 38485 8959
rect 38068 8928 38485 8956
rect 38068 8916 38074 8928
rect 38473 8925 38485 8928
rect 38519 8925 38531 8959
rect 38473 8919 38531 8925
rect 38654 8916 38660 8968
rect 38712 8916 38718 8968
rect 38930 8888 38936 8900
rect 37415 8860 38936 8888
rect 37415 8857 37427 8860
rect 37369 8851 37427 8857
rect 33060 8792 33272 8820
rect 33413 8823 33471 8829
rect 33413 8789 33425 8823
rect 33459 8820 33471 8823
rect 34238 8820 34244 8832
rect 33459 8792 34244 8820
rect 33459 8789 33471 8792
rect 33413 8783 33471 8789
rect 34238 8780 34244 8792
rect 34296 8780 34302 8832
rect 35986 8780 35992 8832
rect 36044 8780 36050 8832
rect 36556 8820 36584 8851
rect 38930 8848 38936 8860
rect 38988 8848 38994 8900
rect 37458 8820 37464 8832
rect 36556 8792 37464 8820
rect 37458 8780 37464 8792
rect 37516 8780 37522 8832
rect 38381 8823 38439 8829
rect 38381 8789 38393 8823
rect 38427 8820 38439 8823
rect 38470 8820 38476 8832
rect 38427 8792 38476 8820
rect 38427 8789 38439 8792
rect 38381 8783 38439 8789
rect 38470 8780 38476 8792
rect 38528 8780 38534 8832
rect 1104 8730 42504 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 42504 8730
rect 1104 8656 42504 8678
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6270 8616 6276 8628
rect 6227 8588 6276 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6365 8619 6423 8625
rect 6365 8585 6377 8619
rect 6411 8616 6423 8619
rect 6638 8616 6644 8628
rect 6411 8588 6644 8616
rect 6411 8585 6423 8588
rect 6365 8579 6423 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 8754 8616 8760 8628
rect 7668 8588 8760 8616
rect 3326 8548 3332 8560
rect 1780 8520 3332 8548
rect 1780 8489 1808 8520
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 3694 8508 3700 8560
rect 3752 8508 3758 8560
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 7668 8548 7696 8588
rect 8754 8576 8760 8588
rect 8812 8616 8818 8628
rect 9490 8616 9496 8628
rect 8812 8588 9496 8616
rect 8812 8576 8818 8588
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10192 8588 10793 8616
rect 10192 8576 10198 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 10781 8579 10839 8585
rect 10873 8619 10931 8625
rect 10873 8585 10885 8619
rect 10919 8585 10931 8619
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 10873 8579 10931 8585
rect 11164 8588 11805 8616
rect 5776 8520 7696 8548
rect 5776 8508 5782 8520
rect 8478 8508 8484 8560
rect 8536 8508 8542 8560
rect 9030 8508 9036 8560
rect 9088 8548 9094 8560
rect 9585 8551 9643 8557
rect 9585 8548 9597 8551
rect 9088 8520 9597 8548
rect 9088 8508 9094 8520
rect 9585 8517 9597 8520
rect 9631 8517 9643 8551
rect 9585 8511 9643 8517
rect 10042 8508 10048 8560
rect 10100 8548 10106 8560
rect 10888 8548 10916 8579
rect 10100 8520 10916 8548
rect 10100 8508 10106 8520
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 2958 8440 2964 8492
rect 3016 8440 3022 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6086 8480 6092 8492
rect 5859 8452 6092 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6512 8452 6561 8480
rect 6512 8440 6518 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7466 8480 7472 8492
rect 6963 8452 7472 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 9306 8480 9312 8492
rect 9263 8452 9312 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9674 8440 9680 8492
rect 9732 8440 9738 8492
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 10318 8440 10324 8492
rect 10376 8480 10382 8492
rect 11164 8489 11192 8588
rect 11793 8585 11805 8588
rect 11839 8616 11851 8619
rect 11882 8616 11888 8628
rect 11839 8588 11888 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 13078 8576 13084 8628
rect 13136 8616 13142 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 13136 8588 13553 8616
rect 13136 8576 13142 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 21085 8619 21143 8625
rect 21085 8616 21097 8619
rect 20404 8588 21097 8616
rect 20404 8576 20410 8588
rect 21085 8585 21097 8588
rect 21131 8616 21143 8619
rect 22281 8619 22339 8625
rect 22281 8616 22293 8619
rect 21131 8588 22293 8616
rect 21131 8585 21143 8588
rect 21085 8579 21143 8585
rect 22281 8585 22293 8588
rect 22327 8585 22339 8619
rect 22281 8579 22339 8585
rect 22370 8576 22376 8628
rect 22428 8576 22434 8628
rect 22462 8576 22468 8628
rect 22520 8576 22526 8628
rect 22830 8576 22836 8628
rect 22888 8616 22894 8628
rect 23293 8619 23351 8625
rect 23293 8616 23305 8619
rect 22888 8588 23305 8616
rect 22888 8576 22894 8588
rect 23293 8585 23305 8588
rect 23339 8585 23351 8619
rect 23293 8579 23351 8585
rect 25130 8576 25136 8628
rect 25188 8576 25194 8628
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 25406 8616 25412 8628
rect 25280 8588 25412 8616
rect 25280 8576 25286 8588
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 26421 8619 26479 8625
rect 26421 8585 26433 8619
rect 26467 8616 26479 8619
rect 26786 8616 26792 8628
rect 26467 8588 26792 8616
rect 26467 8585 26479 8588
rect 26421 8579 26479 8585
rect 26786 8576 26792 8588
rect 26844 8576 26850 8628
rect 27154 8576 27160 8628
rect 27212 8616 27218 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 27212 8588 27353 8616
rect 27212 8576 27218 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 28810 8616 28816 8628
rect 27341 8579 27399 8585
rect 28644 8588 28816 8616
rect 11333 8551 11391 8557
rect 11333 8517 11345 8551
rect 11379 8548 11391 8551
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11379 8520 11713 8548
rect 11379 8517 11391 8520
rect 11333 8511 11391 8517
rect 11701 8517 11713 8520
rect 11747 8548 11759 8551
rect 12066 8548 12072 8560
rect 11747 8520 12072 8548
rect 11747 8517 11759 8520
rect 11701 8511 11759 8517
rect 12066 8508 12072 8520
rect 12124 8508 12130 8560
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 12342 8548 12348 8560
rect 12216 8520 12348 8548
rect 12216 8508 12222 8520
rect 12342 8508 12348 8520
rect 12400 8548 12406 8560
rect 12400 8520 12572 8548
rect 12400 8508 12406 8520
rect 10413 8483 10471 8489
rect 10413 8480 10425 8483
rect 10376 8452 10425 8480
rect 10376 8440 10382 8452
rect 10413 8449 10425 8452
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 1946 8412 1952 8424
rect 1903 8384 1952 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2866 8372 2872 8424
rect 2924 8372 2930 8424
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 2976 8384 3249 8412
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 2976 8344 3004 8384
rect 3237 8381 3249 8384
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 4856 8384 5917 8412
rect 4856 8372 4862 8384
rect 5905 8381 5917 8384
rect 5951 8381 5963 8415
rect 8386 8412 8392 8424
rect 5905 8375 5963 8381
rect 7484 8384 8392 8412
rect 7484 8353 7512 8384
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 8987 8384 9352 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9324 8353 9352 8384
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 10612 8412 10640 8443
rect 10336 8384 10640 8412
rect 11072 8412 11100 8443
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11296 8452 11897 8480
rect 11296 8440 11302 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 12084 8480 12112 8508
rect 12544 8489 12572 8520
rect 12986 8508 12992 8560
rect 13044 8508 13050 8560
rect 14550 8508 14556 8560
rect 14608 8508 14614 8560
rect 18138 8508 18144 8560
rect 18196 8508 18202 8560
rect 20162 8508 20168 8560
rect 20220 8508 20226 8560
rect 22097 8551 22155 8557
rect 22097 8517 22109 8551
rect 22143 8548 22155 8551
rect 25148 8548 25176 8576
rect 22143 8520 22968 8548
rect 25148 8520 25544 8548
rect 22143 8517 22155 8520
rect 22097 8511 22155 8517
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12084 8452 12449 8480
rect 11885 8443 11943 8449
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 22940 8489 22968 8520
rect 22925 8483 22983 8489
rect 22925 8449 22937 8483
rect 22971 8480 22983 8483
rect 23014 8480 23020 8492
rect 22971 8452 23020 8480
rect 22971 8449 22983 8452
rect 22925 8443 22983 8449
rect 23014 8440 23020 8452
rect 23072 8440 23078 8492
rect 25130 8440 25136 8492
rect 25188 8440 25194 8492
rect 25317 8483 25375 8489
rect 25317 8449 25329 8483
rect 25363 8449 25375 8483
rect 25317 8443 25375 8449
rect 11422 8412 11428 8424
rect 11072 8384 11428 8412
rect 10336 8353 10364 8384
rect 2179 8316 3004 8344
rect 7469 8347 7527 8353
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 7469 8313 7481 8347
rect 7515 8313 7527 8347
rect 7469 8307 7527 8313
rect 9309 8347 9367 8353
rect 9309 8313 9321 8347
rect 9355 8313 9367 8347
rect 9309 8307 9367 8313
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8313 10379 8347
rect 10612 8344 10640 8384
rect 11422 8372 11428 8384
rect 11480 8412 11486 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 11480 8384 12081 8412
rect 11480 8372 11486 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 11146 8344 11152 8356
rect 10612 8316 11152 8344
rect 10321 8307 10379 8313
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11388 8316 11529 8344
rect 11388 8304 11394 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 12084 8344 12112 8375
rect 12250 8372 12256 8424
rect 12308 8372 12314 8424
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8412 12403 8415
rect 13096 8412 13124 8440
rect 15013 8415 15071 8421
rect 15013 8412 15025 8415
rect 12391 8384 13124 8412
rect 13372 8384 15025 8412
rect 12391 8381 12403 8384
rect 12345 8375 12403 8381
rect 12360 8344 12388 8375
rect 12434 8344 12440 8356
rect 12084 8316 12440 8344
rect 11517 8307 11575 8313
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 13372 8353 13400 8384
rect 15013 8381 15025 8384
rect 15059 8381 15071 8415
rect 15013 8375 15071 8381
rect 15286 8372 15292 8424
rect 15344 8372 15350 8424
rect 18414 8372 18420 8424
rect 18472 8412 18478 8424
rect 18877 8415 18935 8421
rect 18877 8412 18889 8415
rect 18472 8384 18889 8412
rect 18472 8372 18478 8384
rect 18877 8381 18889 8384
rect 18923 8412 18935 8415
rect 19337 8415 19395 8421
rect 19337 8412 19349 8415
rect 18923 8384 19349 8412
rect 18923 8381 18935 8384
rect 18877 8375 18935 8381
rect 19337 8381 19349 8384
rect 19383 8381 19395 8415
rect 19337 8375 19395 8381
rect 19610 8372 19616 8424
rect 19668 8372 19674 8424
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 22278 8412 22284 8424
rect 20036 8384 22284 8412
rect 20036 8372 20042 8384
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 22738 8372 22744 8424
rect 22796 8412 22802 8424
rect 22833 8415 22891 8421
rect 22833 8412 22845 8415
rect 22796 8384 22845 8412
rect 22796 8372 22802 8384
rect 22833 8381 22845 8384
rect 22879 8381 22891 8415
rect 22833 8375 22891 8381
rect 24394 8372 24400 8424
rect 24452 8412 24458 8424
rect 25222 8412 25228 8424
rect 24452 8384 25228 8412
rect 24452 8372 24458 8384
rect 25222 8372 25228 8384
rect 25280 8372 25286 8424
rect 25332 8412 25360 8443
rect 25406 8440 25412 8492
rect 25464 8440 25470 8492
rect 25516 8489 25544 8520
rect 25501 8483 25559 8489
rect 25501 8449 25513 8483
rect 25547 8449 25559 8483
rect 26326 8480 26332 8492
rect 25501 8443 25559 8449
rect 25608 8452 26332 8480
rect 25608 8412 25636 8452
rect 26326 8440 26332 8452
rect 26384 8480 26390 8492
rect 26878 8480 26884 8492
rect 26384 8452 26884 8480
rect 26384 8440 26390 8452
rect 26878 8440 26884 8452
rect 26936 8440 26942 8492
rect 26970 8440 26976 8492
rect 27028 8440 27034 8492
rect 27154 8440 27160 8492
rect 27212 8440 27218 8492
rect 28644 8466 28672 8588
rect 28810 8576 28816 8588
rect 28868 8616 28874 8628
rect 29638 8616 29644 8628
rect 28868 8588 29644 8616
rect 28868 8576 28874 8588
rect 29638 8576 29644 8588
rect 29696 8576 29702 8628
rect 33042 8616 33048 8628
rect 32140 8588 33048 8616
rect 29730 8508 29736 8560
rect 29788 8508 29794 8560
rect 30009 8483 30067 8489
rect 30009 8449 30021 8483
rect 30055 8480 30067 8483
rect 31754 8480 31760 8492
rect 30055 8452 31760 8480
rect 30055 8449 30067 8452
rect 30009 8443 30067 8449
rect 31754 8440 31760 8452
rect 31812 8480 31818 8492
rect 32140 8489 32168 8588
rect 33042 8576 33048 8588
rect 33100 8576 33106 8628
rect 37093 8619 37151 8625
rect 34164 8588 35572 8616
rect 34164 8548 34192 8588
rect 33626 8520 34192 8548
rect 34238 8508 34244 8560
rect 34296 8508 34302 8560
rect 35544 8548 35572 8588
rect 37093 8585 37105 8619
rect 37139 8616 37151 8619
rect 38010 8616 38016 8628
rect 37139 8588 38016 8616
rect 37139 8585 37151 8588
rect 37093 8579 37151 8585
rect 38010 8576 38016 8588
rect 38068 8576 38074 8628
rect 38470 8576 38476 8628
rect 38528 8616 38534 8628
rect 38528 8588 38884 8616
rect 38528 8576 38534 8588
rect 36262 8548 36268 8560
rect 35466 8520 36268 8548
rect 36262 8508 36268 8520
rect 36320 8508 36326 8560
rect 38286 8508 38292 8560
rect 38344 8508 38350 8560
rect 38856 8557 38884 8588
rect 38841 8551 38899 8557
rect 38841 8517 38853 8551
rect 38887 8517 38899 8551
rect 38841 8511 38899 8517
rect 38930 8508 38936 8560
rect 38988 8548 38994 8560
rect 38988 8520 39160 8548
rect 38988 8508 38994 8520
rect 32125 8483 32183 8489
rect 32125 8480 32137 8483
rect 31812 8452 32137 8480
rect 31812 8440 31818 8452
rect 32125 8449 32137 8452
rect 32171 8449 32183 8483
rect 32125 8443 32183 8449
rect 35989 8483 36047 8489
rect 35989 8449 36001 8483
rect 36035 8480 36047 8483
rect 36078 8480 36084 8492
rect 36035 8452 36084 8480
rect 36035 8449 36047 8452
rect 35989 8443 36047 8449
rect 36078 8440 36084 8452
rect 36136 8440 36142 8492
rect 36173 8483 36231 8489
rect 36173 8449 36185 8483
rect 36219 8449 36231 8483
rect 36173 8443 36231 8449
rect 25332 8384 25636 8412
rect 25777 8415 25835 8421
rect 13357 8347 13415 8353
rect 13357 8313 13369 8347
rect 13403 8313 13415 8347
rect 22649 8347 22707 8353
rect 13357 8307 13415 8313
rect 20640 8316 22048 8344
rect 2222 8236 2228 8288
rect 2280 8236 2286 8288
rect 4706 8236 4712 8288
rect 4764 8236 4770 8288
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 5994 8276 6000 8288
rect 5408 8248 6000 8276
rect 5408 8236 5414 8248
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 6546 8236 6552 8288
rect 6604 8236 6610 8288
rect 11238 8236 11244 8288
rect 11296 8236 11302 8288
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 12802 8276 12808 8288
rect 12759 8248 12808 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 20640 8276 20668 8316
rect 19392 8248 20668 8276
rect 22020 8276 22048 8316
rect 22649 8313 22661 8347
rect 22695 8344 22707 8347
rect 24486 8344 24492 8356
rect 22695 8316 24492 8344
rect 22695 8313 22707 8316
rect 22649 8307 22707 8313
rect 24486 8304 24492 8316
rect 24544 8304 24550 8356
rect 25332 8344 25360 8384
rect 25777 8381 25789 8415
rect 25823 8381 25835 8415
rect 25777 8375 25835 8381
rect 28261 8415 28319 8421
rect 28261 8381 28273 8415
rect 28307 8412 28319 8415
rect 30653 8415 30711 8421
rect 30653 8412 30665 8415
rect 28307 8384 30665 8412
rect 28307 8381 28319 8384
rect 28261 8375 28319 8381
rect 30653 8381 30665 8384
rect 30699 8381 30711 8415
rect 30653 8375 30711 8381
rect 24780 8316 25360 8344
rect 25685 8347 25743 8353
rect 23750 8276 23756 8288
rect 22020 8248 23756 8276
rect 19392 8236 19398 8248
rect 23750 8236 23756 8248
rect 23808 8236 23814 8288
rect 24302 8236 24308 8288
rect 24360 8276 24366 8288
rect 24780 8276 24808 8316
rect 25685 8313 25697 8347
rect 25731 8344 25743 8347
rect 25792 8344 25820 8375
rect 32398 8372 32404 8424
rect 32456 8372 32462 8424
rect 33042 8372 33048 8424
rect 33100 8412 33106 8424
rect 33965 8415 34023 8421
rect 33965 8412 33977 8415
rect 33100 8384 33977 8412
rect 33100 8372 33106 8384
rect 33965 8381 33977 8384
rect 34011 8381 34023 8415
rect 34330 8412 34336 8424
rect 33965 8375 34023 8381
rect 34072 8384 34336 8412
rect 34072 8344 34100 8384
rect 34330 8372 34336 8384
rect 34388 8412 34394 8424
rect 35713 8415 35771 8421
rect 35713 8412 35725 8415
rect 34388 8384 35725 8412
rect 34388 8372 34394 8384
rect 35713 8381 35725 8384
rect 35759 8381 35771 8415
rect 36188 8412 36216 8443
rect 36538 8440 36544 8492
rect 36596 8480 36602 8492
rect 36725 8483 36783 8489
rect 36725 8480 36737 8483
rect 36596 8452 36737 8480
rect 36596 8440 36602 8452
rect 36725 8449 36737 8452
rect 36771 8449 36783 8483
rect 36725 8443 36783 8449
rect 36909 8483 36967 8489
rect 36909 8449 36921 8483
rect 36955 8480 36967 8483
rect 37090 8480 37096 8492
rect 36955 8452 37096 8480
rect 36955 8449 36967 8452
rect 36909 8443 36967 8449
rect 37090 8440 37096 8452
rect 37148 8480 37154 8492
rect 39132 8489 39160 8520
rect 39117 8483 39175 8489
rect 37148 8452 37412 8480
rect 37148 8440 37154 8452
rect 36998 8412 37004 8424
rect 36188 8384 37004 8412
rect 35713 8375 35771 8381
rect 36998 8372 37004 8384
rect 37056 8372 37062 8424
rect 37384 8356 37412 8452
rect 39117 8449 39129 8483
rect 39163 8449 39175 8483
rect 39117 8443 39175 8449
rect 37458 8372 37464 8424
rect 37516 8412 37522 8424
rect 39209 8415 39267 8421
rect 39209 8412 39221 8415
rect 37516 8384 39221 8412
rect 37516 8372 37522 8384
rect 39209 8381 39221 8384
rect 39255 8381 39267 8415
rect 39209 8375 39267 8381
rect 39758 8372 39764 8424
rect 39816 8372 39822 8424
rect 25731 8316 25820 8344
rect 33428 8316 34100 8344
rect 25731 8313 25743 8316
rect 25685 8307 25743 8313
rect 24360 8248 24808 8276
rect 24360 8236 24366 8248
rect 29730 8236 29736 8288
rect 29788 8276 29794 8288
rect 30098 8276 30104 8288
rect 29788 8248 30104 8276
rect 29788 8236 29794 8248
rect 30098 8236 30104 8248
rect 30156 8236 30162 8288
rect 32858 8236 32864 8288
rect 32916 8276 32922 8288
rect 33428 8276 33456 8316
rect 37366 8304 37372 8356
rect 37424 8304 37430 8356
rect 32916 8248 33456 8276
rect 32916 8236 32922 8248
rect 33870 8236 33876 8288
rect 33928 8236 33934 8288
rect 35986 8236 35992 8288
rect 36044 8236 36050 8288
rect 1104 8186 42504 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 42504 8186
rect 1104 8112 42504 8134
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 2924 8044 3157 8072
rect 2924 8032 2930 8044
rect 3145 8041 3157 8044
rect 3191 8072 3203 8075
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 3191 8044 3433 8072
rect 3191 8041 3203 8044
rect 3145 8035 3203 8041
rect 3421 8041 3433 8044
rect 3467 8072 3479 8075
rect 3878 8072 3884 8084
rect 3467 8044 3884 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8072 4123 8075
rect 4614 8072 4620 8084
rect 4111 8044 4620 8072
rect 4111 8041 4123 8044
rect 4065 8035 4123 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 8352 8044 8585 8072
rect 8352 8032 8358 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9493 8075 9551 8081
rect 8803 8044 9444 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 8588 7936 8616 8035
rect 9217 8007 9275 8013
rect 9217 7973 9229 8007
rect 9263 7973 9275 8007
rect 9217 7967 9275 7973
rect 8754 7936 8760 7948
rect 8588 7908 8760 7936
rect 8754 7896 8760 7908
rect 8812 7936 8818 7948
rect 8812 7908 9076 7936
rect 8812 7896 8818 7908
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 2958 7868 2964 7880
rect 2806 7840 2964 7868
rect 2958 7828 2964 7840
rect 3016 7868 3022 7880
rect 3694 7868 3700 7880
rect 3016 7840 3700 7868
rect 3016 7828 3022 7840
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7868 3847 7871
rect 3878 7868 3884 7880
rect 3835 7840 3884 7868
rect 3835 7837 3847 7840
rect 3789 7831 3847 7837
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4706 7868 4712 7880
rect 4203 7840 4712 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7800 1731 7803
rect 1762 7800 1768 7812
rect 1719 7772 1768 7800
rect 1719 7769 1731 7772
rect 1673 7763 1731 7769
rect 1762 7760 1768 7772
rect 1820 7760 1826 7812
rect 3389 7803 3447 7809
rect 3389 7800 3401 7803
rect 3068 7772 3401 7800
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 3068 7732 3096 7772
rect 3389 7769 3401 7772
rect 3435 7769 3447 7803
rect 3389 7763 3447 7769
rect 3602 7760 3608 7812
rect 3660 7800 3666 7812
rect 4172 7800 4200 7831
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 9048 7877 9076 7908
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9033 7871 9091 7877
rect 9033 7837 9045 7871
rect 9079 7837 9091 7871
rect 9232 7868 9260 7967
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 9232 7840 9321 7868
rect 9033 7831 9091 7837
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 9416 7868 9444 8044
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9674 8072 9680 8084
rect 9539 8044 9680 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10318 8032 10324 8084
rect 10376 8032 10382 8084
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 11790 8072 11796 8084
rect 11204 8044 11796 8072
rect 11204 8032 11210 8044
rect 11790 8032 11796 8044
rect 11848 8072 11854 8084
rect 12158 8072 12164 8084
rect 11848 8044 12164 8072
rect 11848 8032 11854 8044
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 19061 8075 19119 8081
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19610 8072 19616 8084
rect 19107 8044 19616 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 19794 8032 19800 8084
rect 19852 8072 19858 8084
rect 19889 8075 19947 8081
rect 19889 8072 19901 8075
rect 19852 8044 19901 8072
rect 19852 8032 19858 8044
rect 19889 8041 19901 8044
rect 19935 8041 19947 8075
rect 25409 8075 25467 8081
rect 25409 8072 25421 8075
rect 19889 8035 19947 8041
rect 24596 8044 25421 8072
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 11238 8004 11244 8016
rect 10008 7976 11244 8004
rect 10008 7964 10014 7976
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9416 7840 9505 7868
rect 9309 7831 9367 7837
rect 9493 7837 9505 7840
rect 9539 7868 9551 7871
rect 10134 7868 10140 7880
rect 9539 7840 10140 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 3660 7772 4200 7800
rect 3660 7760 3666 7772
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 8570 7760 8576 7812
rect 8628 7809 8634 7812
rect 8628 7803 8647 7809
rect 8635 7800 8647 7803
rect 8956 7800 8984 7831
rect 10134 7828 10140 7840
rect 10192 7868 10198 7880
rect 10520 7877 10548 7976
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 20346 8004 20352 8016
rect 18524 7976 20352 8004
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7936 10655 7939
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 10643 7908 11161 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 11882 7936 11888 7948
rect 11379 7908 11888 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 15286 7936 15292 7948
rect 13863 7908 15292 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 10192 7840 10333 7868
rect 10192 7828 10198 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11238 7868 11244 7880
rect 11103 7840 11244 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 11238 7828 11244 7840
rect 11296 7828 11302 7880
rect 11422 7828 11428 7880
rect 11480 7828 11486 7880
rect 11698 7828 11704 7880
rect 11756 7828 11762 7880
rect 11790 7828 11796 7880
rect 11848 7828 11854 7880
rect 18524 7877 18552 7976
rect 20346 7964 20352 7976
rect 20404 7964 20410 8016
rect 24118 7964 24124 8016
rect 24176 8004 24182 8016
rect 24596 8004 24624 8044
rect 25409 8041 25421 8044
rect 25455 8072 25467 8075
rect 26786 8072 26792 8084
rect 25455 8044 26792 8072
rect 25455 8041 25467 8044
rect 25409 8035 25467 8041
rect 26786 8032 26792 8044
rect 26844 8032 26850 8084
rect 26970 8032 26976 8084
rect 27028 8032 27034 8084
rect 29365 8075 29423 8081
rect 29365 8041 29377 8075
rect 29411 8072 29423 8075
rect 29822 8072 29828 8084
rect 29411 8044 29828 8072
rect 29411 8041 29423 8044
rect 29365 8035 29423 8041
rect 29822 8032 29828 8044
rect 29880 8032 29886 8084
rect 32125 8075 32183 8081
rect 32125 8041 32137 8075
rect 32171 8072 32183 8075
rect 32398 8072 32404 8084
rect 32171 8044 32404 8072
rect 32171 8041 32183 8044
rect 32125 8035 32183 8041
rect 32398 8032 32404 8044
rect 32456 8032 32462 8084
rect 33226 8032 33232 8084
rect 33284 8072 33290 8084
rect 33321 8075 33379 8081
rect 33321 8072 33333 8075
rect 33284 8044 33333 8072
rect 33284 8032 33290 8044
rect 33321 8041 33333 8044
rect 33367 8041 33379 8075
rect 33321 8035 33379 8041
rect 38654 8032 38660 8084
rect 38712 8072 38718 8084
rect 38749 8075 38807 8081
rect 38749 8072 38761 8075
rect 38712 8044 38761 8072
rect 38712 8032 38718 8044
rect 38749 8041 38761 8044
rect 38795 8041 38807 8075
rect 38749 8035 38807 8041
rect 24176 7976 24624 8004
rect 24176 7964 24182 7976
rect 19058 7896 19064 7948
rect 19116 7936 19122 7948
rect 19245 7939 19303 7945
rect 19245 7936 19257 7939
rect 19116 7908 19257 7936
rect 19116 7896 19122 7908
rect 19245 7905 19257 7908
rect 19291 7905 19303 7939
rect 19245 7899 19303 7905
rect 19702 7896 19708 7948
rect 19760 7936 19766 7948
rect 22186 7936 22192 7948
rect 19760 7908 20024 7936
rect 19760 7896 19766 7908
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19794 7868 19800 7880
rect 18923 7840 19800 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 19996 7877 20024 7908
rect 20272 7908 22192 7936
rect 20272 7877 20300 7908
rect 22186 7896 22192 7908
rect 22244 7936 22250 7948
rect 24394 7936 24400 7948
rect 22244 7908 24400 7936
rect 22244 7896 22250 7908
rect 24394 7896 24400 7908
rect 24452 7896 24458 7948
rect 24486 7896 24492 7948
rect 24544 7896 24550 7948
rect 19981 7871 20039 7877
rect 19981 7837 19993 7871
rect 20027 7837 20039 7871
rect 20257 7871 20315 7877
rect 20257 7868 20269 7871
rect 19981 7831 20039 7837
rect 20088 7840 20269 7868
rect 9217 7803 9275 7809
rect 9217 7800 9229 7803
rect 8635 7772 8984 7800
rect 9048 7772 9229 7800
rect 8635 7769 8647 7772
rect 8628 7763 8647 7769
rect 8628 7760 8634 7763
rect 2004 7704 3096 7732
rect 2004 7692 2010 7704
rect 3234 7692 3240 7744
rect 3292 7692 3298 7744
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 3881 7735 3939 7741
rect 3881 7732 3893 7735
rect 3844 7704 3893 7732
rect 3844 7692 3850 7704
rect 3881 7701 3893 7704
rect 3927 7701 3939 7735
rect 3881 7695 3939 7701
rect 3970 7692 3976 7744
rect 4028 7692 4034 7744
rect 8404 7732 8432 7760
rect 9048 7744 9076 7772
rect 9217 7769 9229 7772
rect 9263 7769 9275 7803
rect 9217 7763 9275 7769
rect 10965 7803 11023 7809
rect 10965 7769 10977 7803
rect 11011 7800 11023 7803
rect 11011 7772 12204 7800
rect 13110 7772 13492 7800
rect 11011 7769 11023 7772
rect 10965 7763 11023 7769
rect 9030 7732 9036 7744
rect 8404 7704 9036 7732
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 10870 7692 10876 7744
rect 10928 7692 10934 7744
rect 11609 7735 11667 7741
rect 11609 7701 11621 7735
rect 11655 7732 11667 7735
rect 12066 7732 12072 7744
rect 11655 7704 12072 7732
rect 11655 7701 11667 7704
rect 11609 7695 11667 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 12176 7732 12204 7772
rect 12802 7732 12808 7744
rect 12176 7704 12808 7732
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 13464 7732 13492 7772
rect 13538 7760 13544 7812
rect 13596 7760 13602 7812
rect 18690 7760 18696 7812
rect 18748 7760 18754 7812
rect 18785 7803 18843 7809
rect 18785 7769 18797 7803
rect 18831 7800 18843 7803
rect 20088 7800 20116 7840
rect 20257 7837 20269 7840
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7868 20959 7871
rect 22922 7868 22928 7880
rect 20947 7840 22928 7868
rect 20947 7837 20959 7840
rect 20901 7831 20959 7837
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 18831 7772 20116 7800
rect 18831 7769 18843 7772
rect 18785 7763 18843 7769
rect 20162 7760 20168 7812
rect 20220 7760 20226 7812
rect 24504 7800 24532 7896
rect 24596 7877 24624 7976
rect 25593 8007 25651 8013
rect 25593 7973 25605 8007
rect 25639 8004 25651 8007
rect 27154 8004 27160 8016
rect 25639 7976 27160 8004
rect 25639 7973 25651 7976
rect 25593 7967 25651 7973
rect 27154 7964 27160 7976
rect 27212 8004 27218 8016
rect 31662 8004 31668 8016
rect 27212 7976 27292 8004
rect 27212 7964 27218 7976
rect 25130 7896 25136 7948
rect 25188 7936 25194 7948
rect 25188 7908 27016 7936
rect 25188 7896 25194 7908
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 25240 7809 25268 7908
rect 25314 7828 25320 7880
rect 25372 7868 25378 7880
rect 25685 7871 25743 7877
rect 25685 7868 25697 7871
rect 25372 7840 25697 7868
rect 25372 7828 25378 7840
rect 25685 7837 25697 7840
rect 25731 7837 25743 7871
rect 26697 7871 26755 7877
rect 26697 7868 26709 7871
rect 25685 7831 25743 7837
rect 25792 7840 26709 7868
rect 25225 7803 25283 7809
rect 20272 7772 20760 7800
rect 24504 7772 25084 7800
rect 14550 7732 14556 7744
rect 13464 7704 14556 7732
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 20272 7732 20300 7772
rect 18104 7704 20300 7732
rect 18104 7692 18110 7704
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 20732 7741 20760 7772
rect 20717 7735 20775 7741
rect 20717 7701 20729 7735
rect 20763 7732 20775 7735
rect 21266 7732 21272 7744
rect 20763 7704 21272 7732
rect 20763 7701 20775 7704
rect 20717 7695 20775 7701
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 24946 7692 24952 7744
rect 25004 7692 25010 7744
rect 25056 7732 25084 7772
rect 25225 7769 25237 7803
rect 25271 7769 25283 7803
rect 25792 7800 25820 7840
rect 26697 7837 26709 7840
rect 26743 7837 26755 7871
rect 26697 7831 26755 7837
rect 26786 7828 26792 7880
rect 26844 7828 26850 7880
rect 26988 7877 27016 7908
rect 27264 7877 27292 7976
rect 31312 7976 31668 8004
rect 29086 7896 29092 7948
rect 29144 7896 29150 7948
rect 31312 7880 31340 7976
rect 31662 7964 31668 7976
rect 31720 7964 31726 8016
rect 32033 8007 32091 8013
rect 32033 7973 32045 8007
rect 32079 7973 32091 8007
rect 32033 7967 32091 7973
rect 31570 7896 31576 7948
rect 31628 7896 31634 7948
rect 32048 7936 32076 7967
rect 32214 7936 32220 7948
rect 32048 7908 32220 7936
rect 32214 7896 32220 7908
rect 32272 7936 32278 7948
rect 32677 7939 32735 7945
rect 32272 7908 32444 7936
rect 32272 7896 32278 7908
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7837 27307 7871
rect 27249 7831 27307 7837
rect 28997 7871 29055 7877
rect 28997 7837 29009 7871
rect 29043 7868 29055 7871
rect 29043 7840 29500 7868
rect 29043 7837 29055 7840
rect 28997 7831 29055 7837
rect 25225 7763 25283 7769
rect 25516 7772 25820 7800
rect 25425 7735 25483 7741
rect 25425 7732 25437 7735
rect 25056 7704 25437 7732
rect 25425 7701 25437 7704
rect 25471 7732 25483 7735
rect 25516 7732 25544 7772
rect 26234 7760 26240 7812
rect 26292 7800 26298 7812
rect 26418 7800 26424 7812
rect 26292 7772 26424 7800
rect 26292 7760 26298 7772
rect 26418 7760 26424 7772
rect 26476 7760 26482 7812
rect 27080 7800 27108 7831
rect 27430 7800 27436 7812
rect 27080 7772 27436 7800
rect 27430 7760 27436 7772
rect 27488 7760 27494 7812
rect 29472 7744 29500 7840
rect 31294 7828 31300 7880
rect 31352 7828 31358 7880
rect 31665 7871 31723 7877
rect 31665 7837 31677 7871
rect 31711 7837 31723 7871
rect 31665 7831 31723 7837
rect 29638 7760 29644 7812
rect 29696 7800 29702 7812
rect 29696 7772 29854 7800
rect 29696 7760 29702 7772
rect 31018 7760 31024 7812
rect 31076 7760 31082 7812
rect 31680 7800 31708 7831
rect 32122 7828 32128 7880
rect 32180 7868 32186 7880
rect 32416 7877 32444 7908
rect 32677 7905 32689 7939
rect 32723 7936 32735 7939
rect 33244 7936 33272 8032
rect 37369 8007 37427 8013
rect 37369 7973 37381 8007
rect 37415 8004 37427 8007
rect 39758 8004 39764 8016
rect 37415 7976 39764 8004
rect 37415 7973 37427 7976
rect 37369 7967 37427 7973
rect 39758 7964 39764 7976
rect 39816 7964 39822 8016
rect 32723 7908 33272 7936
rect 32723 7905 32735 7908
rect 32677 7899 32735 7905
rect 33870 7896 33876 7948
rect 33928 7896 33934 7948
rect 35342 7896 35348 7948
rect 35400 7936 35406 7948
rect 35621 7939 35679 7945
rect 35621 7936 35633 7939
rect 35400 7908 35633 7936
rect 35400 7896 35406 7908
rect 35621 7905 35633 7908
rect 35667 7936 35679 7939
rect 38930 7936 38936 7948
rect 35667 7908 38936 7936
rect 35667 7905 35679 7908
rect 35621 7899 35679 7905
rect 32309 7871 32367 7877
rect 32309 7868 32321 7871
rect 32180 7840 32321 7868
rect 32180 7828 32186 7840
rect 32309 7837 32321 7840
rect 32355 7837 32367 7871
rect 32309 7831 32367 7837
rect 32401 7871 32459 7877
rect 32401 7837 32413 7871
rect 32447 7837 32459 7871
rect 32858 7868 32864 7880
rect 32401 7831 32459 7837
rect 32692 7840 32864 7868
rect 32692 7800 32720 7840
rect 32858 7828 32864 7840
rect 32916 7828 32922 7880
rect 38396 7877 38424 7908
rect 38930 7896 38936 7908
rect 38988 7896 38994 7948
rect 38381 7871 38439 7877
rect 38381 7837 38393 7871
rect 38427 7837 38439 7871
rect 38381 7831 38439 7837
rect 38654 7828 38660 7880
rect 38712 7828 38718 7880
rect 38841 7871 38899 7877
rect 38841 7837 38853 7871
rect 38887 7837 38899 7871
rect 38841 7831 38899 7837
rect 31680 7772 32720 7800
rect 32766 7760 32772 7812
rect 32824 7800 32830 7812
rect 35158 7800 35164 7812
rect 32824 7772 35164 7800
rect 32824 7760 32830 7772
rect 35158 7760 35164 7772
rect 35216 7760 35222 7812
rect 35894 7760 35900 7812
rect 35952 7760 35958 7812
rect 36354 7760 36360 7812
rect 36412 7760 36418 7812
rect 37366 7760 37372 7812
rect 37424 7800 37430 7812
rect 38856 7800 38884 7831
rect 37424 7772 38884 7800
rect 37424 7760 37430 7772
rect 25471 7704 25544 7732
rect 27157 7735 27215 7741
rect 25471 7701 25483 7704
rect 25425 7695 25483 7701
rect 27157 7701 27169 7735
rect 27203 7732 27215 7735
rect 28166 7732 28172 7744
rect 27203 7704 28172 7732
rect 27203 7701 27215 7704
rect 27157 7695 27215 7701
rect 28166 7692 28172 7704
rect 28224 7692 28230 7744
rect 29454 7692 29460 7744
rect 29512 7732 29518 7744
rect 29549 7735 29607 7741
rect 29549 7732 29561 7735
rect 29512 7704 29561 7732
rect 29512 7692 29518 7704
rect 29549 7701 29561 7704
rect 29595 7701 29607 7735
rect 29549 7695 29607 7701
rect 32122 7692 32128 7744
rect 32180 7732 32186 7744
rect 34882 7732 34888 7744
rect 32180 7704 34888 7732
rect 32180 7692 32186 7704
rect 34882 7692 34888 7704
rect 34940 7732 34946 7744
rect 36170 7732 36176 7744
rect 34940 7704 36176 7732
rect 34940 7692 34946 7704
rect 36170 7692 36176 7704
rect 36228 7692 36234 7744
rect 1104 7642 42504 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 42504 7642
rect 1104 7568 42504 7590
rect 1762 7488 1768 7540
rect 1820 7488 1826 7540
rect 2866 7528 2872 7540
rect 1872 7500 2872 7528
rect 1872 7460 1900 7500
rect 2866 7488 2872 7500
rect 2924 7528 2930 7540
rect 3234 7528 3240 7540
rect 2924 7500 3240 7528
rect 2924 7488 2930 7500
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11296 7500 11529 7528
rect 11296 7488 11302 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 12434 7488 12440 7540
rect 12492 7488 12498 7540
rect 12989 7531 13047 7537
rect 12989 7497 13001 7531
rect 13035 7528 13047 7531
rect 13538 7528 13544 7540
rect 13035 7500 13544 7528
rect 13035 7497 13047 7500
rect 12989 7491 13047 7497
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 18690 7488 18696 7540
rect 18748 7528 18754 7540
rect 20162 7528 20168 7540
rect 18748 7500 20168 7528
rect 18748 7488 18754 7500
rect 20162 7488 20168 7500
rect 20220 7528 20226 7540
rect 22278 7528 22284 7540
rect 20220 7500 22284 7528
rect 20220 7488 20226 7500
rect 22278 7488 22284 7500
rect 22336 7528 22342 7540
rect 22336 7500 23704 7528
rect 22336 7488 22342 7500
rect 1688 7432 1900 7460
rect 1688 7401 1716 7432
rect 2222 7420 2228 7472
rect 2280 7420 2286 7472
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12621 7463 12679 7469
rect 12621 7460 12633 7463
rect 12124 7432 12633 7460
rect 12124 7420 12130 7432
rect 12621 7429 12633 7432
rect 12667 7460 12679 7463
rect 12667 7432 13124 7460
rect 12667 7429 12679 7432
rect 12621 7423 12679 7429
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 1872 7324 1900 7355
rect 1946 7352 1952 7404
rect 2004 7352 2010 7404
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 3602 7392 3608 7404
rect 2087 7364 3608 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11664 7364 11713 7392
rect 11664 7352 11670 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 12158 7352 12164 7404
rect 12216 7392 12222 7404
rect 12345 7395 12403 7401
rect 12345 7392 12357 7395
rect 12216 7364 12357 7392
rect 12216 7352 12222 7364
rect 12345 7361 12357 7364
rect 12391 7361 12403 7395
rect 12345 7355 12403 7361
rect 12713 7395 12771 7401
rect 12713 7361 12725 7395
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 1872 7296 2268 7324
rect 2240 7265 2268 7296
rect 11882 7284 11888 7336
rect 11940 7284 11946 7336
rect 12728 7324 12756 7355
rect 12802 7352 12808 7404
rect 12860 7352 12866 7404
rect 13096 7401 13124 7432
rect 13170 7420 13176 7472
rect 13228 7460 13234 7472
rect 19610 7460 19616 7472
rect 13228 7432 13308 7460
rect 13228 7420 13234 7432
rect 13280 7401 13308 7432
rect 19260 7432 19616 7460
rect 19260 7401 19288 7432
rect 19610 7420 19616 7432
rect 19668 7420 19674 7472
rect 19705 7463 19763 7469
rect 19705 7429 19717 7463
rect 19751 7460 19763 7463
rect 20346 7460 20352 7472
rect 19751 7432 20352 7460
rect 19751 7429 19763 7432
rect 19705 7423 19763 7429
rect 20346 7420 20352 7432
rect 20404 7460 20410 7472
rect 20717 7463 20775 7469
rect 20717 7460 20729 7463
rect 20404 7432 20729 7460
rect 20404 7420 20410 7432
rect 20717 7429 20729 7432
rect 20763 7429 20775 7463
rect 20717 7423 20775 7429
rect 21266 7420 21272 7472
rect 21324 7420 21330 7472
rect 23198 7460 23204 7472
rect 22862 7432 23204 7460
rect 23198 7420 23204 7432
rect 23256 7460 23262 7472
rect 23382 7460 23388 7472
rect 23256 7432 23388 7460
rect 23256 7420 23262 7432
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 23676 7460 23704 7500
rect 23750 7488 23756 7540
rect 23808 7528 23814 7540
rect 23808 7500 24808 7528
rect 23808 7488 23814 7500
rect 24780 7472 24808 7500
rect 27338 7488 27344 7540
rect 27396 7528 27402 7540
rect 28537 7531 28595 7537
rect 28537 7528 28549 7531
rect 27396 7500 28549 7528
rect 27396 7488 27402 7500
rect 28537 7497 28549 7500
rect 28583 7497 28595 7531
rect 30466 7528 30472 7540
rect 28537 7491 28595 7497
rect 29012 7500 30472 7528
rect 24302 7460 24308 7472
rect 23676 7432 24308 7460
rect 24302 7420 24308 7432
rect 24360 7420 24366 7472
rect 24394 7420 24400 7472
rect 24452 7420 24458 7472
rect 24762 7420 24768 7472
rect 24820 7460 24826 7472
rect 24820 7432 26188 7460
rect 24820 7420 24826 7432
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 19245 7395 19303 7401
rect 19245 7361 19257 7395
rect 19291 7361 19303 7395
rect 19245 7355 19303 7361
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 24486 7352 24492 7404
rect 24544 7392 24550 7404
rect 25501 7395 25559 7401
rect 25501 7392 25513 7395
rect 24544 7364 25513 7392
rect 24544 7352 24550 7364
rect 25501 7361 25513 7364
rect 25547 7361 25559 7395
rect 25501 7355 25559 7361
rect 12636 7296 12756 7324
rect 12989 7327 13047 7333
rect 12636 7265 12664 7296
rect 12989 7293 13001 7327
rect 13035 7324 13047 7327
rect 13173 7327 13231 7333
rect 13173 7324 13185 7327
rect 13035 7296 13185 7324
rect 13035 7293 13047 7296
rect 12989 7287 13047 7293
rect 13173 7293 13185 7296
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 19613 7327 19671 7333
rect 19613 7293 19625 7327
rect 19659 7324 19671 7327
rect 19978 7324 19984 7336
rect 19659 7296 19984 7324
rect 19659 7293 19671 7296
rect 19613 7287 19671 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20162 7284 20168 7336
rect 20220 7284 20226 7336
rect 23290 7284 23296 7336
rect 23348 7284 23354 7336
rect 23566 7284 23572 7336
rect 23624 7284 23630 7336
rect 24765 7327 24823 7333
rect 24765 7293 24777 7327
rect 24811 7293 24823 7327
rect 24765 7287 24823 7293
rect 2225 7259 2283 7265
rect 2225 7225 2237 7259
rect 2271 7225 2283 7259
rect 2225 7219 2283 7225
rect 12621 7259 12679 7265
rect 12621 7225 12633 7259
rect 12667 7225 12679 7259
rect 12621 7219 12679 7225
rect 14550 7216 14556 7268
rect 14608 7256 14614 7268
rect 20806 7256 20812 7268
rect 14608 7228 20812 7256
rect 14608 7216 14614 7228
rect 20806 7216 20812 7228
rect 20864 7256 20870 7268
rect 20993 7259 21051 7265
rect 20993 7256 21005 7259
rect 20864 7228 21005 7256
rect 20864 7216 20870 7228
rect 20993 7225 21005 7228
rect 21039 7225 21051 7259
rect 20993 7219 21051 7225
rect 24673 7259 24731 7265
rect 24673 7225 24685 7259
rect 24719 7256 24731 7259
rect 24780 7256 24808 7287
rect 26050 7284 26056 7336
rect 26108 7284 26114 7336
rect 26160 7324 26188 7432
rect 27154 7420 27160 7472
rect 27212 7460 27218 7472
rect 27212 7432 27936 7460
rect 27212 7420 27218 7432
rect 26234 7352 26240 7404
rect 26292 7352 26298 7404
rect 27249 7395 27307 7401
rect 27249 7361 27261 7395
rect 27295 7392 27307 7395
rect 27338 7392 27344 7404
rect 27295 7364 27344 7392
rect 27295 7361 27307 7364
rect 27249 7355 27307 7361
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 27525 7395 27583 7401
rect 27525 7361 27537 7395
rect 27571 7392 27583 7395
rect 27798 7392 27804 7404
rect 27571 7364 27804 7392
rect 27571 7361 27583 7364
rect 27525 7355 27583 7361
rect 27798 7352 27804 7364
rect 27856 7352 27862 7404
rect 27908 7401 27936 7432
rect 28166 7420 28172 7472
rect 28224 7420 28230 7472
rect 29012 7460 29040 7500
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 30653 7531 30711 7537
rect 30653 7497 30665 7531
rect 30699 7528 30711 7531
rect 31018 7528 31024 7540
rect 30699 7500 31024 7528
rect 30699 7497 30711 7500
rect 30653 7491 30711 7497
rect 31018 7488 31024 7500
rect 31076 7488 31082 7540
rect 32398 7488 32404 7540
rect 32456 7528 32462 7540
rect 32493 7531 32551 7537
rect 32493 7528 32505 7531
rect 32456 7500 32505 7528
rect 32456 7488 32462 7500
rect 32493 7497 32505 7500
rect 32539 7528 32551 7531
rect 32674 7528 32680 7540
rect 32539 7500 32680 7528
rect 32539 7497 32551 7500
rect 32493 7491 32551 7497
rect 32674 7488 32680 7500
rect 32732 7488 32738 7540
rect 34441 7531 34499 7537
rect 34441 7528 34453 7531
rect 33888 7500 34453 7528
rect 28368 7432 29040 7460
rect 28368 7401 28396 7432
rect 29086 7420 29092 7472
rect 29144 7460 29150 7472
rect 30837 7463 30895 7469
rect 30837 7460 30849 7463
rect 29144 7432 30849 7460
rect 29144 7420 29150 7432
rect 30837 7429 30849 7432
rect 30883 7429 30895 7463
rect 31386 7460 31392 7472
rect 30837 7423 30895 7429
rect 30944 7432 31392 7460
rect 30944 7404 30972 7432
rect 31386 7420 31392 7432
rect 31444 7420 31450 7472
rect 31570 7420 31576 7472
rect 31628 7460 31634 7472
rect 33888 7460 33916 7500
rect 34441 7497 34453 7500
rect 34487 7497 34499 7531
rect 34441 7491 34499 7497
rect 34698 7488 34704 7540
rect 34756 7488 34762 7540
rect 34974 7488 34980 7540
rect 35032 7528 35038 7540
rect 35434 7528 35440 7540
rect 35032 7500 35440 7528
rect 35032 7488 35038 7500
rect 35434 7488 35440 7500
rect 35492 7528 35498 7540
rect 35805 7531 35863 7537
rect 35805 7528 35817 7531
rect 35492 7500 35817 7528
rect 35492 7488 35498 7500
rect 35805 7497 35817 7500
rect 35851 7497 35863 7531
rect 37642 7528 37648 7540
rect 35805 7491 35863 7497
rect 37476 7500 37648 7528
rect 31628 7432 33916 7460
rect 31628 7420 31634 7432
rect 27893 7395 27951 7401
rect 27893 7361 27905 7395
rect 27939 7361 27951 7395
rect 27893 7355 27951 7361
rect 28077 7395 28135 7401
rect 28077 7361 28089 7395
rect 28123 7392 28135 7395
rect 28353 7395 28411 7401
rect 28353 7392 28365 7395
rect 28123 7364 28365 7392
rect 28123 7361 28135 7364
rect 28077 7355 28135 7361
rect 28353 7361 28365 7364
rect 28399 7361 28411 7395
rect 28353 7355 28411 7361
rect 29365 7395 29423 7401
rect 29365 7361 29377 7395
rect 29411 7392 29423 7395
rect 29454 7392 29460 7404
rect 29411 7364 29460 7392
rect 29411 7361 29423 7364
rect 29365 7355 29423 7361
rect 27157 7327 27215 7333
rect 27157 7324 27169 7327
rect 26160 7296 27169 7324
rect 27157 7293 27169 7296
rect 27203 7293 27215 7327
rect 27157 7287 27215 7293
rect 24719 7228 24808 7256
rect 24719 7225 24731 7228
rect 24673 7219 24731 7225
rect 18690 7148 18696 7200
rect 18748 7188 18754 7200
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 18748 7160 19073 7188
rect 18748 7148 18754 7160
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 21818 7148 21824 7200
rect 21876 7148 21882 7200
rect 25406 7148 25412 7200
rect 25464 7148 25470 7200
rect 26970 7148 26976 7200
rect 27028 7148 27034 7200
rect 27172 7188 27200 7287
rect 27614 7284 27620 7336
rect 27672 7284 27678 7336
rect 27709 7327 27767 7333
rect 27709 7293 27721 7327
rect 27755 7324 27767 7327
rect 28902 7324 28908 7336
rect 27755 7296 28908 7324
rect 27755 7293 27767 7296
rect 27709 7287 27767 7293
rect 27430 7216 27436 7268
rect 27488 7256 27494 7268
rect 27724 7256 27752 7287
rect 28902 7284 28908 7296
rect 28960 7284 28966 7336
rect 29270 7284 29276 7336
rect 29328 7284 29334 7336
rect 27488 7228 27752 7256
rect 27488 7216 27494 7228
rect 28442 7216 28448 7268
rect 28500 7256 28506 7268
rect 28629 7259 28687 7265
rect 28629 7256 28641 7259
rect 28500 7228 28641 7256
rect 28500 7216 28506 7228
rect 28629 7225 28641 7228
rect 28675 7225 28687 7259
rect 28629 7219 28687 7225
rect 29086 7188 29092 7200
rect 27172 7160 29092 7188
rect 29086 7148 29092 7160
rect 29144 7148 29150 7200
rect 29380 7188 29408 7355
rect 29454 7352 29460 7364
rect 29512 7352 29518 7404
rect 29549 7395 29607 7401
rect 29549 7361 29561 7395
rect 29595 7361 29607 7395
rect 29549 7355 29607 7361
rect 29564 7324 29592 7355
rect 29638 7352 29644 7404
rect 29696 7352 29702 7404
rect 29730 7352 29736 7404
rect 29788 7352 29794 7404
rect 30650 7392 30656 7404
rect 29932 7364 30656 7392
rect 29932 7324 29960 7364
rect 30650 7352 30656 7364
rect 30708 7352 30714 7404
rect 30745 7395 30803 7401
rect 30745 7361 30757 7395
rect 30791 7392 30803 7395
rect 30791 7364 30880 7392
rect 30791 7361 30803 7364
rect 30745 7355 30803 7361
rect 29564 7296 29960 7324
rect 30009 7327 30067 7333
rect 30009 7293 30021 7327
rect 30055 7293 30067 7327
rect 30009 7287 30067 7293
rect 29917 7259 29975 7265
rect 29917 7225 29929 7259
rect 29963 7256 29975 7259
rect 30024 7256 30052 7287
rect 29963 7228 30052 7256
rect 30852 7256 30880 7364
rect 30926 7352 30932 7404
rect 30984 7352 30990 7404
rect 31113 7395 31171 7401
rect 31113 7361 31125 7395
rect 31159 7392 31171 7395
rect 31754 7392 31760 7404
rect 31159 7364 31760 7392
rect 31159 7361 31171 7364
rect 31113 7355 31171 7361
rect 31754 7352 31760 7364
rect 31812 7352 31818 7404
rect 32140 7401 32168 7432
rect 33888 7401 33916 7432
rect 34241 7463 34299 7469
rect 34241 7429 34253 7463
rect 34287 7429 34299 7463
rect 34241 7423 34299 7429
rect 32125 7395 32183 7401
rect 32125 7361 32137 7395
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 32218 7395 32276 7401
rect 32218 7361 32230 7395
rect 32264 7361 32276 7395
rect 32218 7355 32276 7361
rect 33873 7395 33931 7401
rect 33873 7361 33885 7395
rect 33919 7361 33931 7395
rect 33873 7355 33931 7361
rect 33965 7395 34023 7401
rect 33965 7361 33977 7395
rect 34011 7361 34023 7395
rect 33965 7355 34023 7361
rect 31018 7284 31024 7336
rect 31076 7324 31082 7336
rect 31205 7327 31263 7333
rect 31205 7324 31217 7327
rect 31076 7296 31217 7324
rect 31076 7284 31082 7296
rect 31205 7293 31217 7296
rect 31251 7293 31263 7327
rect 31205 7287 31263 7293
rect 31294 7284 31300 7336
rect 31352 7284 31358 7336
rect 31386 7284 31392 7336
rect 31444 7284 31450 7336
rect 31573 7327 31631 7333
rect 31573 7293 31585 7327
rect 31619 7324 31631 7327
rect 32232 7324 32260 7355
rect 31619 7296 32260 7324
rect 33980 7324 34008 7355
rect 34146 7352 34152 7404
rect 34204 7392 34210 7404
rect 34256 7392 34284 7423
rect 34790 7420 34796 7472
rect 34848 7460 34854 7472
rect 35253 7463 35311 7469
rect 35253 7460 35265 7463
rect 34848 7432 35265 7460
rect 34848 7420 34854 7432
rect 35253 7429 35265 7432
rect 35299 7429 35311 7463
rect 35253 7423 35311 7429
rect 35360 7432 35940 7460
rect 34204 7364 34284 7392
rect 34204 7352 34210 7364
rect 34882 7352 34888 7404
rect 34940 7352 34946 7404
rect 34974 7352 34980 7404
rect 35032 7352 35038 7404
rect 35158 7352 35164 7404
rect 35216 7392 35222 7404
rect 35360 7401 35388 7432
rect 35345 7395 35403 7401
rect 35345 7392 35357 7395
rect 35216 7364 35357 7392
rect 35216 7352 35222 7364
rect 35345 7361 35357 7364
rect 35391 7361 35403 7395
rect 35345 7355 35403 7361
rect 35437 7395 35495 7401
rect 35437 7361 35449 7395
rect 35483 7392 35495 7395
rect 35621 7395 35679 7401
rect 35483 7364 35572 7392
rect 35483 7361 35495 7364
rect 35437 7355 35495 7361
rect 34330 7324 34336 7336
rect 33980 7296 34336 7324
rect 31619 7293 31631 7296
rect 31573 7287 31631 7293
rect 34330 7284 34336 7296
rect 34388 7284 34394 7336
rect 31312 7256 31340 7284
rect 30852 7228 31340 7256
rect 34149 7259 34207 7265
rect 29963 7225 29975 7228
rect 29917 7219 29975 7225
rect 34149 7225 34161 7259
rect 34195 7256 34207 7259
rect 35544 7256 35572 7364
rect 35621 7361 35633 7395
rect 35667 7361 35679 7395
rect 35912 7392 35940 7432
rect 35986 7420 35992 7472
rect 36044 7420 36050 7472
rect 36173 7463 36231 7469
rect 36173 7429 36185 7463
rect 36219 7460 36231 7463
rect 36538 7460 36544 7472
rect 36219 7432 36544 7460
rect 36219 7429 36231 7432
rect 36173 7423 36231 7429
rect 36538 7420 36544 7432
rect 36596 7460 36602 7472
rect 37476 7469 37504 7500
rect 37642 7488 37648 7500
rect 37700 7528 37706 7540
rect 38930 7528 38936 7540
rect 37700 7500 38936 7528
rect 37700 7488 37706 7500
rect 38930 7488 38936 7500
rect 38988 7488 38994 7540
rect 41414 7528 41420 7540
rect 41386 7488 41420 7528
rect 41472 7488 41478 7540
rect 37461 7463 37519 7469
rect 36596 7432 37412 7460
rect 36596 7420 36602 7432
rect 36354 7392 36360 7404
rect 35912 7364 36360 7392
rect 35621 7355 35679 7361
rect 34195 7228 35572 7256
rect 35636 7256 35664 7355
rect 36354 7352 36360 7364
rect 36412 7352 36418 7404
rect 36446 7352 36452 7404
rect 36504 7352 36510 7404
rect 36633 7395 36691 7401
rect 36633 7361 36645 7395
rect 36679 7361 36691 7395
rect 36633 7355 36691 7361
rect 36538 7284 36544 7336
rect 36596 7324 36602 7336
rect 36648 7324 36676 7355
rect 36722 7352 36728 7404
rect 36780 7352 36786 7404
rect 36814 7352 36820 7404
rect 36872 7352 36878 7404
rect 37182 7392 37188 7404
rect 36924 7364 37188 7392
rect 36924 7324 36952 7364
rect 37182 7352 37188 7364
rect 37240 7352 37246 7404
rect 37384 7392 37412 7432
rect 37461 7429 37473 7463
rect 37507 7429 37519 7463
rect 37461 7423 37519 7429
rect 38194 7420 38200 7472
rect 38252 7420 38258 7472
rect 38654 7460 38660 7472
rect 38396 7432 38660 7460
rect 38396 7392 38424 7432
rect 38654 7420 38660 7432
rect 38712 7420 38718 7472
rect 37384 7364 38424 7392
rect 38473 7395 38531 7401
rect 38473 7361 38485 7395
rect 38519 7361 38531 7395
rect 38473 7355 38531 7361
rect 36596 7296 36952 7324
rect 36596 7284 36602 7296
rect 36998 7284 37004 7336
rect 37056 7324 37062 7336
rect 38289 7327 38347 7333
rect 38289 7324 38301 7327
rect 37056 7296 38301 7324
rect 37056 7284 37062 7296
rect 38289 7293 38301 7296
rect 38335 7293 38347 7327
rect 38289 7287 38347 7293
rect 36078 7256 36084 7268
rect 35636 7228 36084 7256
rect 34195 7225 34207 7228
rect 34149 7219 34207 7225
rect 31018 7188 31024 7200
rect 29380 7160 31024 7188
rect 31018 7148 31024 7160
rect 31076 7148 31082 7200
rect 34330 7148 34336 7200
rect 34388 7188 34394 7200
rect 34425 7191 34483 7197
rect 34425 7188 34437 7191
rect 34388 7160 34437 7188
rect 34388 7148 34394 7160
rect 34425 7157 34437 7160
rect 34471 7157 34483 7191
rect 34425 7151 34483 7157
rect 34609 7191 34667 7197
rect 34609 7157 34621 7191
rect 34655 7188 34667 7191
rect 35636 7188 35664 7228
rect 36078 7216 36084 7228
rect 36136 7256 36142 7268
rect 38488 7256 38516 7355
rect 38746 7352 38752 7404
rect 38804 7392 38810 7404
rect 39666 7392 39672 7404
rect 38804 7364 39672 7392
rect 38804 7352 38810 7364
rect 39666 7352 39672 7364
rect 39724 7352 39730 7404
rect 36136 7228 38516 7256
rect 36136 7216 36142 7228
rect 38838 7216 38844 7268
rect 38896 7256 38902 7268
rect 38933 7259 38991 7265
rect 38933 7256 38945 7259
rect 38896 7228 38945 7256
rect 38896 7216 38902 7228
rect 38933 7225 38945 7228
rect 38979 7256 38991 7259
rect 41386 7256 41414 7488
rect 38979 7228 41414 7256
rect 38979 7225 38991 7228
rect 38933 7219 38991 7225
rect 34655 7160 35664 7188
rect 34655 7157 34667 7160
rect 34609 7151 34667 7157
rect 35986 7148 35992 7200
rect 36044 7188 36050 7200
rect 36357 7191 36415 7197
rect 36357 7188 36369 7191
rect 36044 7160 36369 7188
rect 36044 7148 36050 7160
rect 36357 7157 36369 7160
rect 36403 7188 36415 7191
rect 36630 7188 36636 7200
rect 36403 7160 36636 7188
rect 36403 7157 36415 7160
rect 36357 7151 36415 7157
rect 36630 7148 36636 7160
rect 36688 7148 36694 7200
rect 37001 7191 37059 7197
rect 37001 7157 37013 7191
rect 37047 7188 37059 7191
rect 37366 7188 37372 7200
rect 37047 7160 37372 7188
rect 37047 7157 37059 7160
rect 37001 7151 37059 7157
rect 37366 7148 37372 7160
rect 37424 7148 37430 7200
rect 1104 7098 42504 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 42504 7098
rect 1104 7024 42504 7046
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 4430 6984 4436 6996
rect 3016 6956 4436 6984
rect 3016 6944 3022 6956
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6086 6984 6092 6996
rect 5592 6956 6092 6984
rect 5592 6944 5598 6956
rect 6086 6944 6092 6956
rect 6144 6984 6150 6996
rect 6641 6987 6699 6993
rect 6641 6984 6653 6987
rect 6144 6956 6653 6984
rect 6144 6944 6150 6956
rect 6641 6953 6653 6956
rect 6687 6953 6699 6987
rect 6641 6947 6699 6953
rect 8570 6944 8576 6996
rect 8628 6944 8634 6996
rect 8754 6944 8760 6996
rect 8812 6944 8818 6996
rect 8941 6987 8999 6993
rect 8941 6953 8953 6987
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 10400 6987 10458 6993
rect 10400 6953 10412 6987
rect 10446 6984 10458 6987
rect 10870 6984 10876 6996
rect 10446 6956 10876 6984
rect 10446 6953 10458 6956
rect 10400 6947 10458 6953
rect 3050 6876 3056 6928
rect 3108 6916 3114 6928
rect 3786 6916 3792 6928
rect 3108 6888 3792 6916
rect 3108 6876 3114 6888
rect 3528 6857 3556 6888
rect 3786 6876 3792 6888
rect 3844 6876 3850 6928
rect 3988 6888 4752 6916
rect 3513 6851 3571 6857
rect 2608 6820 3188 6848
rect 2608 6789 2636 6820
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6749 2651 6783
rect 2593 6743 2651 6749
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 2792 6712 2820 6743
rect 2866 6740 2872 6792
rect 2924 6740 2930 6792
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 3160 6721 3188 6820
rect 3513 6817 3525 6851
rect 3559 6817 3571 6851
rect 3988 6848 4016 6888
rect 3513 6811 3571 6817
rect 3804 6820 4016 6848
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3804 6789 3832 6820
rect 3329 6783 3387 6789
rect 3329 6780 3341 6783
rect 3292 6752 3341 6780
rect 3292 6740 3298 6752
rect 3329 6749 3341 6752
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2792 6684 2973 6712
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 3145 6715 3203 6721
rect 3145 6681 3157 6715
rect 3191 6712 3203 6715
rect 3804 6712 3832 6743
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4028 6752 4476 6780
rect 4028 6740 4034 6752
rect 3191 6684 3832 6712
rect 3191 6681 3203 6684
rect 3145 6675 3203 6681
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 2685 6647 2743 6653
rect 2685 6644 2697 6647
rect 1728 6616 2697 6644
rect 1728 6604 1734 6616
rect 2685 6613 2697 6616
rect 2731 6613 2743 6647
rect 2685 6607 2743 6613
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3384 6616 3893 6644
rect 3384 6604 3390 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 4448 6644 4476 6752
rect 4614 6740 4620 6792
rect 4672 6740 4678 6792
rect 4724 6780 4752 6888
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 7101 6919 7159 6925
rect 7101 6916 7113 6919
rect 6052 6888 7113 6916
rect 6052 6876 6058 6888
rect 7101 6885 7113 6888
rect 7147 6885 7159 6919
rect 7101 6879 7159 6885
rect 7837 6919 7895 6925
rect 7837 6885 7849 6919
rect 7883 6885 7895 6919
rect 8588 6916 8616 6944
rect 8956 6916 8984 6947
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11882 6944 11888 6996
rect 11940 6944 11946 6996
rect 19610 6944 19616 6996
rect 19668 6944 19674 6996
rect 20530 6944 20536 6996
rect 20588 6984 20594 6996
rect 21097 6987 21155 6993
rect 21097 6984 21109 6987
rect 20588 6956 21109 6984
rect 20588 6944 20594 6956
rect 21097 6953 21109 6956
rect 21143 6953 21155 6987
rect 21097 6947 21155 6953
rect 24118 6944 24124 6996
rect 24176 6984 24182 6996
rect 24397 6987 24455 6993
rect 24397 6984 24409 6987
rect 24176 6956 24409 6984
rect 24176 6944 24182 6956
rect 24397 6953 24409 6956
rect 24443 6953 24455 6987
rect 24397 6947 24455 6953
rect 25406 6944 25412 6996
rect 25464 6984 25470 6996
rect 25881 6987 25939 6993
rect 25881 6984 25893 6987
rect 25464 6956 25893 6984
rect 25464 6944 25470 6956
rect 25881 6953 25893 6956
rect 25927 6953 25939 6987
rect 25881 6947 25939 6953
rect 26500 6987 26558 6993
rect 26500 6953 26512 6987
rect 26546 6984 26558 6987
rect 26970 6984 26976 6996
rect 26546 6956 26976 6984
rect 26546 6953 26558 6956
rect 26500 6947 26558 6953
rect 26970 6944 26976 6956
rect 27028 6944 27034 6996
rect 27798 6944 27804 6996
rect 27856 6984 27862 6996
rect 28905 6987 28963 6993
rect 28905 6984 28917 6987
rect 27856 6956 28917 6984
rect 27856 6944 27862 6956
rect 28905 6953 28917 6956
rect 28951 6953 28963 6987
rect 28905 6947 28963 6953
rect 8588 6888 8984 6916
rect 7837 6879 7895 6885
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5902 6848 5908 6860
rect 5307 6820 5908 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5902 6808 5908 6820
rect 5960 6848 5966 6860
rect 6546 6848 6552 6860
rect 5960 6820 6552 6848
rect 5960 6808 5966 6820
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 7653 6851 7711 6857
rect 6871 6820 7052 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 4724 6752 5457 6780
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 5718 6780 5724 6792
rect 5583 6752 5724 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 5718 6740 5724 6752
rect 5776 6780 5782 6792
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 5776 6752 6469 6780
rect 5776 6740 5782 6752
rect 6457 6749 6469 6752
rect 6503 6780 6515 6783
rect 6641 6783 6699 6789
rect 6641 6780 6653 6783
rect 6503 6752 6653 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 6641 6749 6653 6752
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 5813 6715 5871 6721
rect 5813 6681 5825 6715
rect 5859 6712 5871 6715
rect 5994 6712 6000 6724
rect 5859 6684 6000 6712
rect 5859 6681 5871 6684
rect 5813 6675 5871 6681
rect 5994 6672 6000 6684
rect 6052 6712 6058 6724
rect 6932 6712 6960 6743
rect 6052 6684 6960 6712
rect 7024 6712 7052 6820
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 7852 6848 7880 6879
rect 7699 6820 7880 6848
rect 8205 6851 8263 6857
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 8386 6848 8392 6860
rect 8251 6820 8392 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 9030 6808 9036 6860
rect 9088 6808 9094 6860
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 11054 6848 11060 6860
rect 10183 6820 11060 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 18414 6808 18420 6860
rect 18472 6848 18478 6860
rect 21361 6851 21419 6857
rect 21361 6848 21373 6851
rect 18472 6820 21373 6848
rect 18472 6808 18478 6820
rect 21361 6817 21373 6820
rect 21407 6848 21419 6851
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21407 6820 21465 6848
rect 21407 6817 21419 6820
rect 21361 6811 21419 6817
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 23566 6808 23572 6860
rect 23624 6848 23630 6860
rect 26145 6851 26203 6857
rect 26145 6848 26157 6851
rect 23624 6820 26157 6848
rect 23624 6808 23630 6820
rect 26145 6817 26157 6820
rect 26191 6848 26203 6851
rect 26234 6848 26240 6860
rect 26191 6820 26240 6848
rect 26191 6817 26203 6820
rect 26145 6811 26203 6817
rect 26234 6808 26240 6820
rect 26292 6848 26298 6860
rect 28718 6848 28724 6860
rect 26292 6820 28724 6848
rect 26292 6808 26298 6820
rect 28718 6808 28724 6820
rect 28776 6808 28782 6860
rect 7098 6740 7104 6792
rect 7156 6780 7162 6792
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 7156 6752 7205 6780
rect 7156 6740 7162 6752
rect 7193 6749 7205 6752
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 7466 6740 7472 6792
rect 7524 6740 7530 6792
rect 9122 6780 9128 6792
rect 8404 6752 9128 6780
rect 8404 6721 8432 6752
rect 9122 6740 9128 6752
rect 9180 6780 9186 6792
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 9180 6752 9229 6780
rect 9180 6740 9186 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 23750 6740 23756 6792
rect 23808 6740 23814 6792
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6749 23903 6783
rect 23845 6743 23903 6749
rect 24121 6783 24179 6789
rect 24121 6749 24133 6783
rect 24167 6780 24179 6783
rect 24486 6780 24492 6792
rect 24167 6752 24492 6780
rect 24167 6749 24179 6752
rect 24121 6743 24179 6749
rect 7285 6715 7343 6721
rect 7285 6712 7297 6715
rect 7024 6684 7297 6712
rect 6052 6672 6058 6684
rect 5534 6644 5540 6656
rect 4448 6616 5540 6644
rect 3881 6607 3939 6613
rect 5534 6604 5540 6616
rect 5592 6644 5598 6656
rect 5629 6647 5687 6653
rect 5629 6644 5641 6647
rect 5592 6616 5641 6644
rect 5592 6604 5598 6616
rect 5629 6613 5641 6616
rect 5675 6613 5687 6647
rect 5629 6607 5687 6613
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 5776 6616 5917 6644
rect 5776 6604 5782 6616
rect 5905 6613 5917 6616
rect 5951 6613 5963 6647
rect 5905 6607 5963 6613
rect 6362 6604 6368 6656
rect 6420 6644 6426 6656
rect 7024 6644 7052 6684
rect 7285 6681 7297 6684
rect 7331 6681 7343 6715
rect 7285 6675 7343 6681
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6681 8447 6715
rect 8389 6675 8447 6681
rect 8605 6715 8663 6721
rect 8605 6681 8617 6715
rect 8651 6712 8663 6715
rect 8941 6715 8999 6721
rect 8941 6712 8953 6715
rect 8651 6684 8953 6712
rect 8651 6681 8663 6684
rect 8605 6675 8663 6681
rect 8941 6681 8953 6684
rect 8987 6712 8999 6715
rect 9306 6712 9312 6724
rect 8987 6684 9312 6712
rect 8987 6681 8999 6684
rect 8941 6675 8999 6681
rect 9306 6672 9312 6684
rect 9364 6672 9370 6724
rect 10318 6672 10324 6724
rect 10376 6712 10382 6724
rect 21174 6712 21180 6724
rect 10376 6684 10902 6712
rect 20654 6684 21180 6712
rect 10376 6672 10382 6684
rect 21174 6672 21180 6684
rect 21232 6672 21238 6724
rect 21726 6672 21732 6724
rect 21784 6672 21790 6724
rect 23382 6712 23388 6724
rect 22954 6684 23388 6712
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 6420 6616 7052 6644
rect 6420 6604 6426 6616
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7432 6616 7757 6644
rect 7432 6604 7438 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 7745 6607 7803 6613
rect 9398 6604 9404 6656
rect 9456 6604 9462 6656
rect 22462 6604 22468 6656
rect 22520 6644 22526 6656
rect 23014 6644 23020 6656
rect 22520 6616 23020 6644
rect 22520 6604 22526 6616
rect 23014 6604 23020 6616
rect 23072 6644 23078 6656
rect 23201 6647 23259 6653
rect 23201 6644 23213 6647
rect 23072 6616 23213 6644
rect 23072 6604 23078 6616
rect 23201 6613 23213 6616
rect 23247 6613 23259 6647
rect 23201 6607 23259 6613
rect 23474 6604 23480 6656
rect 23532 6644 23538 6656
rect 23569 6647 23627 6653
rect 23569 6644 23581 6647
rect 23532 6616 23581 6644
rect 23532 6604 23538 6616
rect 23569 6613 23581 6616
rect 23615 6613 23627 6647
rect 23860 6644 23888 6743
rect 24486 6740 24492 6752
rect 24544 6740 24550 6792
rect 28261 6783 28319 6789
rect 28261 6780 28273 6783
rect 28000 6752 28273 6780
rect 24210 6672 24216 6724
rect 24268 6672 24274 6724
rect 25590 6712 25596 6724
rect 25438 6684 25596 6712
rect 25590 6672 25596 6684
rect 25648 6672 25654 6724
rect 27798 6712 27804 6724
rect 27738 6684 27804 6712
rect 27798 6672 27804 6684
rect 27856 6672 27862 6724
rect 24946 6644 24952 6656
rect 23860 6616 24952 6644
rect 23569 6607 23627 6613
rect 24946 6604 24952 6616
rect 25004 6604 25010 6656
rect 28000 6653 28028 6752
rect 28261 6749 28273 6752
rect 28307 6749 28319 6783
rect 28920 6780 28948 6947
rect 29270 6944 29276 6996
rect 29328 6984 29334 6996
rect 29549 6987 29607 6993
rect 29549 6984 29561 6987
rect 29328 6956 29561 6984
rect 29328 6944 29334 6956
rect 29549 6953 29561 6956
rect 29595 6953 29607 6987
rect 29549 6947 29607 6953
rect 29638 6944 29644 6996
rect 29696 6984 29702 6996
rect 30834 6984 30840 6996
rect 29696 6956 30840 6984
rect 29696 6944 29702 6956
rect 30834 6944 30840 6956
rect 30892 6944 30898 6996
rect 31754 6984 31760 6996
rect 31036 6956 31760 6984
rect 29454 6876 29460 6928
rect 29512 6916 29518 6928
rect 30282 6916 30288 6928
rect 29512 6888 30288 6916
rect 29512 6876 29518 6888
rect 30282 6876 30288 6888
rect 30340 6876 30346 6928
rect 31036 6925 31064 6956
rect 31754 6944 31760 6956
rect 31812 6984 31818 6996
rect 32766 6984 32772 6996
rect 31812 6956 32772 6984
rect 31812 6944 31818 6956
rect 32766 6944 32772 6956
rect 32824 6944 32830 6996
rect 33032 6987 33090 6993
rect 33032 6953 33044 6987
rect 33078 6984 33090 6987
rect 34698 6984 34704 6996
rect 33078 6956 34704 6984
rect 33078 6953 33090 6956
rect 33032 6947 33090 6953
rect 34698 6944 34704 6956
rect 34756 6944 34762 6996
rect 36446 6944 36452 6996
rect 36504 6944 36510 6996
rect 36814 6944 36820 6996
rect 36872 6984 36878 6996
rect 37185 6987 37243 6993
rect 37185 6984 37197 6987
rect 36872 6956 37197 6984
rect 36872 6944 36878 6956
rect 37185 6953 37197 6956
rect 37231 6953 37243 6987
rect 37185 6947 37243 6953
rect 31021 6919 31079 6925
rect 31021 6885 31033 6919
rect 31067 6885 31079 6919
rect 31021 6879 31079 6885
rect 31570 6876 31576 6928
rect 31628 6876 31634 6928
rect 36722 6916 36728 6928
rect 35820 6888 36728 6916
rect 28994 6808 29000 6860
rect 29052 6848 29058 6860
rect 29052 6820 30144 6848
rect 29052 6808 29058 6820
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 28920 6752 29745 6780
rect 28261 6743 28319 6749
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 29914 6740 29920 6792
rect 29972 6740 29978 6792
rect 30116 6789 30144 6820
rect 30466 6808 30472 6860
rect 30524 6848 30530 6860
rect 30926 6848 30932 6860
rect 30524 6820 30932 6848
rect 30524 6808 30530 6820
rect 30926 6808 30932 6820
rect 30984 6808 30990 6860
rect 31202 6808 31208 6860
rect 31260 6848 31266 6860
rect 32769 6851 32827 6857
rect 32769 6848 32781 6851
rect 31260 6820 32781 6848
rect 31260 6808 31266 6820
rect 32769 6817 32781 6820
rect 32815 6817 32827 6851
rect 32769 6811 32827 6817
rect 34517 6851 34575 6857
rect 34517 6817 34529 6851
rect 34563 6848 34575 6851
rect 34885 6851 34943 6857
rect 34885 6848 34897 6851
rect 34563 6820 34897 6848
rect 34563 6817 34575 6820
rect 34517 6811 34575 6817
rect 34885 6817 34897 6820
rect 34931 6817 34943 6851
rect 34885 6811 34943 6817
rect 30101 6783 30159 6789
rect 30101 6749 30113 6783
rect 30147 6749 30159 6783
rect 30101 6743 30159 6749
rect 30561 6783 30619 6789
rect 30561 6749 30573 6783
rect 30607 6780 30619 6783
rect 31294 6780 31300 6792
rect 30607 6752 31300 6780
rect 30607 6749 30619 6752
rect 30561 6743 30619 6749
rect 31294 6740 31300 6752
rect 31352 6740 31358 6792
rect 31386 6740 31392 6792
rect 31444 6740 31450 6792
rect 34606 6740 34612 6792
rect 34664 6780 34670 6792
rect 35820 6780 35848 6888
rect 36722 6876 36728 6888
rect 36780 6876 36786 6928
rect 35897 6851 35955 6857
rect 35897 6817 35909 6851
rect 35943 6848 35955 6851
rect 36170 6848 36176 6860
rect 35943 6820 36176 6848
rect 35943 6817 35955 6820
rect 35897 6811 35955 6817
rect 36170 6808 36176 6820
rect 36228 6808 36234 6860
rect 36265 6851 36323 6857
rect 36265 6817 36277 6851
rect 36311 6848 36323 6851
rect 36832 6848 36860 6944
rect 36311 6820 36860 6848
rect 36311 6817 36323 6820
rect 36265 6811 36323 6817
rect 34664 6752 35848 6780
rect 34664 6740 34670 6752
rect 35986 6740 35992 6792
rect 36044 6740 36050 6792
rect 36354 6740 36360 6792
rect 36412 6740 36418 6792
rect 36998 6740 37004 6792
rect 37056 6740 37062 6792
rect 37734 6740 37740 6792
rect 37792 6740 37798 6792
rect 38838 6740 38844 6792
rect 38896 6740 38902 6792
rect 29362 6672 29368 6724
rect 29420 6712 29426 6724
rect 29825 6715 29883 6721
rect 29825 6712 29837 6715
rect 29420 6684 29837 6712
rect 29420 6672 29426 6684
rect 29825 6681 29837 6684
rect 29871 6681 29883 6715
rect 29825 6675 29883 6681
rect 31018 6672 31024 6724
rect 31076 6712 31082 6724
rect 31205 6715 31263 6721
rect 31205 6712 31217 6715
rect 31076 6684 31217 6712
rect 31076 6672 31082 6684
rect 31205 6681 31217 6684
rect 31251 6681 31263 6715
rect 34330 6712 34336 6724
rect 34270 6684 34336 6712
rect 31205 6675 31263 6681
rect 34330 6672 34336 6684
rect 34388 6672 34394 6724
rect 35434 6672 35440 6724
rect 35492 6712 35498 6724
rect 35492 6684 35756 6712
rect 35492 6672 35498 6684
rect 27985 6647 28043 6653
rect 27985 6613 27997 6647
rect 28031 6613 28043 6647
rect 27985 6607 28043 6613
rect 30190 6604 30196 6656
rect 30248 6604 30254 6656
rect 31294 6604 31300 6656
rect 31352 6604 31358 6656
rect 34790 6604 34796 6656
rect 34848 6644 34854 6656
rect 35728 6653 35756 6684
rect 36262 6672 36268 6724
rect 36320 6712 36326 6724
rect 37921 6715 37979 6721
rect 37921 6712 37933 6715
rect 36320 6684 37933 6712
rect 36320 6672 36326 6684
rect 37921 6681 37933 6684
rect 37967 6681 37979 6715
rect 37921 6675 37979 6681
rect 38286 6672 38292 6724
rect 38344 6712 38350 6724
rect 38473 6715 38531 6721
rect 38473 6712 38485 6715
rect 38344 6684 38485 6712
rect 38344 6672 38350 6684
rect 38473 6681 38485 6684
rect 38519 6681 38531 6715
rect 38473 6675 38531 6681
rect 35529 6647 35587 6653
rect 35529 6644 35541 6647
rect 34848 6616 35541 6644
rect 34848 6604 34854 6616
rect 35529 6613 35541 6616
rect 35575 6613 35587 6647
rect 35529 6607 35587 6613
rect 35713 6647 35771 6653
rect 35713 6613 35725 6647
rect 35759 6613 35771 6647
rect 35713 6607 35771 6613
rect 1104 6554 42504 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 42504 6554
rect 1104 6480 42504 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 4614 6440 4620 6452
rect 1452 6412 4620 6440
rect 1452 6400 1458 6412
rect 1670 6332 1676 6384
rect 1728 6332 1734 6384
rect 2958 6372 2964 6384
rect 2898 6344 2964 6372
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 3234 6332 3240 6384
rect 3292 6372 3298 6384
rect 3481 6375 3539 6381
rect 3481 6372 3493 6375
rect 3292 6344 3493 6372
rect 3292 6332 3298 6344
rect 3481 6341 3493 6344
rect 3527 6341 3539 6375
rect 3481 6335 3539 6341
rect 3697 6375 3755 6381
rect 3697 6341 3709 6375
rect 3743 6372 3755 6375
rect 3786 6372 3792 6384
rect 3743 6344 3792 6372
rect 3743 6341 3755 6344
rect 3697 6335 3755 6341
rect 1394 6264 1400 6316
rect 1452 6264 1458 6316
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3712 6236 3740 6335
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 3878 6264 3884 6316
rect 3936 6264 3942 6316
rect 4062 6264 4068 6316
rect 4120 6264 4126 6316
rect 4172 6313 4200 6412
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 6733 6443 6791 6449
rect 6733 6409 6745 6443
rect 6779 6440 6791 6443
rect 8386 6440 8392 6452
rect 6779 6412 8392 6440
rect 6779 6409 6791 6412
rect 6733 6403 6791 6409
rect 8386 6400 8392 6412
rect 8444 6440 8450 6452
rect 8846 6440 8852 6452
rect 8444 6412 8852 6440
rect 8444 6400 8450 6412
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 10376 6412 10609 6440
rect 10376 6400 10382 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 11057 6443 11115 6449
rect 11057 6409 11069 6443
rect 11103 6409 11115 6443
rect 11057 6403 11115 6409
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 4706 6372 4712 6384
rect 4488 6344 4712 6372
rect 4488 6332 4494 6344
rect 4706 6332 4712 6344
rect 4764 6372 4770 6384
rect 4764 6344 4922 6372
rect 4764 6332 4770 6344
rect 6362 6332 6368 6384
rect 6420 6332 6426 6384
rect 6546 6332 6552 6384
rect 6604 6381 6610 6384
rect 6604 6375 6639 6381
rect 6627 6372 6639 6375
rect 7006 6372 7012 6384
rect 6627 6344 7012 6372
rect 6627 6341 6639 6344
rect 6604 6335 6639 6341
rect 6604 6332 6610 6335
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 7101 6375 7159 6381
rect 7101 6341 7113 6375
rect 7147 6372 7159 6375
rect 7374 6372 7380 6384
rect 7147 6344 7380 6372
rect 7147 6341 7159 6344
rect 7101 6335 7159 6341
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 8478 6372 8484 6384
rect 8326 6344 8484 6372
rect 8478 6332 8484 6344
rect 8536 6372 8542 6384
rect 10336 6372 10364 6400
rect 8536 6344 10364 6372
rect 8536 6332 8542 6344
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 10778 6372 10784 6384
rect 10560 6344 10784 6372
rect 10560 6332 10566 6344
rect 10778 6332 10784 6344
rect 10836 6372 10842 6384
rect 11072 6372 11100 6403
rect 20162 6400 20168 6452
rect 20220 6400 20226 6452
rect 23382 6400 23388 6452
rect 23440 6440 23446 6452
rect 24949 6443 25007 6449
rect 23440 6412 24808 6440
rect 23440 6400 23446 6412
rect 10836 6344 11100 6372
rect 10836 6332 10842 6344
rect 18690 6332 18696 6384
rect 18748 6332 18754 6384
rect 20806 6332 20812 6384
rect 20864 6332 20870 6384
rect 21174 6332 21180 6384
rect 21232 6332 21238 6384
rect 23566 6372 23572 6384
rect 23216 6344 23572 6372
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 8895 6276 9321 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 9309 6273 9321 6276
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 9456 6276 9873 6304
rect 9456 6264 9462 6276
rect 9861 6273 9873 6276
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 17954 6304 17960 6316
rect 11287 6276 17960 6304
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 18414 6264 18420 6316
rect 18472 6264 18478 6316
rect 21192 6304 21220 6332
rect 19826 6276 21220 6304
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 23216 6313 23244 6344
rect 23566 6332 23572 6344
rect 23624 6332 23630 6384
rect 24780 6372 24808 6412
rect 24949 6409 24961 6443
rect 24995 6440 25007 6443
rect 26050 6440 26056 6452
rect 24995 6412 26056 6440
rect 24995 6409 25007 6412
rect 24949 6403 25007 6409
rect 26050 6400 26056 6412
rect 26108 6400 26114 6452
rect 26973 6443 27031 6449
rect 26973 6409 26985 6443
rect 27019 6440 27031 6443
rect 27430 6440 27436 6452
rect 27019 6412 27436 6440
rect 27019 6409 27031 6412
rect 26973 6403 27031 6409
rect 27430 6400 27436 6412
rect 27488 6400 27494 6452
rect 27798 6400 27804 6452
rect 27856 6440 27862 6452
rect 29546 6440 29552 6452
rect 27856 6412 29552 6440
rect 27856 6400 27862 6412
rect 25133 6375 25191 6381
rect 25133 6372 25145 6375
rect 24702 6344 25145 6372
rect 25133 6341 25145 6344
rect 25179 6372 25191 6375
rect 25590 6372 25596 6384
rect 25179 6344 25596 6372
rect 25179 6341 25191 6344
rect 25133 6335 25191 6341
rect 25590 6332 25596 6344
rect 25648 6332 25654 6384
rect 28092 6372 28120 6412
rect 29546 6400 29552 6412
rect 29604 6400 29610 6452
rect 31846 6440 31852 6452
rect 31496 6412 31852 6440
rect 28014 6344 28120 6372
rect 28442 6332 28448 6384
rect 28500 6332 28506 6384
rect 30190 6372 30196 6384
rect 29104 6344 30196 6372
rect 29104 6313 29132 6344
rect 30190 6332 30196 6344
rect 30248 6332 30254 6384
rect 30650 6332 30656 6384
rect 30708 6372 30714 6384
rect 30929 6375 30987 6381
rect 30929 6372 30941 6375
rect 30708 6344 30941 6372
rect 30708 6332 30714 6344
rect 30929 6341 30941 6344
rect 30975 6372 30987 6375
rect 31496 6372 31524 6412
rect 31846 6400 31852 6412
rect 31904 6400 31910 6452
rect 33042 6400 33048 6452
rect 33100 6440 33106 6452
rect 34330 6440 34336 6452
rect 33100 6412 34336 6440
rect 33100 6400 33106 6412
rect 34330 6400 34336 6412
rect 34388 6440 34394 6452
rect 36262 6440 36268 6452
rect 34388 6412 36268 6440
rect 34388 6400 34394 6412
rect 32674 6372 32680 6384
rect 30975 6344 31524 6372
rect 31588 6344 32680 6372
rect 30975 6341 30987 6344
rect 30929 6335 30987 6341
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21876 6276 22017 6304
rect 21876 6264 21882 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 23201 6307 23259 6313
rect 23201 6273 23213 6307
rect 23247 6273 23259 6307
rect 23201 6267 23259 6273
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6273 25559 6307
rect 25501 6267 25559 6273
rect 29089 6307 29147 6313
rect 29089 6273 29101 6307
rect 29135 6273 29147 6307
rect 29089 6267 29147 6273
rect 29365 6307 29423 6313
rect 29365 6273 29377 6307
rect 29411 6304 29423 6307
rect 30469 6307 30527 6313
rect 30469 6304 30481 6307
rect 29411 6276 30481 6304
rect 29411 6273 29423 6276
rect 29365 6267 29423 6273
rect 30469 6273 30481 6276
rect 30515 6304 30527 6307
rect 30745 6307 30803 6313
rect 30745 6304 30757 6307
rect 30515 6276 30757 6304
rect 30515 6273 30527 6276
rect 30469 6267 30527 6273
rect 30745 6273 30757 6276
rect 30791 6273 30803 6307
rect 30745 6267 30803 6273
rect 3191 6208 3740 6236
rect 3973 6239 4031 6245
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4433 6239 4491 6245
rect 4433 6236 4445 6239
rect 4019 6208 4445 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4433 6205 4445 6208
rect 4479 6205 4491 6239
rect 4433 6199 4491 6205
rect 5902 6196 5908 6248
rect 5960 6196 5966 6248
rect 6822 6196 6828 6248
rect 6880 6196 6886 6248
rect 8938 6196 8944 6248
rect 8996 6196 9002 6248
rect 23474 6196 23480 6248
rect 23532 6196 23538 6248
rect 25516 6236 25544 6267
rect 30834 6264 30840 6316
rect 30892 6264 30898 6316
rect 31113 6307 31171 6313
rect 31113 6273 31125 6307
rect 31159 6304 31171 6307
rect 31294 6304 31300 6316
rect 31159 6276 31300 6304
rect 31159 6273 31171 6276
rect 31113 6267 31171 6273
rect 31294 6264 31300 6276
rect 31352 6264 31358 6316
rect 31588 6313 31616 6344
rect 32674 6332 32680 6344
rect 32732 6332 32738 6384
rect 34348 6372 34376 6400
rect 35342 6372 35348 6384
rect 34270 6344 34376 6372
rect 35176 6344 35348 6372
rect 31573 6307 31631 6313
rect 31573 6273 31585 6307
rect 31619 6273 31631 6307
rect 31573 6267 31631 6273
rect 31662 6264 31668 6316
rect 31720 6264 31726 6316
rect 31757 6307 31815 6313
rect 31757 6273 31769 6307
rect 31803 6304 31815 6307
rect 31846 6304 31852 6316
rect 31803 6276 31852 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 31846 6264 31852 6276
rect 31904 6264 31910 6316
rect 31938 6264 31944 6316
rect 31996 6264 32002 6316
rect 32398 6264 32404 6316
rect 32456 6264 32462 6316
rect 32582 6264 32588 6316
rect 32640 6304 32646 6316
rect 35176 6313 35204 6344
rect 35342 6332 35348 6344
rect 35400 6332 35406 6384
rect 35434 6332 35440 6384
rect 35492 6332 35498 6384
rect 35820 6372 35848 6412
rect 36262 6400 36268 6412
rect 36320 6400 36326 6452
rect 36909 6443 36967 6449
rect 36909 6409 36921 6443
rect 36955 6440 36967 6443
rect 37734 6440 37740 6452
rect 36955 6412 37740 6440
rect 36955 6409 36967 6412
rect 36909 6403 36967 6409
rect 37734 6400 37740 6412
rect 37792 6400 37798 6452
rect 35820 6344 35926 6372
rect 32769 6307 32827 6313
rect 32769 6304 32781 6307
rect 32640 6276 32781 6304
rect 32640 6264 32646 6276
rect 32769 6273 32781 6276
rect 32815 6273 32827 6307
rect 32769 6267 32827 6273
rect 34977 6307 35035 6313
rect 34977 6273 34989 6307
rect 35023 6304 35035 6307
rect 35161 6307 35219 6313
rect 35161 6304 35173 6307
rect 35023 6276 35173 6304
rect 35023 6273 35035 6276
rect 34977 6267 35035 6273
rect 35161 6273 35173 6276
rect 35207 6273 35219 6307
rect 35161 6267 35219 6273
rect 37277 6307 37335 6313
rect 37277 6273 37289 6307
rect 37323 6304 37335 6307
rect 41966 6304 41972 6316
rect 37323 6276 41972 6304
rect 37323 6273 37335 6276
rect 37277 6267 37335 6273
rect 25516 6208 28672 6236
rect 5920 6168 5948 6196
rect 5460 6140 5948 6168
rect 9217 6171 9275 6177
rect 3329 6103 3387 6109
rect 3329 6069 3341 6103
rect 3375 6100 3387 6103
rect 3418 6100 3424 6112
rect 3375 6072 3424 6100
rect 3375 6069 3387 6072
rect 3329 6063 3387 6069
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 3970 6100 3976 6112
rect 3568 6072 3976 6100
rect 3568 6060 3574 6072
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 5460 6100 5488 6140
rect 9217 6137 9229 6171
rect 9263 6168 9275 6171
rect 10778 6168 10784 6180
rect 9263 6140 10784 6168
rect 9263 6137 9275 6140
rect 9217 6131 9275 6137
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 28644 6168 28672 6208
rect 28718 6196 28724 6248
rect 28776 6196 28782 6248
rect 28997 6239 29055 6245
rect 28997 6205 29009 6239
rect 29043 6205 29055 6239
rect 28997 6199 29055 6205
rect 29012 6168 29040 6199
rect 29454 6196 29460 6248
rect 29512 6196 29518 6248
rect 29914 6196 29920 6248
rect 29972 6196 29978 6248
rect 30006 6196 30012 6248
rect 30064 6236 30070 6248
rect 32309 6239 32367 6245
rect 32309 6236 32321 6239
rect 30064 6208 32321 6236
rect 30064 6196 30070 6208
rect 32309 6205 32321 6208
rect 32355 6205 32367 6239
rect 32309 6199 32367 6205
rect 34698 6196 34704 6248
rect 34756 6196 34762 6248
rect 29086 6168 29092 6180
rect 28644 6140 28948 6168
rect 29012 6140 29092 6168
rect 4120 6072 5488 6100
rect 4120 6060 4126 6072
rect 5810 6060 5816 6112
rect 5868 6100 5874 6112
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 5868 6072 5917 6100
rect 5868 6060 5874 6072
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 6549 6103 6607 6109
rect 6549 6069 6561 6103
rect 6595 6100 6607 6103
rect 7466 6100 7472 6112
rect 6595 6072 7472 6100
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 7466 6060 7472 6072
rect 7524 6100 7530 6112
rect 8570 6100 8576 6112
rect 7524 6072 8576 6100
rect 7524 6060 7530 6072
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 22646 6060 22652 6112
rect 22704 6060 22710 6112
rect 28442 6060 28448 6112
rect 28500 6100 28506 6112
rect 28813 6103 28871 6109
rect 28813 6100 28825 6103
rect 28500 6072 28825 6100
rect 28500 6060 28506 6072
rect 28813 6069 28825 6072
rect 28859 6069 28871 6103
rect 28920 6100 28948 6140
rect 29086 6128 29092 6140
rect 29144 6168 29150 6180
rect 30024 6168 30052 6196
rect 29144 6140 30052 6168
rect 31389 6171 31447 6177
rect 29144 6128 29150 6140
rect 31389 6137 31401 6171
rect 31435 6168 31447 6171
rect 31478 6168 31484 6180
rect 31435 6140 31484 6168
rect 31435 6137 31447 6140
rect 31389 6131 31447 6137
rect 31478 6128 31484 6140
rect 31536 6128 31542 6180
rect 31588 6140 33732 6168
rect 30466 6100 30472 6112
rect 28920 6072 30472 6100
rect 28813 6063 28871 6069
rect 30466 6060 30472 6072
rect 30524 6060 30530 6112
rect 30558 6060 30564 6112
rect 30616 6060 30622 6112
rect 30742 6060 30748 6112
rect 30800 6100 30806 6112
rect 31588 6100 31616 6140
rect 30800 6072 31616 6100
rect 30800 6060 30806 6072
rect 32122 6060 32128 6112
rect 32180 6060 32186 6112
rect 33226 6060 33232 6112
rect 33284 6060 33290 6112
rect 33704 6100 33732 6140
rect 37292 6100 37320 6267
rect 41966 6264 41972 6276
rect 42024 6264 42030 6316
rect 37458 6128 37464 6180
rect 37516 6168 37522 6180
rect 38746 6168 38752 6180
rect 37516 6140 38752 6168
rect 37516 6128 37522 6140
rect 38746 6128 38752 6140
rect 38804 6128 38810 6180
rect 33704 6072 37320 6100
rect 1104 6010 42504 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 42504 6010
rect 1104 5936 42504 5958
rect 3510 5856 3516 5908
rect 3568 5856 3574 5908
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 4062 5896 4068 5908
rect 3835 5868 4068 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 4764 5868 7236 5896
rect 4764 5856 4770 5868
rect 3878 5788 3884 5840
rect 3936 5828 3942 5840
rect 5721 5831 5779 5837
rect 5721 5828 5733 5831
rect 3936 5800 5733 5828
rect 3936 5788 3942 5800
rect 5721 5797 5733 5800
rect 5767 5797 5779 5831
rect 5721 5791 5779 5797
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1765 5763 1823 5769
rect 1765 5760 1777 5763
rect 1452 5732 1777 5760
rect 1452 5720 1458 5732
rect 1765 5729 1777 5732
rect 1811 5729 1823 5763
rect 1765 5723 1823 5729
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5760 2099 5763
rect 3234 5760 3240 5772
rect 2087 5732 3240 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3476 5732 4077 5760
rect 3476 5720 3482 5732
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 3108 5664 3174 5692
rect 3108 5652 3114 5664
rect 4080 5624 4108 5723
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 4614 5760 4620 5772
rect 4396 5732 4620 5760
rect 4396 5720 4402 5732
rect 4614 5720 4620 5732
rect 4672 5760 4678 5772
rect 5905 5763 5963 5769
rect 5905 5760 5917 5763
rect 4672 5732 5917 5760
rect 4672 5720 4678 5732
rect 5905 5729 5917 5732
rect 5951 5760 5963 5763
rect 6822 5760 6828 5772
rect 5951 5732 6828 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 7208 5704 7236 5868
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8996 5868 9045 5896
rect 8996 5856 9002 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 9306 5856 9312 5908
rect 9364 5856 9370 5908
rect 21726 5856 21732 5908
rect 21784 5896 21790 5908
rect 21821 5899 21879 5905
rect 21821 5896 21833 5899
rect 21784 5868 21833 5896
rect 21784 5856 21790 5868
rect 21821 5865 21833 5868
rect 21867 5865 21879 5899
rect 21821 5859 21879 5865
rect 22557 5899 22615 5905
rect 22557 5865 22569 5899
rect 22603 5896 22615 5899
rect 23290 5896 23296 5908
rect 22603 5868 23296 5896
rect 22603 5865 22615 5868
rect 22557 5859 22615 5865
rect 23290 5856 23296 5868
rect 23348 5856 23354 5908
rect 31294 5856 31300 5908
rect 31352 5856 31358 5908
rect 32674 5856 32680 5908
rect 32732 5896 32738 5908
rect 33229 5899 33287 5905
rect 33229 5896 33241 5899
rect 32732 5868 33241 5896
rect 32732 5856 32738 5868
rect 33229 5865 33241 5868
rect 33275 5865 33287 5899
rect 33229 5859 33287 5865
rect 35897 5899 35955 5905
rect 35897 5865 35909 5899
rect 35943 5896 35955 5899
rect 36998 5896 37004 5908
rect 35943 5868 37004 5896
rect 35943 5865 35955 5868
rect 35897 5859 35955 5865
rect 36998 5856 37004 5868
rect 37056 5856 37062 5908
rect 41966 5856 41972 5908
rect 42024 5856 42030 5908
rect 10410 5760 10416 5772
rect 7576 5732 10416 5760
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4798 5692 4804 5704
rect 4203 5664 4804 5692
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 4908 5664 5457 5692
rect 4908 5624 4936 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 5718 5652 5724 5704
rect 5776 5652 5782 5704
rect 7190 5652 7196 5704
rect 7248 5692 7254 5704
rect 7248 5664 7314 5692
rect 7248 5652 7254 5664
rect 4080 5596 4936 5624
rect 5353 5627 5411 5633
rect 5353 5593 5365 5627
rect 5399 5624 5411 5627
rect 5399 5596 6132 5624
rect 5399 5593 5411 5596
rect 5353 5587 5411 5593
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 6104 5556 6132 5596
rect 6178 5584 6184 5636
rect 6236 5584 6242 5636
rect 7576 5556 7604 5732
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 10778 5720 10784 5772
rect 10836 5720 10842 5772
rect 11054 5720 11060 5772
rect 11112 5720 11118 5772
rect 22741 5763 22799 5769
rect 22741 5729 22753 5763
rect 22787 5760 22799 5763
rect 23750 5760 23756 5772
rect 22787 5732 23756 5760
rect 22787 5729 22799 5732
rect 22741 5723 22799 5729
rect 23750 5720 23756 5732
rect 23808 5720 23814 5772
rect 28718 5720 28724 5772
rect 28776 5760 28782 5772
rect 29549 5763 29607 5769
rect 29549 5760 29561 5763
rect 28776 5732 29561 5760
rect 28776 5720 28782 5732
rect 29549 5729 29561 5732
rect 29595 5729 29607 5763
rect 29549 5723 29607 5729
rect 29825 5763 29883 5769
rect 29825 5729 29837 5763
rect 29871 5760 29883 5763
rect 30558 5760 30564 5772
rect 29871 5732 30564 5760
rect 29871 5729 29883 5732
rect 29825 5723 29883 5729
rect 30558 5720 30564 5732
rect 30616 5720 30622 5772
rect 31665 5763 31723 5769
rect 31665 5729 31677 5763
rect 31711 5760 31723 5763
rect 32122 5760 32128 5772
rect 31711 5732 32128 5760
rect 31711 5729 31723 5732
rect 31665 5723 31723 5729
rect 32122 5720 32128 5732
rect 32180 5720 32186 5772
rect 33137 5763 33195 5769
rect 33137 5729 33149 5763
rect 33183 5760 33195 5763
rect 33781 5763 33839 5769
rect 33781 5760 33793 5763
rect 33183 5732 33793 5760
rect 33183 5729 33195 5732
rect 33137 5723 33195 5729
rect 33781 5729 33793 5732
rect 33827 5729 33839 5763
rect 33781 5723 33839 5729
rect 37366 5720 37372 5772
rect 37424 5720 37430 5772
rect 37642 5720 37648 5772
rect 37700 5720 37706 5772
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 8772 5624 8800 5655
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8904 5664 8953 5692
rect 8904 5652 8910 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9122 5652 9128 5704
rect 9180 5652 9186 5704
rect 22370 5652 22376 5704
rect 22428 5652 22434 5704
rect 22830 5652 22836 5704
rect 22888 5652 22894 5704
rect 23201 5695 23259 5701
rect 23201 5661 23213 5695
rect 23247 5692 23259 5695
rect 24210 5692 24216 5704
rect 23247 5664 24216 5692
rect 23247 5661 23259 5664
rect 23201 5655 23259 5661
rect 24210 5652 24216 5664
rect 24268 5652 24274 5704
rect 31202 5652 31208 5704
rect 31260 5692 31266 5704
rect 31389 5695 31447 5701
rect 31389 5692 31401 5695
rect 31260 5664 31401 5692
rect 31260 5652 31266 5664
rect 31389 5661 31401 5664
rect 31435 5661 31447 5695
rect 31389 5655 31447 5661
rect 33226 5652 33232 5704
rect 33284 5692 33290 5704
rect 34146 5692 34152 5704
rect 33284 5664 34152 5692
rect 33284 5652 33290 5664
rect 34146 5652 34152 5664
rect 34204 5692 34210 5704
rect 34701 5695 34759 5701
rect 34701 5692 34713 5695
rect 34204 5664 34713 5692
rect 34204 5652 34210 5664
rect 34701 5661 34713 5664
rect 34747 5661 34759 5695
rect 34701 5655 34759 5661
rect 9140 5624 9168 5652
rect 8772 5596 9168 5624
rect 10318 5584 10324 5636
rect 10376 5624 10382 5636
rect 10376 5596 10456 5624
rect 10376 5584 10382 5596
rect 6104 5528 7604 5556
rect 7650 5516 7656 5568
rect 7708 5516 7714 5568
rect 8113 5559 8171 5565
rect 8113 5525 8125 5559
rect 8159 5556 8171 5559
rect 8386 5556 8392 5568
rect 8159 5528 8392 5556
rect 8159 5525 8171 5528
rect 8113 5519 8171 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 10428 5556 10456 5596
rect 22094 5584 22100 5636
rect 22152 5624 22158 5636
rect 22646 5624 22652 5636
rect 22152 5596 22652 5624
rect 22152 5584 22158 5596
rect 22646 5584 22652 5596
rect 22704 5624 22710 5636
rect 23109 5627 23167 5633
rect 23109 5624 23121 5627
rect 22704 5596 23121 5624
rect 22704 5584 22710 5596
rect 23109 5593 23121 5596
rect 23155 5593 23167 5627
rect 23109 5587 23167 5593
rect 29546 5584 29552 5636
rect 29604 5624 29610 5636
rect 33042 5624 33048 5636
rect 29604 5596 30314 5624
rect 32890 5596 33048 5624
rect 29604 5584 29610 5596
rect 33042 5584 33048 5596
rect 33100 5584 33106 5636
rect 38286 5624 38292 5636
rect 36938 5596 38292 5624
rect 38286 5584 38292 5596
rect 38344 5584 38350 5636
rect 42058 5584 42064 5636
rect 42116 5584 42122 5636
rect 9548 5528 10456 5556
rect 9548 5516 9554 5528
rect 22922 5516 22928 5568
rect 22980 5556 22986 5568
rect 30742 5556 30748 5568
rect 22980 5528 30748 5556
rect 22980 5516 22986 5528
rect 30742 5516 30748 5528
rect 30800 5516 30806 5568
rect 30834 5516 30840 5568
rect 30892 5556 30898 5568
rect 31662 5556 31668 5568
rect 30892 5528 31668 5556
rect 30892 5516 30898 5528
rect 31662 5516 31668 5528
rect 31720 5556 31726 5568
rect 34606 5556 34612 5568
rect 31720 5528 34612 5556
rect 31720 5516 31726 5528
rect 34606 5516 34612 5528
rect 34664 5516 34670 5568
rect 35250 5516 35256 5568
rect 35308 5556 35314 5568
rect 35345 5559 35403 5565
rect 35345 5556 35357 5559
rect 35308 5528 35357 5556
rect 35308 5516 35314 5528
rect 35345 5525 35357 5528
rect 35391 5525 35403 5559
rect 35345 5519 35403 5525
rect 1104 5466 42504 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 42504 5466
rect 1104 5392 42504 5414
rect 3234 5312 3240 5364
rect 3292 5312 3298 5364
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5994 5352 6000 5364
rect 5592 5324 6000 5352
rect 5592 5312 5598 5324
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 9122 5312 9128 5364
rect 9180 5352 9186 5364
rect 9585 5355 9643 5361
rect 9585 5352 9597 5355
rect 9180 5324 9597 5352
rect 9180 5312 9186 5324
rect 9585 5321 9597 5324
rect 9631 5321 9643 5355
rect 9585 5315 9643 5321
rect 29914 5312 29920 5364
rect 29972 5312 29978 5364
rect 31938 5312 31944 5364
rect 31996 5352 32002 5364
rect 32125 5355 32183 5361
rect 32125 5352 32137 5355
rect 31996 5324 32137 5352
rect 31996 5312 32002 5324
rect 32125 5321 32137 5324
rect 32171 5321 32183 5355
rect 32125 5315 32183 5321
rect 34698 5312 34704 5364
rect 34756 5312 34762 5364
rect 3418 5284 3424 5296
rect 3160 5256 3424 5284
rect 3160 5225 3188 5256
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 4338 5284 4344 5296
rect 3804 5256 4344 5284
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 3804 5225 3832 5256
rect 4338 5244 4344 5256
rect 4396 5244 4402 5296
rect 4706 5244 4712 5296
rect 4764 5244 4770 5296
rect 9490 5284 9496 5296
rect 9338 5256 9496 5284
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 22186 5244 22192 5296
rect 22244 5244 22250 5296
rect 22278 5244 22284 5296
rect 22336 5244 22342 5296
rect 28718 5284 28724 5296
rect 28184 5256 28724 5284
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 5859 5188 6745 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 6880 5188 7849 5216
rect 6880 5176 6886 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 22094 5176 22100 5228
rect 22152 5176 22158 5228
rect 22462 5176 22468 5228
rect 22520 5176 22526 5228
rect 28184 5225 28212 5256
rect 28718 5244 28724 5256
rect 28776 5244 28782 5296
rect 30650 5244 30656 5296
rect 30708 5284 30714 5296
rect 30837 5287 30895 5293
rect 30837 5284 30849 5287
rect 30708 5256 30849 5284
rect 30708 5244 30714 5256
rect 30837 5253 30849 5256
rect 30883 5253 30895 5287
rect 30837 5247 30895 5253
rect 31021 5287 31079 5293
rect 31021 5253 31033 5287
rect 31067 5284 31079 5287
rect 31067 5256 34560 5284
rect 31067 5253 31079 5256
rect 31021 5247 31079 5253
rect 28169 5219 28227 5225
rect 28169 5185 28181 5219
rect 28215 5185 28227 5219
rect 28169 5179 28227 5185
rect 29546 5176 29552 5228
rect 29604 5216 29610 5228
rect 30285 5219 30343 5225
rect 30285 5216 30297 5219
rect 29604 5188 30297 5216
rect 29604 5176 29610 5188
rect 30285 5185 30297 5188
rect 30331 5185 30343 5219
rect 30285 5179 30343 5185
rect 4062 5108 4068 5160
rect 4120 5108 4126 5160
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 6178 5108 6184 5160
rect 6236 5108 6242 5160
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 6638 5148 6644 5160
rect 6420 5120 6644 5148
rect 6420 5108 6426 5120
rect 6638 5108 6644 5120
rect 6696 5148 6702 5160
rect 7285 5151 7343 5157
rect 7285 5148 7297 5151
rect 6696 5120 7297 5148
rect 6696 5108 6702 5120
rect 7285 5117 7297 5120
rect 7331 5148 7343 5151
rect 7650 5148 7656 5160
rect 7331 5120 7656 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 8110 5108 8116 5160
rect 8168 5108 8174 5160
rect 28442 5108 28448 5160
rect 28500 5108 28506 5160
rect 32766 5108 32772 5160
rect 32824 5148 32830 5160
rect 32950 5148 32956 5160
rect 32824 5120 32956 5148
rect 32824 5108 32830 5120
rect 32950 5108 32956 5120
rect 33008 5108 33014 5160
rect 34532 5148 34560 5256
rect 34606 5244 34612 5296
rect 34664 5284 34670 5296
rect 34977 5287 35035 5293
rect 34977 5284 34989 5287
rect 34664 5256 34989 5284
rect 34664 5244 34670 5256
rect 34977 5253 34989 5256
rect 35023 5253 35035 5287
rect 34977 5247 35035 5253
rect 35069 5287 35127 5293
rect 35069 5253 35081 5287
rect 35115 5284 35127 5287
rect 36538 5284 36544 5296
rect 35115 5256 36544 5284
rect 35115 5253 35127 5256
rect 35069 5247 35127 5253
rect 36538 5244 36544 5256
rect 36596 5244 36602 5296
rect 34790 5176 34796 5228
rect 34848 5216 34854 5228
rect 34885 5219 34943 5225
rect 34885 5216 34897 5219
rect 34848 5188 34897 5216
rect 34848 5176 34854 5188
rect 34885 5185 34897 5188
rect 34931 5185 34943 5219
rect 34885 5179 34943 5185
rect 35250 5176 35256 5228
rect 35308 5176 35314 5228
rect 37458 5148 37464 5160
rect 34532 5120 37464 5148
rect 37458 5108 37464 5120
rect 37516 5108 37522 5160
rect 21913 5083 21971 5089
rect 21913 5049 21925 5083
rect 21959 5080 21971 5083
rect 22370 5080 22376 5092
rect 21959 5052 22376 5080
rect 21959 5049 21971 5052
rect 21913 5043 21971 5049
rect 22370 5040 22376 5052
rect 22428 5040 22434 5092
rect 1104 4922 42504 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 42504 4922
rect 1104 4848 42504 4870
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 4856 4780 4905 4808
rect 4856 4768 4862 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 4893 4771 4951 4777
rect 5626 4768 5632 4820
rect 5684 4768 5690 4820
rect 7190 4768 7196 4820
rect 7248 4768 7254 4820
rect 8021 4811 8079 4817
rect 8021 4777 8033 4811
rect 8067 4808 8079 4811
rect 8110 4808 8116 4820
rect 8067 4780 8116 4808
rect 8067 4777 8079 4780
rect 8021 4771 8079 4777
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 32950 4768 32956 4820
rect 33008 4768 33014 4820
rect 5994 4740 6000 4752
rect 5552 4712 6000 4740
rect 5552 4681 5580 4712
rect 5994 4700 6000 4712
rect 6052 4740 6058 4752
rect 6181 4743 6239 4749
rect 6181 4740 6193 4743
rect 6052 4712 6193 4740
rect 6052 4700 6058 4712
rect 6181 4709 6193 4712
rect 6227 4709 6239 4743
rect 6181 4703 6239 4709
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4641 5595 4675
rect 5537 4635 5595 4641
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 8846 4672 8852 4684
rect 8527 4644 8852 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 31202 4632 31208 4684
rect 31260 4632 31266 4684
rect 31478 4632 31484 4684
rect 31536 4632 31542 4684
rect 5810 4564 5816 4616
rect 5868 4564 5874 4616
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 6638 4604 6644 4616
rect 5951 4576 6644 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 8386 4564 8392 4616
rect 8444 4564 8450 4616
rect 5997 4539 6055 4545
rect 5997 4505 6009 4539
rect 6043 4536 6055 4539
rect 6086 4536 6092 4548
rect 6043 4508 6092 4536
rect 6043 4505 6055 4508
rect 5997 4499 6055 4505
rect 6086 4496 6092 4508
rect 6144 4496 6150 4548
rect 7469 4539 7527 4545
rect 7469 4505 7481 4539
rect 7515 4536 7527 4539
rect 10502 4536 10508 4548
rect 7515 4508 10508 4536
rect 7515 4505 7527 4508
rect 7469 4499 7527 4505
rect 10502 4496 10508 4508
rect 10560 4496 10566 4548
rect 33042 4536 33048 4548
rect 32706 4508 33048 4536
rect 33042 4496 33048 4508
rect 33100 4496 33106 4548
rect 1104 4378 42504 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 42504 4378
rect 1104 4304 42504 4326
rect 1104 3834 42504 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 42504 3834
rect 1104 3760 42504 3782
rect 1104 3290 42504 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 42504 3290
rect 1104 3216 42504 3238
rect 1104 2746 42504 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 42504 2746
rect 1104 2672 42504 2694
rect 11422 2388 11428 2440
rect 11480 2428 11486 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11480 2400 11713 2428
rect 11480 2388 11486 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 1104 2202 42504 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 42504 2202
rect 1104 2128 42504 2150
<< via1 >>
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 35594 43494 35646 43546
rect 35658 43494 35710 43546
rect 35722 43494 35774 43546
rect 35786 43494 35838 43546
rect 35850 43494 35902 43546
rect 20260 43435 20312 43444
rect 20260 43401 20269 43435
rect 20269 43401 20303 43435
rect 20303 43401 20312 43435
rect 20260 43392 20312 43401
rect 20536 43392 20588 43444
rect 21548 43435 21600 43444
rect 21548 43401 21557 43435
rect 21557 43401 21591 43435
rect 21591 43401 21600 43435
rect 21548 43392 21600 43401
rect 22744 43435 22796 43444
rect 22744 43401 22753 43435
rect 22753 43401 22787 43435
rect 22787 43401 22796 43435
rect 22744 43392 22796 43401
rect 24032 43435 24084 43444
rect 24032 43401 24041 43435
rect 24041 43401 24075 43435
rect 24075 43401 24084 43435
rect 24032 43392 24084 43401
rect 19892 43256 19944 43308
rect 20904 43256 20956 43308
rect 21088 43299 21140 43308
rect 21088 43265 21097 43299
rect 21097 43265 21131 43299
rect 21131 43265 21140 43299
rect 21088 43256 21140 43265
rect 21640 43324 21692 43376
rect 21180 43188 21232 43240
rect 23112 43256 23164 43308
rect 23756 43256 23808 43308
rect 26240 43188 26292 43240
rect 33876 43188 33928 43240
rect 21548 43052 21600 43104
rect 25872 43095 25924 43104
rect 25872 43061 25881 43095
rect 25881 43061 25915 43095
rect 25915 43061 25924 43095
rect 25872 43052 25924 43061
rect 33784 43095 33836 43104
rect 33784 43061 33793 43095
rect 33793 43061 33827 43095
rect 33827 43061 33836 43095
rect 33784 43052 33836 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 33140 42848 33192 42900
rect 33876 42891 33928 42900
rect 33876 42857 33885 42891
rect 33885 42857 33919 42891
rect 33919 42857 33928 42891
rect 33876 42848 33928 42857
rect 17868 42780 17920 42832
rect 23572 42780 23624 42832
rect 29552 42755 29604 42764
rect 29552 42721 29561 42755
rect 29561 42721 29595 42755
rect 29595 42721 29604 42755
rect 29552 42712 29604 42721
rect 31760 42712 31812 42764
rect 34336 42712 34388 42764
rect 20168 42644 20220 42696
rect 21456 42687 21508 42696
rect 21456 42653 21465 42687
rect 21465 42653 21499 42687
rect 21499 42653 21508 42687
rect 21456 42644 21508 42653
rect 19432 42576 19484 42628
rect 23940 42644 23992 42696
rect 24676 42644 24728 42696
rect 25872 42644 25924 42696
rect 32128 42687 32180 42696
rect 32128 42653 32137 42687
rect 32137 42653 32171 42687
rect 32171 42653 32180 42687
rect 32128 42644 32180 42653
rect 33508 42644 33560 42696
rect 33968 42687 34020 42696
rect 33968 42653 33977 42687
rect 33977 42653 34011 42687
rect 34011 42653 34020 42687
rect 33968 42644 34020 42653
rect 22008 42619 22060 42628
rect 22008 42585 22017 42619
rect 22017 42585 22051 42619
rect 22051 42585 22060 42619
rect 22008 42576 22060 42585
rect 23296 42576 23348 42628
rect 27620 42576 27672 42628
rect 28724 42576 28776 42628
rect 29828 42619 29880 42628
rect 29828 42585 29837 42619
rect 29837 42585 29871 42619
rect 29871 42585 29880 42619
rect 29828 42576 29880 42585
rect 30472 42576 30524 42628
rect 19524 42508 19576 42560
rect 19616 42551 19668 42560
rect 19616 42517 19625 42551
rect 19625 42517 19659 42551
rect 19659 42517 19668 42551
rect 19616 42508 19668 42517
rect 19800 42508 19852 42560
rect 20444 42508 20496 42560
rect 23480 42551 23532 42560
rect 23480 42517 23489 42551
rect 23489 42517 23523 42551
rect 23523 42517 23532 42551
rect 23480 42508 23532 42517
rect 24584 42508 24636 42560
rect 25872 42508 25924 42560
rect 26056 42551 26108 42560
rect 26056 42517 26065 42551
rect 26065 42517 26099 42551
rect 26099 42517 26108 42551
rect 26056 42508 26108 42517
rect 26424 42551 26476 42560
rect 26424 42517 26433 42551
rect 26433 42517 26467 42551
rect 26467 42517 26476 42551
rect 26424 42508 26476 42517
rect 26792 42508 26844 42560
rect 29000 42508 29052 42560
rect 31392 42551 31444 42560
rect 31392 42517 31401 42551
rect 31401 42517 31435 42551
rect 31435 42517 31444 42551
rect 31392 42508 31444 42517
rect 33232 42508 33284 42560
rect 34060 42619 34112 42628
rect 34060 42585 34069 42619
rect 34069 42585 34103 42619
rect 34103 42585 34112 42619
rect 34060 42576 34112 42585
rect 34152 42576 34204 42628
rect 35348 42551 35400 42560
rect 35348 42517 35357 42551
rect 35357 42517 35391 42551
rect 35391 42517 35400 42551
rect 35348 42508 35400 42517
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 35594 42406 35646 42458
rect 35658 42406 35710 42458
rect 35722 42406 35774 42458
rect 35786 42406 35838 42458
rect 35850 42406 35902 42458
rect 21456 42304 21508 42356
rect 19800 42236 19852 42288
rect 20260 42236 20312 42288
rect 21088 42236 21140 42288
rect 19432 42211 19484 42220
rect 19432 42177 19441 42211
rect 19441 42177 19475 42211
rect 19475 42177 19484 42211
rect 19432 42168 19484 42177
rect 21640 42168 21692 42220
rect 23940 42236 23992 42288
rect 26240 42304 26292 42356
rect 26424 42304 26476 42356
rect 27620 42347 27672 42356
rect 27620 42313 27629 42347
rect 27629 42313 27663 42347
rect 27663 42313 27672 42347
rect 27620 42304 27672 42313
rect 29828 42304 29880 42356
rect 31392 42304 31444 42356
rect 31484 42304 31536 42356
rect 24584 42279 24636 42288
rect 24584 42245 24593 42279
rect 24593 42245 24627 42279
rect 24627 42245 24636 42279
rect 24584 42236 24636 42245
rect 26884 42236 26936 42288
rect 24308 42211 24360 42220
rect 24308 42177 24317 42211
rect 24317 42177 24351 42211
rect 24351 42177 24360 42211
rect 24308 42168 24360 42177
rect 25688 42168 25740 42220
rect 26700 42168 26752 42220
rect 29000 42211 29052 42220
rect 29000 42177 29009 42211
rect 29009 42177 29043 42211
rect 29043 42177 29052 42211
rect 29000 42168 29052 42177
rect 30840 42168 30892 42220
rect 31208 42211 31260 42220
rect 31208 42177 31217 42211
rect 31217 42177 31251 42211
rect 31251 42177 31260 42211
rect 31208 42168 31260 42177
rect 22468 42143 22520 42152
rect 22468 42109 22477 42143
rect 22477 42109 22511 42143
rect 22511 42109 22520 42143
rect 22468 42100 22520 42109
rect 26240 42143 26292 42152
rect 26240 42109 26249 42143
rect 26249 42109 26283 42143
rect 26283 42109 26292 42143
rect 26240 42100 26292 42109
rect 27712 42100 27764 42152
rect 27896 42032 27948 42084
rect 30104 42100 30156 42152
rect 31300 42100 31352 42152
rect 31576 42211 31628 42220
rect 31576 42177 31585 42211
rect 31585 42177 31619 42211
rect 31619 42177 31628 42211
rect 31576 42168 31628 42177
rect 31760 42211 31812 42220
rect 31760 42177 31769 42211
rect 31769 42177 31803 42211
rect 31803 42177 31812 42211
rect 31760 42168 31812 42177
rect 33140 42347 33192 42356
rect 33140 42313 33149 42347
rect 33149 42313 33183 42347
rect 33183 42313 33192 42347
rect 33140 42304 33192 42313
rect 33784 42304 33836 42356
rect 33968 42347 34020 42356
rect 33968 42313 33977 42347
rect 33977 42313 34011 42347
rect 34011 42313 34020 42347
rect 33968 42304 34020 42313
rect 34152 42236 34204 42288
rect 33876 42168 33928 42220
rect 34336 42168 34388 42220
rect 31852 42100 31904 42152
rect 33600 42143 33652 42152
rect 33600 42109 33609 42143
rect 33609 42109 33643 42143
rect 33643 42109 33652 42143
rect 33600 42100 33652 42109
rect 30656 42032 30708 42084
rect 34704 42100 34756 42152
rect 37464 42100 37516 42152
rect 38568 42100 38620 42152
rect 35992 42032 36044 42084
rect 21916 41964 21968 42016
rect 22560 41964 22612 42016
rect 24676 41964 24728 42016
rect 27068 42007 27120 42016
rect 27068 41973 27077 42007
rect 27077 41973 27111 42007
rect 27111 41973 27120 42007
rect 27068 41964 27120 41973
rect 31576 41964 31628 42016
rect 31852 41964 31904 42016
rect 37740 42007 37792 42016
rect 37740 41973 37749 42007
rect 37749 41973 37783 42007
rect 37783 41973 37792 42007
rect 37740 41964 37792 41973
rect 39488 42007 39540 42016
rect 39488 41973 39497 42007
rect 39497 41973 39531 42007
rect 39531 41973 39540 42007
rect 39488 41964 39540 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19616 41760 19668 41812
rect 22468 41760 22520 41812
rect 23940 41760 23992 41812
rect 25688 41760 25740 41812
rect 26240 41760 26292 41812
rect 28724 41760 28776 41812
rect 30472 41760 30524 41812
rect 31208 41760 31260 41812
rect 31484 41803 31536 41812
rect 31484 41769 31493 41803
rect 31493 41769 31527 41803
rect 31527 41769 31536 41803
rect 31484 41760 31536 41769
rect 34060 41803 34112 41812
rect 34060 41769 34069 41803
rect 34069 41769 34103 41803
rect 34103 41769 34112 41803
rect 34060 41760 34112 41769
rect 34704 41803 34756 41812
rect 34704 41769 34713 41803
rect 34713 41769 34747 41803
rect 34747 41769 34756 41803
rect 34704 41760 34756 41769
rect 19524 41667 19576 41676
rect 19524 41633 19533 41667
rect 19533 41633 19567 41667
rect 19567 41633 19576 41667
rect 19524 41624 19576 41633
rect 21088 41624 21140 41676
rect 21456 41624 21508 41676
rect 23572 41692 23624 41744
rect 24584 41692 24636 41744
rect 28080 41692 28132 41744
rect 29000 41692 29052 41744
rect 31116 41692 31168 41744
rect 31668 41692 31720 41744
rect 23480 41624 23532 41676
rect 23848 41624 23900 41676
rect 24308 41624 24360 41676
rect 26056 41624 26108 41676
rect 17132 41531 17184 41540
rect 17132 41497 17141 41531
rect 17141 41497 17175 41531
rect 17175 41497 17184 41531
rect 17132 41488 17184 41497
rect 21916 41599 21968 41608
rect 21916 41565 21925 41599
rect 21925 41565 21959 41599
rect 21959 41565 21968 41599
rect 21916 41556 21968 41565
rect 22560 41599 22612 41608
rect 22560 41565 22569 41599
rect 22569 41565 22603 41599
rect 22603 41565 22612 41599
rect 22560 41556 22612 41565
rect 23296 41556 23348 41608
rect 24400 41599 24452 41608
rect 24400 41565 24409 41599
rect 24409 41565 24443 41599
rect 24443 41565 24452 41599
rect 24400 41556 24452 41565
rect 24676 41599 24728 41608
rect 24676 41565 24685 41599
rect 24685 41565 24719 41599
rect 24719 41565 24728 41599
rect 24676 41556 24728 41565
rect 26884 41556 26936 41608
rect 18604 41463 18656 41472
rect 18604 41429 18613 41463
rect 18613 41429 18647 41463
rect 18647 41429 18656 41463
rect 18604 41420 18656 41429
rect 19432 41488 19484 41540
rect 19984 41488 20036 41540
rect 21548 41488 21600 41540
rect 22376 41488 22428 41540
rect 20260 41420 20312 41472
rect 21088 41420 21140 41472
rect 22560 41463 22612 41472
rect 22560 41429 22569 41463
rect 22569 41429 22603 41463
rect 22603 41429 22612 41463
rect 22560 41420 22612 41429
rect 22928 41488 22980 41540
rect 23572 41488 23624 41540
rect 25688 41488 25740 41540
rect 23480 41463 23532 41472
rect 23480 41429 23489 41463
rect 23489 41429 23523 41463
rect 23523 41429 23532 41463
rect 23480 41420 23532 41429
rect 24768 41420 24820 41472
rect 26700 41488 26752 41540
rect 28172 41599 28224 41608
rect 28172 41565 28181 41599
rect 28181 41565 28215 41599
rect 28215 41565 28224 41599
rect 29552 41624 29604 41676
rect 29736 41667 29788 41676
rect 29736 41633 29745 41667
rect 29745 41633 29779 41667
rect 29779 41633 29788 41667
rect 29736 41624 29788 41633
rect 31300 41624 31352 41676
rect 28172 41556 28224 41565
rect 29276 41556 29328 41608
rect 31484 41556 31536 41608
rect 31760 41624 31812 41676
rect 32864 41624 32916 41676
rect 33324 41624 33376 41676
rect 31852 41599 31904 41608
rect 31852 41565 31861 41599
rect 31861 41565 31895 41599
rect 31895 41565 31904 41599
rect 31852 41556 31904 41565
rect 26608 41463 26660 41472
rect 26608 41429 26617 41463
rect 26617 41429 26651 41463
rect 26651 41429 26660 41463
rect 26608 41420 26660 41429
rect 28632 41463 28684 41472
rect 28632 41429 28641 41463
rect 28641 41429 28675 41463
rect 28675 41429 28684 41463
rect 28632 41420 28684 41429
rect 29184 41531 29236 41540
rect 29184 41497 29193 41531
rect 29193 41497 29227 41531
rect 29227 41497 29236 41531
rect 29184 41488 29236 41497
rect 30012 41531 30064 41540
rect 30012 41497 30021 41531
rect 30021 41497 30055 41531
rect 30055 41497 30064 41531
rect 30012 41488 30064 41497
rect 30472 41488 30524 41540
rect 33232 41599 33284 41608
rect 33232 41565 33241 41599
rect 33241 41565 33275 41599
rect 33275 41565 33284 41599
rect 33232 41556 33284 41565
rect 33876 41624 33928 41676
rect 34428 41735 34480 41744
rect 34428 41701 34437 41735
rect 34437 41701 34471 41735
rect 34471 41701 34480 41735
rect 34428 41692 34480 41701
rect 33416 41488 33468 41540
rect 34152 41599 34204 41608
rect 34152 41565 34161 41599
rect 34161 41565 34195 41599
rect 34195 41565 34204 41599
rect 34152 41556 34204 41565
rect 38016 41624 38068 41676
rect 39028 41624 39080 41676
rect 37464 41599 37516 41608
rect 37464 41565 37473 41599
rect 37473 41565 37507 41599
rect 37507 41565 37516 41599
rect 37464 41556 37516 41565
rect 33968 41488 34020 41540
rect 35348 41488 35400 41540
rect 37648 41488 37700 41540
rect 37832 41488 37884 41540
rect 38108 41488 38160 41540
rect 39396 41531 39448 41540
rect 39396 41497 39405 41531
rect 39405 41497 39439 41531
rect 39439 41497 39448 41531
rect 39396 41488 39448 41497
rect 30840 41420 30892 41472
rect 31484 41420 31536 41472
rect 31668 41420 31720 41472
rect 32772 41463 32824 41472
rect 32772 41429 32781 41463
rect 32781 41429 32815 41463
rect 32815 41429 32824 41463
rect 32772 41420 32824 41429
rect 35164 41463 35216 41472
rect 35164 41429 35173 41463
rect 35173 41429 35207 41463
rect 35207 41429 35216 41463
rect 35164 41420 35216 41429
rect 37464 41463 37516 41472
rect 37464 41429 37473 41463
rect 37473 41429 37507 41463
rect 37507 41429 37516 41463
rect 37464 41420 37516 41429
rect 37924 41463 37976 41472
rect 37924 41429 37933 41463
rect 37933 41429 37967 41463
rect 37967 41429 37976 41463
rect 37924 41420 37976 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 35594 41318 35646 41370
rect 35658 41318 35710 41370
rect 35722 41318 35774 41370
rect 35786 41318 35838 41370
rect 35850 41318 35902 41370
rect 17132 41216 17184 41268
rect 17224 41148 17276 41200
rect 18604 41080 18656 41132
rect 18788 41080 18840 41132
rect 22008 41216 22060 41268
rect 23572 41216 23624 41268
rect 21088 41123 21140 41132
rect 16856 41055 16908 41064
rect 16856 41021 16865 41055
rect 16865 41021 16899 41055
rect 16899 41021 16908 41055
rect 16856 41012 16908 41021
rect 17776 41012 17828 41064
rect 18052 41055 18104 41064
rect 18052 41021 18061 41055
rect 18061 41021 18095 41055
rect 18095 41021 18104 41055
rect 18052 41012 18104 41021
rect 21088 41089 21096 41123
rect 21096 41089 21130 41123
rect 21130 41089 21140 41123
rect 21088 41080 21140 41089
rect 18880 40944 18932 40996
rect 20352 40987 20404 40996
rect 20352 40953 20361 40987
rect 20361 40953 20395 40987
rect 20395 40953 20404 40987
rect 20352 40944 20404 40953
rect 20536 40944 20588 40996
rect 20812 40987 20864 40996
rect 20812 40953 20821 40987
rect 20821 40953 20855 40987
rect 20855 40953 20864 40987
rect 20812 40944 20864 40953
rect 21272 40987 21324 40996
rect 21272 40953 21281 40987
rect 21281 40953 21315 40987
rect 21315 40953 21324 40987
rect 21272 40944 21324 40953
rect 21548 41123 21600 41132
rect 21548 41089 21557 41123
rect 21557 41089 21591 41123
rect 21591 41089 21600 41123
rect 21548 41080 21600 41089
rect 21640 41080 21692 41132
rect 23480 41080 23532 41132
rect 23848 41191 23900 41200
rect 23848 41157 23857 41191
rect 23857 41157 23891 41191
rect 23891 41157 23900 41191
rect 23848 41148 23900 41157
rect 26148 41216 26200 41268
rect 26240 41216 26292 41268
rect 28172 41216 28224 41268
rect 28264 41216 28316 41268
rect 28908 41216 28960 41268
rect 30840 41216 30892 41268
rect 31484 41216 31536 41268
rect 33600 41216 33652 41268
rect 35164 41259 35216 41268
rect 35164 41225 35173 41259
rect 35173 41225 35207 41259
rect 35207 41225 35216 41259
rect 35164 41216 35216 41225
rect 37740 41216 37792 41268
rect 39396 41216 39448 41268
rect 39488 41216 39540 41268
rect 21916 41012 21968 41064
rect 22744 41012 22796 41064
rect 23572 41012 23624 41064
rect 24768 41080 24820 41132
rect 21456 40944 21508 40996
rect 22376 40944 22428 40996
rect 24400 40944 24452 40996
rect 26240 41123 26292 41132
rect 26240 41089 26249 41123
rect 26249 41089 26283 41123
rect 26283 41089 26292 41123
rect 26240 41080 26292 41089
rect 26608 41080 26660 41132
rect 27804 41123 27856 41132
rect 27804 41089 27813 41123
rect 27813 41089 27847 41123
rect 27847 41089 27856 41123
rect 27804 41080 27856 41089
rect 29184 41148 29236 41200
rect 28080 41080 28132 41132
rect 28540 41123 28592 41132
rect 28540 41089 28549 41123
rect 28549 41089 28583 41123
rect 28583 41089 28592 41123
rect 28540 41080 28592 41089
rect 28356 41055 28408 41064
rect 28356 41021 28365 41055
rect 28365 41021 28399 41055
rect 28399 41021 28408 41055
rect 28356 41012 28408 41021
rect 27068 40944 27120 40996
rect 28264 40944 28316 40996
rect 28908 41080 28960 41132
rect 29092 41123 29144 41132
rect 29092 41089 29101 41123
rect 29101 41089 29135 41123
rect 29135 41089 29144 41123
rect 29092 41080 29144 41089
rect 29736 41080 29788 41132
rect 30932 41123 30984 41132
rect 30932 41089 30941 41123
rect 30941 41089 30975 41123
rect 30975 41089 30984 41123
rect 30932 41080 30984 41089
rect 31576 41123 31628 41132
rect 31576 41089 31585 41123
rect 31585 41089 31619 41123
rect 31619 41089 31628 41123
rect 31576 41080 31628 41089
rect 31760 41123 31812 41132
rect 31760 41089 31769 41123
rect 31769 41089 31803 41123
rect 31803 41089 31812 41123
rect 31760 41080 31812 41089
rect 32864 41148 32916 41200
rect 31116 40944 31168 40996
rect 33140 41123 33192 41132
rect 33140 41089 33149 41123
rect 33149 41089 33183 41123
rect 33183 41089 33192 41123
rect 33140 41080 33192 41089
rect 33232 41080 33284 41132
rect 33416 41080 33468 41132
rect 34796 41148 34848 41200
rect 37372 41148 37424 41200
rect 37556 41148 37608 41200
rect 37832 41148 37884 41200
rect 37924 41148 37976 41200
rect 33048 41012 33100 41064
rect 34428 41012 34480 41064
rect 35440 41080 35492 41132
rect 38568 41148 38620 41200
rect 33324 40944 33376 40996
rect 34704 40944 34756 40996
rect 37832 41055 37884 41064
rect 37832 41021 37841 41055
rect 37841 41021 37875 41055
rect 37875 41021 37884 41055
rect 37832 41012 37884 41021
rect 38292 41123 38344 41132
rect 38292 41089 38301 41123
rect 38301 41089 38335 41123
rect 38335 41089 38344 41123
rect 38292 41080 38344 41089
rect 39580 41080 39632 41132
rect 40224 41123 40276 41132
rect 40224 41089 40233 41123
rect 40233 41089 40267 41123
rect 40267 41089 40276 41123
rect 40224 41080 40276 41089
rect 38844 41055 38896 41064
rect 38844 41021 38853 41055
rect 38853 41021 38887 41055
rect 38887 41021 38896 41055
rect 38844 41012 38896 41021
rect 17040 40876 17092 40928
rect 21180 40876 21232 40928
rect 26056 40919 26108 40928
rect 26056 40885 26065 40919
rect 26065 40885 26099 40919
rect 26099 40885 26108 40919
rect 26056 40876 26108 40885
rect 26424 40919 26476 40928
rect 26424 40885 26433 40919
rect 26433 40885 26467 40919
rect 26467 40885 26476 40919
rect 26424 40876 26476 40885
rect 28448 40876 28500 40928
rect 28632 40876 28684 40928
rect 29276 40876 29328 40928
rect 30472 40876 30524 40928
rect 32588 40919 32640 40928
rect 32588 40885 32597 40919
rect 32597 40885 32631 40919
rect 32631 40885 32640 40919
rect 32588 40876 32640 40885
rect 36820 40919 36872 40928
rect 36820 40885 36829 40919
rect 36829 40885 36863 40919
rect 36863 40885 36872 40919
rect 36820 40876 36872 40885
rect 37188 40876 37240 40928
rect 37280 40919 37332 40928
rect 37280 40885 37289 40919
rect 37289 40885 37323 40919
rect 37323 40885 37332 40919
rect 37280 40876 37332 40885
rect 39304 41012 39356 41064
rect 40132 41012 40184 41064
rect 39856 40944 39908 40996
rect 37648 40876 37700 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 16856 40672 16908 40724
rect 17776 40715 17828 40724
rect 17776 40681 17785 40715
rect 17785 40681 17819 40715
rect 17819 40681 17828 40715
rect 17776 40672 17828 40681
rect 20352 40672 20404 40724
rect 20536 40604 20588 40656
rect 26056 40647 26108 40656
rect 26056 40613 26065 40647
rect 26065 40613 26099 40647
rect 26099 40613 26108 40647
rect 26056 40604 26108 40613
rect 17408 40536 17460 40588
rect 14740 40468 14792 40520
rect 18788 40511 18840 40520
rect 18788 40477 18797 40511
rect 18797 40477 18831 40511
rect 18831 40477 18840 40511
rect 18788 40468 18840 40477
rect 18880 40511 18932 40520
rect 18880 40477 18889 40511
rect 18889 40477 18923 40511
rect 18923 40477 18932 40511
rect 18880 40468 18932 40477
rect 24860 40536 24912 40588
rect 15660 40443 15712 40452
rect 15660 40409 15669 40443
rect 15669 40409 15703 40443
rect 15703 40409 15712 40443
rect 15660 40400 15712 40409
rect 16120 40400 16172 40452
rect 18696 40400 18748 40452
rect 17776 40332 17828 40384
rect 18236 40375 18288 40384
rect 18236 40341 18245 40375
rect 18245 40341 18279 40375
rect 18279 40341 18288 40375
rect 18236 40332 18288 40341
rect 18880 40332 18932 40384
rect 19524 40443 19576 40452
rect 19524 40409 19533 40443
rect 19533 40409 19567 40443
rect 19567 40409 19576 40443
rect 19524 40400 19576 40409
rect 19432 40332 19484 40384
rect 20352 40400 20404 40452
rect 20996 40511 21048 40520
rect 20996 40477 21005 40511
rect 21005 40477 21039 40511
rect 21039 40477 21048 40511
rect 20996 40468 21048 40477
rect 21272 40511 21324 40520
rect 21272 40477 21281 40511
rect 21281 40477 21315 40511
rect 21315 40477 21324 40511
rect 21272 40468 21324 40477
rect 22560 40468 22612 40520
rect 24584 40468 24636 40520
rect 25136 40511 25188 40520
rect 25136 40477 25145 40511
rect 25145 40477 25179 40511
rect 25179 40477 25188 40511
rect 25136 40468 25188 40477
rect 25412 40511 25464 40520
rect 25412 40477 25421 40511
rect 25421 40477 25455 40511
rect 25455 40477 25464 40511
rect 25412 40468 25464 40477
rect 26424 40511 26476 40520
rect 26424 40477 26433 40511
rect 26433 40477 26467 40511
rect 26467 40477 26476 40511
rect 27896 40672 27948 40724
rect 28172 40672 28224 40724
rect 28724 40647 28776 40656
rect 28724 40613 28733 40647
rect 28733 40613 28767 40647
rect 28767 40613 28776 40647
rect 28724 40604 28776 40613
rect 30012 40672 30064 40724
rect 31484 40672 31536 40724
rect 34704 40672 34756 40724
rect 37280 40672 37332 40724
rect 37372 40672 37424 40724
rect 38292 40672 38344 40724
rect 40040 40672 40092 40724
rect 40224 40672 40276 40724
rect 31116 40647 31168 40656
rect 31116 40613 31125 40647
rect 31125 40613 31159 40647
rect 31159 40613 31168 40647
rect 31116 40604 31168 40613
rect 33048 40647 33100 40656
rect 33048 40613 33057 40647
rect 33057 40613 33091 40647
rect 33091 40613 33100 40647
rect 33048 40604 33100 40613
rect 38016 40604 38068 40656
rect 40132 40604 40184 40656
rect 28540 40536 28592 40588
rect 26424 40468 26476 40477
rect 27804 40468 27856 40520
rect 27988 40511 28040 40520
rect 27988 40477 27996 40511
rect 27996 40477 28030 40511
rect 28030 40477 28040 40511
rect 27988 40468 28040 40477
rect 28080 40511 28132 40520
rect 28080 40477 28089 40511
rect 28089 40477 28123 40511
rect 28123 40477 28132 40511
rect 28080 40468 28132 40477
rect 28908 40468 28960 40520
rect 30656 40579 30708 40588
rect 30656 40545 30665 40579
rect 30665 40545 30699 40579
rect 30699 40545 30708 40579
rect 30656 40536 30708 40545
rect 31760 40536 31812 40588
rect 32864 40579 32916 40588
rect 32864 40545 32873 40579
rect 32873 40545 32907 40579
rect 32907 40545 32916 40579
rect 32864 40536 32916 40545
rect 35992 40579 36044 40588
rect 35992 40545 36001 40579
rect 36001 40545 36035 40579
rect 36035 40545 36044 40579
rect 35992 40536 36044 40545
rect 20720 40332 20772 40384
rect 22560 40375 22612 40384
rect 22560 40341 22569 40375
rect 22569 40341 22603 40375
rect 22603 40341 22612 40375
rect 22560 40332 22612 40341
rect 26056 40332 26108 40384
rect 27620 40332 27672 40384
rect 27896 40332 27948 40384
rect 28356 40332 28408 40384
rect 28908 40332 28960 40384
rect 30472 40511 30524 40520
rect 30472 40477 30481 40511
rect 30481 40477 30515 40511
rect 30515 40477 30524 40511
rect 30472 40468 30524 40477
rect 32772 40511 32824 40520
rect 32772 40477 32781 40511
rect 32781 40477 32815 40511
rect 32815 40477 32824 40511
rect 32772 40468 32824 40477
rect 33232 40511 33284 40520
rect 33232 40477 33271 40511
rect 33271 40477 33284 40511
rect 33232 40468 33284 40477
rect 33416 40511 33468 40520
rect 33416 40477 33425 40511
rect 33425 40477 33459 40511
rect 33459 40477 33468 40511
rect 33416 40468 33468 40477
rect 39212 40511 39264 40520
rect 39212 40477 39221 40511
rect 39221 40477 39255 40511
rect 39255 40477 39264 40511
rect 39212 40468 39264 40477
rect 38108 40400 38160 40452
rect 40132 40400 40184 40452
rect 30564 40375 30616 40384
rect 30564 40341 30573 40375
rect 30573 40341 30607 40375
rect 30607 40341 30616 40375
rect 30564 40332 30616 40341
rect 32404 40375 32456 40384
rect 32404 40341 32413 40375
rect 32413 40341 32447 40375
rect 32447 40341 32456 40375
rect 32404 40332 32456 40341
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 35594 40230 35646 40282
rect 35658 40230 35710 40282
rect 35722 40230 35774 40282
rect 35786 40230 35838 40282
rect 35850 40230 35902 40282
rect 15660 40128 15712 40180
rect 17040 40171 17092 40180
rect 17040 40137 17049 40171
rect 17049 40137 17083 40171
rect 17083 40137 17092 40171
rect 17040 40128 17092 40137
rect 18236 40128 18288 40180
rect 24400 40128 24452 40180
rect 27988 40128 28040 40180
rect 28540 40128 28592 40180
rect 32864 40128 32916 40180
rect 39304 40171 39356 40180
rect 39304 40137 39313 40171
rect 39313 40137 39347 40171
rect 39347 40137 39356 40171
rect 39304 40128 39356 40137
rect 39580 40128 39632 40180
rect 17776 40060 17828 40112
rect 18788 40060 18840 40112
rect 21180 40060 21232 40112
rect 19432 39992 19484 40044
rect 20720 40035 20772 40044
rect 20720 40001 20729 40035
rect 20729 40001 20763 40035
rect 20763 40001 20772 40035
rect 20720 39992 20772 40001
rect 23388 40103 23440 40112
rect 23388 40069 23397 40103
rect 23397 40069 23431 40103
rect 23431 40069 23440 40103
rect 23388 40060 23440 40069
rect 22100 39992 22152 40044
rect 24308 39992 24360 40044
rect 24584 40035 24636 40044
rect 24584 40001 24593 40035
rect 24593 40001 24627 40035
rect 24627 40001 24636 40035
rect 24584 39992 24636 40001
rect 24860 39992 24912 40044
rect 27620 40060 27672 40112
rect 17316 39967 17368 39976
rect 17316 39933 17325 39967
rect 17325 39933 17359 39967
rect 17359 39933 17368 39967
rect 17316 39924 17368 39933
rect 17868 39924 17920 39976
rect 17408 39856 17460 39908
rect 18880 39924 18932 39976
rect 20812 39967 20864 39976
rect 20812 39933 20821 39967
rect 20821 39933 20855 39967
rect 20855 39933 20864 39967
rect 20812 39924 20864 39933
rect 22560 39924 22612 39976
rect 23020 39967 23072 39976
rect 23020 39933 23029 39967
rect 23029 39933 23063 39967
rect 23063 39933 23072 39967
rect 23020 39924 23072 39933
rect 21088 39899 21140 39908
rect 21088 39865 21097 39899
rect 21097 39865 21131 39899
rect 21131 39865 21140 39899
rect 25228 39992 25280 40044
rect 32404 40103 32456 40112
rect 32404 40069 32413 40103
rect 32413 40069 32447 40103
rect 32447 40069 32456 40103
rect 32404 40060 32456 40069
rect 33140 40060 33192 40112
rect 31116 39992 31168 40044
rect 32036 39992 32088 40044
rect 36820 40060 36872 40112
rect 38292 40103 38344 40112
rect 38292 40069 38301 40103
rect 38301 40069 38335 40103
rect 38335 40069 38344 40103
rect 38292 40060 38344 40069
rect 38844 40060 38896 40112
rect 26056 39967 26108 39976
rect 26056 39933 26065 39967
rect 26065 39933 26099 39967
rect 26099 39933 26108 39967
rect 26056 39924 26108 39933
rect 26976 39924 27028 39976
rect 27896 39967 27948 39976
rect 27896 39933 27905 39967
rect 27905 39933 27939 39967
rect 27939 39933 27948 39967
rect 27896 39924 27948 39933
rect 21088 39856 21140 39865
rect 18788 39788 18840 39840
rect 22100 39788 22152 39840
rect 24768 39831 24820 39840
rect 24768 39797 24777 39831
rect 24777 39797 24811 39831
rect 24811 39797 24820 39831
rect 24768 39788 24820 39797
rect 25320 39856 25372 39908
rect 28356 39899 28408 39908
rect 28356 39865 28365 39899
rect 28365 39865 28399 39899
rect 28399 39865 28408 39899
rect 28356 39856 28408 39865
rect 32496 39856 32548 39908
rect 37464 39992 37516 40044
rect 39212 39924 39264 39976
rect 39856 39967 39908 39976
rect 39856 39933 39865 39967
rect 39865 39933 39899 39967
rect 39899 39933 39908 39967
rect 39856 39924 39908 39933
rect 32404 39831 32456 39840
rect 32404 39797 32413 39831
rect 32413 39797 32447 39831
rect 32447 39797 32456 39831
rect 32404 39788 32456 39797
rect 32680 39788 32732 39840
rect 35348 39788 35400 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 30104 39584 30156 39636
rect 30564 39584 30616 39636
rect 32036 39584 32088 39636
rect 32220 39584 32272 39636
rect 32588 39584 32640 39636
rect 33508 39584 33560 39636
rect 34888 39584 34940 39636
rect 35256 39584 35308 39636
rect 24584 39516 24636 39568
rect 31116 39516 31168 39568
rect 18788 39491 18840 39500
rect 18788 39457 18797 39491
rect 18797 39457 18831 39491
rect 18831 39457 18840 39491
rect 18788 39448 18840 39457
rect 22192 39448 22244 39500
rect 18696 39423 18748 39432
rect 18696 39389 18705 39423
rect 18705 39389 18739 39423
rect 18739 39389 18748 39423
rect 18696 39380 18748 39389
rect 22100 39380 22152 39432
rect 30840 39448 30892 39500
rect 31484 39491 31536 39500
rect 31484 39457 31493 39491
rect 31493 39457 31527 39491
rect 31527 39457 31536 39491
rect 31484 39448 31536 39457
rect 32036 39448 32088 39500
rect 32680 39491 32732 39500
rect 32680 39457 32689 39491
rect 32689 39457 32723 39491
rect 32723 39457 32732 39491
rect 32680 39448 32732 39457
rect 34612 39516 34664 39568
rect 21824 39312 21876 39364
rect 24308 39380 24360 39432
rect 24768 39423 24820 39432
rect 24768 39389 24777 39423
rect 24777 39389 24811 39423
rect 24811 39389 24820 39423
rect 24768 39380 24820 39389
rect 25228 39423 25280 39432
rect 25228 39389 25237 39423
rect 25237 39389 25271 39423
rect 25271 39389 25280 39423
rect 25228 39380 25280 39389
rect 25320 39423 25372 39432
rect 25320 39389 25330 39423
rect 25330 39389 25364 39423
rect 25364 39389 25372 39423
rect 25320 39380 25372 39389
rect 31852 39380 31904 39432
rect 32220 39380 32272 39432
rect 32312 39380 32364 39432
rect 30932 39312 30984 39364
rect 31944 39355 31996 39364
rect 31944 39321 31953 39355
rect 31953 39321 31987 39355
rect 31987 39321 31996 39355
rect 32588 39423 32640 39432
rect 32588 39389 32597 39423
rect 32597 39389 32631 39423
rect 32631 39389 32640 39423
rect 32588 39380 32640 39389
rect 31944 39312 31996 39321
rect 19708 39244 19760 39296
rect 22652 39244 22704 39296
rect 25596 39244 25648 39296
rect 30564 39244 30616 39296
rect 32220 39287 32272 39296
rect 32220 39253 32229 39287
rect 32229 39253 32263 39287
rect 32263 39253 32272 39287
rect 32220 39244 32272 39253
rect 34244 39423 34296 39432
rect 34244 39389 34253 39423
rect 34253 39389 34287 39423
rect 34287 39389 34296 39423
rect 34244 39380 34296 39389
rect 34520 39355 34572 39364
rect 34520 39321 34529 39355
rect 34529 39321 34563 39355
rect 34563 39321 34572 39355
rect 34520 39312 34572 39321
rect 34796 39380 34848 39432
rect 35348 39448 35400 39500
rect 38568 39516 38620 39568
rect 40224 39448 40276 39500
rect 35164 39312 35216 39364
rect 36820 39380 36872 39432
rect 36636 39312 36688 39364
rect 37372 39380 37424 39432
rect 39672 39423 39724 39432
rect 39672 39389 39681 39423
rect 39681 39389 39715 39423
rect 39715 39389 39724 39423
rect 39672 39380 39724 39389
rect 38200 39312 38252 39364
rect 39396 39355 39448 39364
rect 39396 39321 39405 39355
rect 39405 39321 39439 39355
rect 39439 39321 39448 39355
rect 40960 39380 41012 39432
rect 42156 39423 42208 39432
rect 42156 39389 42165 39423
rect 42165 39389 42199 39423
rect 42199 39389 42208 39423
rect 42156 39380 42208 39389
rect 39396 39312 39448 39321
rect 34336 39244 34388 39296
rect 34428 39244 34480 39296
rect 35440 39287 35492 39296
rect 35440 39253 35449 39287
rect 35449 39253 35483 39287
rect 35483 39253 35492 39287
rect 35440 39244 35492 39253
rect 37648 39244 37700 39296
rect 39580 39287 39632 39296
rect 39580 39253 39589 39287
rect 39589 39253 39623 39287
rect 39623 39253 39632 39287
rect 39580 39244 39632 39253
rect 39764 39244 39816 39296
rect 40316 39287 40368 39296
rect 40316 39253 40325 39287
rect 40325 39253 40359 39287
rect 40359 39253 40368 39287
rect 40316 39244 40368 39253
rect 41420 39244 41472 39296
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 17224 39040 17276 39092
rect 18696 39040 18748 39092
rect 16580 38972 16632 39024
rect 14740 38947 14792 38956
rect 14740 38913 14749 38947
rect 14749 38913 14783 38947
rect 14783 38913 14792 38947
rect 14740 38904 14792 38913
rect 16120 38904 16172 38956
rect 20260 39015 20312 39024
rect 16488 38836 16540 38888
rect 17592 38743 17644 38752
rect 17592 38709 17601 38743
rect 17601 38709 17635 38743
rect 17635 38709 17644 38743
rect 17592 38700 17644 38709
rect 18420 38700 18472 38752
rect 19708 38947 19760 38956
rect 19708 38913 19718 38947
rect 19718 38913 19752 38947
rect 19752 38913 19760 38947
rect 20260 38981 20271 39015
rect 20271 38981 20312 39015
rect 20260 38972 20312 38981
rect 20352 38972 20404 39024
rect 21088 38972 21140 39024
rect 22100 39015 22152 39024
rect 22100 38981 22109 39015
rect 22109 38981 22143 39015
rect 22143 38981 22152 39015
rect 22100 38972 22152 38981
rect 19708 38904 19760 38913
rect 20812 38947 20864 38956
rect 20812 38913 20821 38947
rect 20821 38913 20855 38947
rect 20855 38913 20864 38947
rect 20812 38904 20864 38913
rect 21456 38947 21508 38956
rect 21456 38913 21465 38947
rect 21465 38913 21499 38947
rect 21499 38913 21508 38947
rect 21456 38904 21508 38913
rect 21824 38947 21876 38956
rect 21824 38913 21833 38947
rect 21833 38913 21867 38947
rect 21867 38913 21876 38947
rect 21824 38904 21876 38913
rect 23480 39040 23532 39092
rect 24308 39040 24360 39092
rect 25320 39040 25372 39092
rect 23940 38972 23992 39024
rect 24860 38904 24912 38956
rect 19340 38768 19392 38820
rect 20628 38811 20680 38820
rect 20628 38777 20637 38811
rect 20637 38777 20671 38811
rect 20671 38777 20680 38811
rect 20628 38768 20680 38777
rect 20076 38743 20128 38752
rect 20076 38709 20085 38743
rect 20085 38709 20119 38743
rect 20119 38709 20128 38743
rect 20076 38700 20128 38709
rect 20536 38700 20588 38752
rect 22468 38879 22520 38888
rect 22468 38845 22477 38879
rect 22477 38845 22511 38879
rect 22511 38845 22520 38879
rect 22468 38836 22520 38845
rect 25044 38947 25096 38956
rect 25044 38913 25053 38947
rect 25053 38913 25087 38947
rect 25087 38913 25096 38947
rect 25044 38904 25096 38913
rect 25596 39015 25648 39024
rect 25596 38981 25605 39015
rect 25605 38981 25639 39015
rect 25639 38981 25648 39015
rect 25596 38972 25648 38981
rect 25320 38904 25372 38956
rect 25412 38947 25464 38956
rect 25412 38913 25421 38947
rect 25421 38913 25455 38947
rect 25455 38913 25464 38947
rect 25412 38904 25464 38913
rect 28540 39040 28592 39092
rect 28724 38972 28776 39024
rect 24124 38768 24176 38820
rect 25228 38768 25280 38820
rect 22560 38700 22612 38752
rect 24032 38743 24084 38752
rect 24032 38709 24041 38743
rect 24041 38709 24075 38743
rect 24075 38709 24084 38743
rect 24032 38700 24084 38709
rect 24400 38700 24452 38752
rect 28356 38947 28408 38956
rect 28356 38913 28365 38947
rect 28365 38913 28399 38947
rect 28399 38913 28408 38947
rect 28356 38904 28408 38913
rect 31944 39040 31996 39092
rect 32128 39040 32180 39092
rect 33968 39040 34020 39092
rect 36176 39040 36228 39092
rect 28816 38836 28868 38888
rect 31392 38904 31444 38956
rect 31852 38836 31904 38888
rect 26700 38700 26752 38752
rect 26976 38700 27028 38752
rect 28448 38743 28500 38752
rect 28448 38709 28457 38743
rect 28457 38709 28491 38743
rect 28491 38709 28500 38743
rect 28448 38700 28500 38709
rect 28724 38700 28776 38752
rect 30380 38700 30432 38752
rect 31116 38743 31168 38752
rect 31116 38709 31125 38743
rect 31125 38709 31159 38743
rect 31159 38709 31168 38743
rect 31116 38700 31168 38709
rect 31944 38700 31996 38752
rect 32128 38947 32180 38956
rect 32128 38913 32137 38947
rect 32137 38913 32171 38947
rect 32171 38913 32180 38947
rect 32128 38904 32180 38913
rect 33508 38904 33560 38956
rect 32128 38768 32180 38820
rect 34888 38972 34940 39024
rect 33968 38947 34020 38956
rect 33968 38913 33977 38947
rect 33977 38913 34011 38947
rect 34011 38913 34020 38947
rect 33968 38904 34020 38913
rect 40224 39040 40276 39092
rect 38568 38972 38620 39024
rect 34612 38836 34664 38888
rect 35256 38836 35308 38888
rect 36636 38947 36688 38956
rect 36636 38913 36645 38947
rect 36645 38913 36679 38947
rect 36679 38913 36688 38947
rect 36636 38904 36688 38913
rect 37648 38947 37700 38956
rect 37648 38913 37657 38947
rect 37657 38913 37691 38947
rect 37691 38913 37700 38947
rect 37648 38904 37700 38913
rect 38108 38947 38160 38956
rect 38108 38913 38117 38947
rect 38117 38913 38151 38947
rect 38151 38913 38160 38947
rect 38108 38904 38160 38913
rect 38200 38947 38252 38956
rect 38200 38913 38209 38947
rect 38209 38913 38243 38947
rect 38243 38913 38252 38947
rect 38200 38904 38252 38913
rect 38384 38947 38436 38956
rect 38384 38913 38393 38947
rect 38393 38913 38427 38947
rect 38427 38913 38436 38947
rect 39764 38972 39816 39024
rect 40132 38972 40184 39024
rect 40960 39083 41012 39092
rect 40960 39049 40969 39083
rect 40969 39049 41003 39083
rect 41003 39049 41012 39083
rect 40960 39040 41012 39049
rect 41420 39083 41472 39092
rect 41420 39049 41429 39083
rect 41429 39049 41463 39083
rect 41463 39049 41472 39083
rect 41420 39040 41472 39049
rect 41236 38972 41288 39024
rect 38384 38904 38436 38913
rect 35716 38811 35768 38820
rect 35716 38777 35725 38811
rect 35725 38777 35759 38811
rect 35759 38777 35768 38811
rect 35716 38768 35768 38777
rect 39212 38879 39264 38888
rect 39212 38845 39221 38879
rect 39221 38845 39255 38879
rect 39255 38845 39264 38879
rect 39212 38836 39264 38845
rect 41328 38836 41380 38888
rect 37372 38768 37424 38820
rect 38016 38768 38068 38820
rect 33876 38743 33928 38752
rect 33876 38709 33885 38743
rect 33885 38709 33919 38743
rect 33919 38709 33928 38743
rect 33876 38700 33928 38709
rect 34428 38700 34480 38752
rect 34888 38700 34940 38752
rect 35624 38700 35676 38752
rect 35992 38700 36044 38752
rect 37832 38700 37884 38752
rect 41052 38743 41104 38752
rect 41052 38709 41061 38743
rect 41061 38709 41095 38743
rect 41095 38709 41104 38743
rect 41052 38700 41104 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 16488 38496 16540 38548
rect 17408 38496 17460 38548
rect 20996 38496 21048 38548
rect 21456 38496 21508 38548
rect 16580 38471 16632 38480
rect 16580 38437 16589 38471
rect 16589 38437 16623 38471
rect 16623 38437 16632 38471
rect 16580 38428 16632 38437
rect 21272 38428 21324 38480
rect 22468 38539 22520 38548
rect 22468 38505 22477 38539
rect 22477 38505 22511 38539
rect 22511 38505 22520 38539
rect 22468 38496 22520 38505
rect 24860 38539 24912 38548
rect 24860 38505 24869 38539
rect 24869 38505 24903 38539
rect 24903 38505 24912 38539
rect 24860 38496 24912 38505
rect 25320 38496 25372 38548
rect 17316 38403 17368 38412
rect 17316 38369 17325 38403
rect 17325 38369 17359 38403
rect 17359 38369 17368 38403
rect 17316 38360 17368 38369
rect 20076 38360 20128 38412
rect 14832 38335 14884 38344
rect 14832 38301 14841 38335
rect 14841 38301 14875 38335
rect 14875 38301 14884 38335
rect 14832 38292 14884 38301
rect 17500 38335 17552 38344
rect 17500 38301 17509 38335
rect 17509 38301 17543 38335
rect 17543 38301 17552 38335
rect 17500 38292 17552 38301
rect 19340 38292 19392 38344
rect 21088 38360 21140 38412
rect 20536 38335 20588 38344
rect 20536 38301 20545 38335
rect 20545 38301 20579 38335
rect 20579 38301 20588 38335
rect 20536 38292 20588 38301
rect 15108 38267 15160 38276
rect 15108 38233 15117 38267
rect 15117 38233 15151 38267
rect 15151 38233 15160 38267
rect 15108 38224 15160 38233
rect 16120 38224 16172 38276
rect 17592 38224 17644 38276
rect 18144 38224 18196 38276
rect 18788 38267 18840 38276
rect 18788 38233 18797 38267
rect 18797 38233 18831 38267
rect 18831 38233 18840 38267
rect 18788 38224 18840 38233
rect 20260 38267 20312 38276
rect 20260 38233 20269 38267
rect 20269 38233 20303 38267
rect 20303 38233 20312 38267
rect 20260 38224 20312 38233
rect 20352 38224 20404 38276
rect 17132 38199 17184 38208
rect 17132 38165 17141 38199
rect 17141 38165 17175 38199
rect 17175 38165 17184 38199
rect 17132 38156 17184 38165
rect 17684 38199 17736 38208
rect 17684 38165 17693 38199
rect 17693 38165 17727 38199
rect 17727 38165 17736 38199
rect 17684 38156 17736 38165
rect 19064 38156 19116 38208
rect 19708 38156 19760 38208
rect 20720 38224 20772 38276
rect 21456 38292 21508 38344
rect 21916 38292 21968 38344
rect 23020 38428 23072 38480
rect 31852 38496 31904 38548
rect 32128 38539 32180 38548
rect 32128 38505 32137 38539
rect 32137 38505 32171 38539
rect 32171 38505 32180 38539
rect 32128 38496 32180 38505
rect 34244 38496 34296 38548
rect 34796 38496 34848 38548
rect 39580 38496 39632 38548
rect 40132 38496 40184 38548
rect 41144 38496 41196 38548
rect 41420 38496 41472 38548
rect 42156 38539 42208 38548
rect 42156 38505 42165 38539
rect 42165 38505 42199 38539
rect 42199 38505 42208 38539
rect 42156 38496 42208 38505
rect 22652 38403 22704 38412
rect 22652 38369 22661 38403
rect 22661 38369 22695 38403
rect 22695 38369 22704 38403
rect 22652 38360 22704 38369
rect 24032 38360 24084 38412
rect 22560 38292 22612 38344
rect 22836 38292 22888 38344
rect 24400 38335 24452 38344
rect 24400 38301 24409 38335
rect 24409 38301 24443 38335
rect 24443 38301 24452 38335
rect 24400 38292 24452 38301
rect 24584 38335 24636 38344
rect 24584 38301 24593 38335
rect 24593 38301 24627 38335
rect 24627 38301 24636 38335
rect 24584 38292 24636 38301
rect 25596 38360 25648 38412
rect 25044 38292 25096 38344
rect 27252 38428 27304 38480
rect 27528 38403 27580 38412
rect 27528 38369 27537 38403
rect 27537 38369 27571 38403
rect 27571 38369 27580 38403
rect 27528 38360 27580 38369
rect 28356 38360 28408 38412
rect 28632 38403 28684 38412
rect 28632 38369 28641 38403
rect 28641 38369 28675 38403
rect 28675 38369 28684 38403
rect 28632 38360 28684 38369
rect 20996 38156 21048 38208
rect 21180 38156 21232 38208
rect 23020 38267 23072 38276
rect 23020 38233 23029 38267
rect 23029 38233 23063 38267
rect 23063 38233 23072 38267
rect 23020 38224 23072 38233
rect 26700 38335 26752 38344
rect 26700 38301 26709 38335
rect 26709 38301 26743 38335
rect 26743 38301 26752 38335
rect 26700 38292 26752 38301
rect 26976 38335 27028 38344
rect 26976 38301 26985 38335
rect 26985 38301 27019 38335
rect 27019 38301 27028 38335
rect 26976 38292 27028 38301
rect 25688 38267 25740 38276
rect 25688 38233 25697 38267
rect 25697 38233 25731 38267
rect 25731 38233 25740 38267
rect 25688 38224 25740 38233
rect 28264 38292 28316 38344
rect 28448 38292 28500 38344
rect 28816 38224 28868 38276
rect 34520 38428 34572 38480
rect 35072 38428 35124 38480
rect 38200 38471 38252 38480
rect 38200 38437 38209 38471
rect 38209 38437 38243 38471
rect 38243 38437 38252 38471
rect 38200 38428 38252 38437
rect 38384 38428 38436 38480
rect 32220 38360 32272 38412
rect 32680 38403 32732 38412
rect 32680 38369 32689 38403
rect 32689 38369 32723 38403
rect 32723 38369 32732 38403
rect 32680 38360 32732 38369
rect 33968 38360 34020 38412
rect 32404 38335 32456 38344
rect 32404 38301 32413 38335
rect 32413 38301 32447 38335
rect 32447 38301 32456 38335
rect 32404 38292 32456 38301
rect 33876 38292 33928 38344
rect 34244 38292 34296 38344
rect 34336 38267 34388 38276
rect 34336 38233 34345 38267
rect 34345 38233 34379 38267
rect 34379 38233 34388 38267
rect 34336 38224 34388 38233
rect 34612 38224 34664 38276
rect 34796 38335 34848 38344
rect 34796 38301 34805 38335
rect 34805 38301 34839 38335
rect 34839 38301 34848 38335
rect 34796 38292 34848 38301
rect 34888 38335 34940 38344
rect 34888 38301 34897 38335
rect 34897 38301 34931 38335
rect 34931 38301 34940 38335
rect 34888 38292 34940 38301
rect 35072 38335 35124 38344
rect 35072 38301 35081 38335
rect 35081 38301 35115 38335
rect 35115 38301 35124 38335
rect 35072 38292 35124 38301
rect 38016 38360 38068 38412
rect 37740 38335 37792 38344
rect 37740 38301 37749 38335
rect 37749 38301 37783 38335
rect 37783 38301 37792 38335
rect 37740 38292 37792 38301
rect 38108 38335 38160 38344
rect 38108 38301 38117 38335
rect 38117 38301 38151 38335
rect 38151 38301 38160 38335
rect 38108 38292 38160 38301
rect 39212 38360 39264 38412
rect 41052 38360 41104 38412
rect 38660 38292 38712 38344
rect 39396 38335 39448 38344
rect 39396 38301 39405 38335
rect 39405 38301 39439 38335
rect 39439 38301 39448 38335
rect 39396 38292 39448 38301
rect 39580 38292 39632 38344
rect 39672 38335 39724 38344
rect 39672 38301 39681 38335
rect 39681 38301 39715 38335
rect 39715 38301 39724 38335
rect 39672 38292 39724 38301
rect 40040 38335 40092 38344
rect 40040 38301 40049 38335
rect 40049 38301 40083 38335
rect 40083 38301 40092 38335
rect 40040 38292 40092 38301
rect 24584 38156 24636 38208
rect 25596 38199 25648 38208
rect 25596 38165 25605 38199
rect 25605 38165 25639 38199
rect 25639 38165 25648 38199
rect 25596 38156 25648 38165
rect 27160 38156 27212 38208
rect 28448 38199 28500 38208
rect 28448 38165 28457 38199
rect 28457 38165 28491 38199
rect 28491 38165 28500 38199
rect 28448 38156 28500 38165
rect 29552 38156 29604 38208
rect 31944 38156 31996 38208
rect 32588 38156 32640 38208
rect 34888 38156 34940 38208
rect 35440 38156 35492 38208
rect 35716 38224 35768 38276
rect 37188 38199 37240 38208
rect 37188 38165 37197 38199
rect 37197 38165 37231 38199
rect 37231 38165 37240 38199
rect 37188 38156 37240 38165
rect 37924 38199 37976 38208
rect 37924 38165 37933 38199
rect 37933 38165 37967 38199
rect 37967 38165 37976 38199
rect 37924 38156 37976 38165
rect 40132 38156 40184 38208
rect 41144 38224 41196 38276
rect 42156 38156 42208 38208
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 15108 37952 15160 38004
rect 17684 37952 17736 38004
rect 15752 37816 15804 37868
rect 16028 37816 16080 37868
rect 16212 37816 16264 37868
rect 13360 37791 13412 37800
rect 13360 37757 13369 37791
rect 13369 37757 13403 37791
rect 13403 37757 13412 37791
rect 13360 37748 13412 37757
rect 13636 37791 13688 37800
rect 13636 37757 13645 37791
rect 13645 37757 13679 37791
rect 13679 37757 13688 37791
rect 16856 37884 16908 37936
rect 17316 37884 17368 37936
rect 17408 37927 17460 37936
rect 17408 37893 17417 37927
rect 17417 37893 17451 37927
rect 17451 37893 17460 37927
rect 17408 37884 17460 37893
rect 18420 37927 18472 37936
rect 18420 37893 18429 37927
rect 18429 37893 18463 37927
rect 18463 37893 18472 37927
rect 18420 37884 18472 37893
rect 19064 37927 19116 37936
rect 19064 37893 19073 37927
rect 19073 37893 19107 37927
rect 19107 37893 19116 37927
rect 19064 37884 19116 37893
rect 20628 37884 20680 37936
rect 21916 37884 21968 37936
rect 28264 37995 28316 38004
rect 28264 37961 28273 37995
rect 28273 37961 28307 37995
rect 28307 37961 28316 37995
rect 28264 37952 28316 37961
rect 29552 37995 29604 38004
rect 29552 37961 29561 37995
rect 29561 37961 29595 37995
rect 29595 37961 29604 37995
rect 29552 37952 29604 37961
rect 35440 37952 35492 38004
rect 37188 37952 37240 38004
rect 39672 37952 39724 38004
rect 40316 37995 40368 38004
rect 40316 37961 40325 37995
rect 40325 37961 40359 37995
rect 40359 37961 40368 37995
rect 40316 37952 40368 37961
rect 41328 37952 41380 38004
rect 26424 37884 26476 37936
rect 18328 37859 18380 37868
rect 18328 37825 18337 37859
rect 18337 37825 18371 37859
rect 18371 37825 18380 37859
rect 18328 37816 18380 37825
rect 13636 37748 13688 37757
rect 16580 37748 16632 37800
rect 18144 37748 18196 37800
rect 18696 37680 18748 37732
rect 17592 37612 17644 37664
rect 20076 37748 20128 37800
rect 20536 37816 20588 37868
rect 20996 37816 21048 37868
rect 21180 37859 21232 37868
rect 21180 37825 21189 37859
rect 21189 37825 21223 37859
rect 21223 37825 21232 37859
rect 21180 37816 21232 37825
rect 21272 37859 21324 37868
rect 21272 37825 21281 37859
rect 21281 37825 21315 37859
rect 21315 37825 21324 37859
rect 21272 37816 21324 37825
rect 25504 37816 25556 37868
rect 27160 37859 27212 37868
rect 27160 37825 27169 37859
rect 27169 37825 27203 37859
rect 27203 37825 27212 37859
rect 27160 37816 27212 37825
rect 27252 37859 27304 37868
rect 27252 37825 27261 37859
rect 27261 37825 27295 37859
rect 27295 37825 27304 37859
rect 27252 37816 27304 37825
rect 21456 37748 21508 37800
rect 23020 37791 23072 37800
rect 23020 37757 23029 37791
rect 23029 37757 23063 37791
rect 23063 37757 23072 37791
rect 23020 37748 23072 37757
rect 34796 37884 34848 37936
rect 40868 37884 40920 37936
rect 20812 37680 20864 37732
rect 27896 37748 27948 37800
rect 19432 37612 19484 37664
rect 20536 37655 20588 37664
rect 20536 37621 20545 37655
rect 20545 37621 20579 37655
rect 20579 37621 20588 37655
rect 20536 37612 20588 37621
rect 20904 37612 20956 37664
rect 23664 37612 23716 37664
rect 24768 37612 24820 37664
rect 26516 37612 26568 37664
rect 27620 37612 27672 37664
rect 28540 37859 28592 37868
rect 28540 37825 28549 37859
rect 28549 37825 28583 37859
rect 28583 37825 28592 37859
rect 28540 37816 28592 37825
rect 33968 37816 34020 37868
rect 35992 37816 36044 37868
rect 37832 37859 37884 37868
rect 37832 37825 37841 37859
rect 37841 37825 37875 37859
rect 37875 37825 37884 37859
rect 37832 37816 37884 37825
rect 40040 37816 40092 37868
rect 40132 37859 40184 37868
rect 40132 37825 40141 37859
rect 40141 37825 40175 37859
rect 40175 37825 40184 37859
rect 40132 37816 40184 37825
rect 41144 37816 41196 37868
rect 28816 37748 28868 37800
rect 29000 37748 29052 37800
rect 30472 37791 30524 37800
rect 30472 37757 30481 37791
rect 30481 37757 30515 37791
rect 30515 37757 30524 37791
rect 30472 37748 30524 37757
rect 34152 37748 34204 37800
rect 38568 37791 38620 37800
rect 38568 37757 38577 37791
rect 38577 37757 38611 37791
rect 38611 37757 38620 37791
rect 38568 37748 38620 37757
rect 39856 37748 39908 37800
rect 41696 37791 41748 37800
rect 41696 37757 41705 37791
rect 41705 37757 41739 37791
rect 41739 37757 41748 37791
rect 41696 37748 41748 37757
rect 28632 37680 28684 37732
rect 30748 37680 30800 37732
rect 35072 37680 35124 37732
rect 38660 37680 38712 37732
rect 28816 37612 28868 37664
rect 33600 37612 33652 37664
rect 35256 37612 35308 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16212 37451 16264 37460
rect 16212 37417 16221 37451
rect 16221 37417 16255 37451
rect 16255 37417 16264 37451
rect 16212 37408 16264 37417
rect 17132 37408 17184 37460
rect 17408 37408 17460 37460
rect 18328 37408 18380 37460
rect 22468 37408 22520 37460
rect 23020 37408 23072 37460
rect 19524 37340 19576 37392
rect 19984 37340 20036 37392
rect 17592 37315 17644 37324
rect 17592 37281 17601 37315
rect 17601 37281 17635 37315
rect 17635 37281 17644 37315
rect 17592 37272 17644 37281
rect 19432 37272 19484 37324
rect 20904 37315 20956 37324
rect 20904 37281 20913 37315
rect 20913 37281 20947 37315
rect 20947 37281 20956 37315
rect 20904 37272 20956 37281
rect 23020 37315 23072 37324
rect 23020 37281 23029 37315
rect 23029 37281 23063 37315
rect 23063 37281 23072 37315
rect 23020 37272 23072 37281
rect 24768 37272 24820 37324
rect 24860 37315 24912 37324
rect 24860 37281 24869 37315
rect 24869 37281 24903 37315
rect 24903 37281 24912 37315
rect 24860 37272 24912 37281
rect 27068 37408 27120 37460
rect 12900 37204 12952 37256
rect 13360 37204 13412 37256
rect 14832 37247 14884 37256
rect 14832 37213 14841 37247
rect 14841 37213 14875 37247
rect 14875 37213 14884 37247
rect 14832 37204 14884 37213
rect 16580 37204 16632 37256
rect 17132 37204 17184 37256
rect 19524 37204 19576 37256
rect 20168 37204 20220 37256
rect 26516 37315 26568 37324
rect 26516 37281 26525 37315
rect 26525 37281 26559 37315
rect 26559 37281 26568 37315
rect 26516 37272 26568 37281
rect 32036 37315 32088 37324
rect 32036 37281 32045 37315
rect 32045 37281 32079 37315
rect 32079 37281 32088 37315
rect 32036 37272 32088 37281
rect 33692 37315 33744 37324
rect 33692 37281 33701 37315
rect 33701 37281 33735 37315
rect 33735 37281 33744 37315
rect 33692 37272 33744 37281
rect 33968 37272 34020 37324
rect 34152 37315 34204 37324
rect 34152 37281 34161 37315
rect 34161 37281 34195 37315
rect 34195 37281 34204 37315
rect 34152 37272 34204 37281
rect 34796 37272 34848 37324
rect 15108 37136 15160 37188
rect 20076 37136 20128 37188
rect 16028 37068 16080 37120
rect 19524 37068 19576 37120
rect 19892 37068 19944 37120
rect 25044 37204 25096 37256
rect 25688 37204 25740 37256
rect 27620 37204 27672 37256
rect 30656 37204 30708 37256
rect 31116 37204 31168 37256
rect 31208 37204 31260 37256
rect 31484 37247 31536 37256
rect 31484 37213 31493 37247
rect 31493 37213 31527 37247
rect 31527 37213 31536 37247
rect 31484 37204 31536 37213
rect 34980 37204 35032 37256
rect 20812 37136 20864 37188
rect 21456 37136 21508 37188
rect 20720 37068 20772 37120
rect 23020 37068 23072 37120
rect 23204 37111 23256 37120
rect 23204 37077 23213 37111
rect 23213 37077 23247 37111
rect 23247 37077 23256 37111
rect 23204 37068 23256 37077
rect 23388 37068 23440 37120
rect 23664 37068 23716 37120
rect 30380 37136 30432 37188
rect 31760 37136 31812 37188
rect 32772 37136 32824 37188
rect 33968 37179 34020 37188
rect 33968 37145 33977 37179
rect 33977 37145 34011 37179
rect 34011 37145 34020 37179
rect 33968 37136 34020 37145
rect 35256 37247 35308 37256
rect 35256 37213 35265 37247
rect 35265 37213 35299 37247
rect 35299 37213 35308 37247
rect 35256 37204 35308 37213
rect 37464 37204 37516 37256
rect 37648 37204 37700 37256
rect 37924 37204 37976 37256
rect 42156 37247 42208 37256
rect 42156 37213 42165 37247
rect 42165 37213 42199 37247
rect 42199 37213 42208 37247
rect 42156 37204 42208 37213
rect 35348 37136 35400 37188
rect 27896 37068 27948 37120
rect 31300 37068 31352 37120
rect 31576 37068 31628 37120
rect 32496 37111 32548 37120
rect 32496 37077 32505 37111
rect 32505 37077 32539 37111
rect 32539 37077 32548 37111
rect 32496 37068 32548 37077
rect 36360 37068 36412 37120
rect 37280 37068 37332 37120
rect 41052 37068 41104 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 3240 36660 3292 36712
rect 5448 36796 5500 36848
rect 7288 36839 7340 36848
rect 7288 36805 7297 36839
rect 7297 36805 7331 36839
rect 7331 36805 7340 36839
rect 7288 36796 7340 36805
rect 8116 36771 8168 36780
rect 8116 36737 8125 36771
rect 8125 36737 8159 36771
rect 8159 36737 8168 36771
rect 8116 36728 8168 36737
rect 15936 36771 15988 36780
rect 15936 36737 15945 36771
rect 15945 36737 15979 36771
rect 15979 36737 15988 36771
rect 15936 36728 15988 36737
rect 16764 36728 16816 36780
rect 20260 36864 20312 36916
rect 23204 36907 23256 36916
rect 23204 36873 23213 36907
rect 23213 36873 23247 36907
rect 23247 36873 23256 36907
rect 23204 36864 23256 36873
rect 23940 36864 23992 36916
rect 25044 36907 25096 36916
rect 25044 36873 25053 36907
rect 25053 36873 25087 36907
rect 25087 36873 25096 36907
rect 25044 36864 25096 36873
rect 25596 36864 25648 36916
rect 4068 36703 4120 36712
rect 4068 36669 4077 36703
rect 4077 36669 4111 36703
rect 4111 36669 4120 36703
rect 4068 36660 4120 36669
rect 15568 36703 15620 36712
rect 15568 36669 15577 36703
rect 15577 36669 15611 36703
rect 15611 36669 15620 36703
rect 15568 36660 15620 36669
rect 16856 36660 16908 36712
rect 17040 36660 17092 36712
rect 18788 36771 18840 36780
rect 18788 36737 18797 36771
rect 18797 36737 18831 36771
rect 18831 36737 18840 36771
rect 18788 36728 18840 36737
rect 19064 36728 19116 36780
rect 22836 36796 22888 36848
rect 18144 36592 18196 36644
rect 19340 36592 19392 36644
rect 19892 36728 19944 36780
rect 19616 36592 19668 36644
rect 21364 36728 21416 36780
rect 23480 36796 23532 36848
rect 23664 36796 23716 36848
rect 20812 36703 20864 36712
rect 20812 36669 20821 36703
rect 20821 36669 20855 36703
rect 20855 36669 20864 36703
rect 20812 36660 20864 36669
rect 21180 36660 21232 36712
rect 22652 36703 22704 36712
rect 22652 36669 22661 36703
rect 22661 36669 22695 36703
rect 22695 36669 22704 36703
rect 22652 36660 22704 36669
rect 23020 36660 23072 36712
rect 29000 36864 29052 36916
rect 31392 36864 31444 36916
rect 32036 36864 32088 36916
rect 29092 36796 29144 36848
rect 27344 36660 27396 36712
rect 28816 36703 28868 36712
rect 28816 36669 28825 36703
rect 28825 36669 28859 36703
rect 28859 36669 28868 36703
rect 28816 36660 28868 36669
rect 28908 36660 28960 36712
rect 21640 36592 21692 36644
rect 4804 36524 4856 36576
rect 15016 36567 15068 36576
rect 15016 36533 15025 36567
rect 15025 36533 15059 36567
rect 15059 36533 15068 36567
rect 15016 36524 15068 36533
rect 15292 36524 15344 36576
rect 16672 36567 16724 36576
rect 16672 36533 16681 36567
rect 16681 36533 16715 36567
rect 16715 36533 16724 36567
rect 16672 36524 16724 36533
rect 17224 36524 17276 36576
rect 18052 36524 18104 36576
rect 19892 36524 19944 36576
rect 20168 36567 20220 36576
rect 20168 36533 20177 36567
rect 20177 36533 20211 36567
rect 20211 36533 20220 36567
rect 20168 36524 20220 36533
rect 25320 36524 25372 36576
rect 25780 36592 25832 36644
rect 27620 36592 27672 36644
rect 30656 36771 30708 36780
rect 30656 36737 30665 36771
rect 30665 36737 30699 36771
rect 30699 36737 30708 36771
rect 30656 36728 30708 36737
rect 31484 36796 31536 36848
rect 33692 36864 33744 36916
rect 34980 36864 35032 36916
rect 37464 36864 37516 36916
rect 38660 36864 38712 36916
rect 41052 36907 41104 36916
rect 41052 36873 41061 36907
rect 41061 36873 41095 36907
rect 41095 36873 41104 36907
rect 41052 36864 41104 36873
rect 35256 36796 35308 36848
rect 31116 36771 31168 36780
rect 31116 36737 31125 36771
rect 31125 36737 31159 36771
rect 31159 36737 31168 36771
rect 31116 36728 31168 36737
rect 31576 36771 31628 36780
rect 31576 36737 31585 36771
rect 31585 36737 31619 36771
rect 31619 36737 31628 36771
rect 31576 36728 31628 36737
rect 32128 36771 32180 36780
rect 32128 36737 32137 36771
rect 32137 36737 32171 36771
rect 32171 36737 32180 36771
rect 32128 36728 32180 36737
rect 33508 36728 33560 36780
rect 31300 36660 31352 36712
rect 32404 36703 32456 36712
rect 32404 36669 32413 36703
rect 32413 36669 32447 36703
rect 32447 36669 32456 36703
rect 32404 36660 32456 36669
rect 32864 36660 32916 36712
rect 34796 36703 34848 36712
rect 34796 36669 34805 36703
rect 34805 36669 34839 36703
rect 34839 36669 34848 36703
rect 34796 36660 34848 36669
rect 31208 36592 31260 36644
rect 29920 36524 29972 36576
rect 30472 36524 30524 36576
rect 33784 36524 33836 36576
rect 33968 36567 34020 36576
rect 33968 36533 33977 36567
rect 33977 36533 34011 36567
rect 34011 36533 34020 36567
rect 33968 36524 34020 36533
rect 35348 36728 35400 36780
rect 36360 36771 36412 36780
rect 36360 36737 36369 36771
rect 36369 36737 36403 36771
rect 36403 36737 36412 36771
rect 36360 36728 36412 36737
rect 37372 36728 37424 36780
rect 37648 36771 37700 36780
rect 37648 36737 37657 36771
rect 37657 36737 37691 36771
rect 37691 36737 37700 36771
rect 37648 36728 37700 36737
rect 36452 36703 36504 36712
rect 36452 36669 36461 36703
rect 36461 36669 36495 36703
rect 36495 36669 36504 36703
rect 36452 36660 36504 36669
rect 37924 36771 37976 36780
rect 37924 36737 37933 36771
rect 37933 36737 37967 36771
rect 37967 36737 37976 36771
rect 37924 36728 37976 36737
rect 38108 36771 38160 36780
rect 38108 36737 38118 36771
rect 38118 36737 38152 36771
rect 38152 36737 38160 36771
rect 38108 36728 38160 36737
rect 39028 36728 39080 36780
rect 39580 36660 39632 36712
rect 35716 36635 35768 36644
rect 35716 36601 35725 36635
rect 35725 36601 35759 36635
rect 35759 36601 35768 36635
rect 35716 36592 35768 36601
rect 35992 36635 36044 36644
rect 35992 36601 36001 36635
rect 36001 36601 36035 36635
rect 36035 36601 36044 36635
rect 35992 36592 36044 36601
rect 37556 36635 37608 36644
rect 37556 36601 37565 36635
rect 37565 36601 37599 36635
rect 37599 36601 37608 36635
rect 39948 36660 40000 36712
rect 42156 36728 42208 36780
rect 41144 36703 41196 36712
rect 41144 36669 41153 36703
rect 41153 36669 41187 36703
rect 41187 36669 41196 36703
rect 41144 36660 41196 36669
rect 41236 36703 41288 36712
rect 41236 36669 41245 36703
rect 41245 36669 41279 36703
rect 41279 36669 41288 36703
rect 41236 36660 41288 36669
rect 37556 36592 37608 36601
rect 40316 36592 40368 36644
rect 41328 36592 41380 36644
rect 37188 36524 37240 36576
rect 37464 36524 37516 36576
rect 38568 36524 38620 36576
rect 40684 36567 40736 36576
rect 40684 36533 40693 36567
rect 40693 36533 40727 36567
rect 40727 36533 40736 36567
rect 40684 36524 40736 36533
rect 40776 36524 40828 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4068 36320 4120 36372
rect 13912 36320 13964 36372
rect 3976 36184 4028 36236
rect 3884 36116 3936 36168
rect 4252 36091 4304 36100
rect 4252 36057 4261 36091
rect 4261 36057 4295 36091
rect 4295 36057 4304 36091
rect 4252 36048 4304 36057
rect 4620 36252 4672 36304
rect 5448 36252 5500 36304
rect 7288 36252 7340 36304
rect 16488 36252 16540 36304
rect 16764 36363 16816 36372
rect 16764 36329 16773 36363
rect 16773 36329 16807 36363
rect 16807 36329 16816 36363
rect 16764 36320 16816 36329
rect 19892 36363 19944 36372
rect 19892 36329 19901 36363
rect 19901 36329 19935 36363
rect 19935 36329 19944 36363
rect 19892 36320 19944 36329
rect 20444 36320 20496 36372
rect 25504 36320 25556 36372
rect 4712 36116 4764 36168
rect 6736 36116 6788 36168
rect 11060 36184 11112 36236
rect 12900 36184 12952 36236
rect 7012 36116 7064 36168
rect 8668 36159 8720 36168
rect 8668 36125 8677 36159
rect 8677 36125 8711 36159
rect 8711 36125 8720 36159
rect 8668 36116 8720 36125
rect 5540 36048 5592 36100
rect 4804 35980 4856 36032
rect 5356 35980 5408 36032
rect 6828 35980 6880 36032
rect 6920 36023 6972 36032
rect 6920 35989 6929 36023
rect 6929 35989 6963 36023
rect 6963 35989 6972 36023
rect 6920 35980 6972 35989
rect 7104 35980 7156 36032
rect 8392 36091 8444 36100
rect 8392 36057 8401 36091
rect 8401 36057 8435 36091
rect 8435 36057 8444 36091
rect 8392 36048 8444 36057
rect 13452 36116 13504 36168
rect 14096 36159 14148 36168
rect 14096 36125 14105 36159
rect 14105 36125 14139 36159
rect 14139 36125 14148 36159
rect 14096 36116 14148 36125
rect 14464 36116 14516 36168
rect 18052 36184 18104 36236
rect 16948 36159 17000 36168
rect 16948 36125 16958 36159
rect 16958 36125 16992 36159
rect 16992 36125 17000 36159
rect 16948 36116 17000 36125
rect 17132 36116 17184 36168
rect 8944 36023 8996 36032
rect 8944 35989 8953 36023
rect 8953 35989 8987 36023
rect 8987 35989 8996 36023
rect 8944 35980 8996 35989
rect 10324 36048 10376 36100
rect 10416 36091 10468 36100
rect 10416 36057 10425 36091
rect 10425 36057 10459 36091
rect 10459 36057 10468 36091
rect 10416 36048 10468 36057
rect 13728 35980 13780 36032
rect 14188 35980 14240 36032
rect 15292 36091 15344 36100
rect 15292 36057 15301 36091
rect 15301 36057 15335 36091
rect 15335 36057 15344 36091
rect 15292 36048 15344 36057
rect 15752 36048 15804 36100
rect 15936 35980 15988 36032
rect 18512 35980 18564 36032
rect 21180 36227 21232 36236
rect 21180 36193 21189 36227
rect 21189 36193 21223 36227
rect 21223 36193 21232 36227
rect 21180 36184 21232 36193
rect 21640 36184 21692 36236
rect 22652 36184 22704 36236
rect 23020 36184 23072 36236
rect 23388 36227 23440 36236
rect 23388 36193 23397 36227
rect 23397 36193 23431 36227
rect 23431 36193 23440 36227
rect 23388 36184 23440 36193
rect 21456 36116 21508 36168
rect 20904 36023 20956 36032
rect 20904 35989 20913 36023
rect 20913 35989 20947 36023
rect 20947 35989 20956 36023
rect 20904 35980 20956 35989
rect 21364 35980 21416 36032
rect 23480 36048 23532 36100
rect 24400 36116 24452 36168
rect 27068 36116 27120 36168
rect 30472 36320 30524 36372
rect 30656 36320 30708 36372
rect 30104 36252 30156 36304
rect 31116 36320 31168 36372
rect 32404 36320 32456 36372
rect 29092 36116 29144 36168
rect 30104 36159 30156 36168
rect 30104 36125 30113 36159
rect 30113 36125 30147 36159
rect 30147 36125 30156 36159
rect 30104 36116 30156 36125
rect 31024 36116 31076 36168
rect 31208 36159 31260 36168
rect 31208 36125 31217 36159
rect 31217 36125 31251 36159
rect 31251 36125 31260 36159
rect 31208 36116 31260 36125
rect 32496 36184 32548 36236
rect 34152 36320 34204 36372
rect 34796 36320 34848 36372
rect 36452 36320 36504 36372
rect 37188 36363 37240 36372
rect 37188 36329 37197 36363
rect 37197 36329 37231 36363
rect 37231 36329 37240 36363
rect 37188 36320 37240 36329
rect 33968 36252 34020 36304
rect 34888 36252 34940 36304
rect 37924 36320 37976 36372
rect 39028 36363 39080 36372
rect 39028 36329 39037 36363
rect 39037 36329 39071 36363
rect 39071 36329 39080 36363
rect 39028 36320 39080 36329
rect 39948 36363 40000 36372
rect 39948 36329 39957 36363
rect 39957 36329 39991 36363
rect 39991 36329 40000 36363
rect 39948 36320 40000 36329
rect 40224 36320 40276 36372
rect 41236 36320 41288 36372
rect 42156 36363 42208 36372
rect 42156 36329 42165 36363
rect 42165 36329 42199 36363
rect 42199 36329 42208 36363
rect 42156 36320 42208 36329
rect 37464 36252 37516 36304
rect 37648 36252 37700 36304
rect 33784 36184 33836 36236
rect 36176 36184 36228 36236
rect 25320 36091 25372 36100
rect 25320 36057 25329 36091
rect 25329 36057 25363 36091
rect 25363 36057 25372 36091
rect 25320 36048 25372 36057
rect 23940 35980 23992 36032
rect 25136 35980 25188 36032
rect 25780 36048 25832 36100
rect 27804 36048 27856 36100
rect 28908 36048 28960 36100
rect 27344 35980 27396 36032
rect 29552 36023 29604 36032
rect 29552 35989 29561 36023
rect 29561 35989 29595 36023
rect 29595 35989 29604 36023
rect 29552 35980 29604 35989
rect 30472 36091 30524 36100
rect 30472 36057 30481 36091
rect 30481 36057 30515 36091
rect 30515 36057 30524 36091
rect 30472 36048 30524 36057
rect 31484 36091 31536 36100
rect 31484 36057 31493 36091
rect 31493 36057 31527 36091
rect 31527 36057 31536 36091
rect 31484 36048 31536 36057
rect 31668 36048 31720 36100
rect 33416 36048 33468 36100
rect 31208 35980 31260 36032
rect 35256 36116 35308 36168
rect 37280 36116 37332 36168
rect 37372 36159 37424 36168
rect 37372 36125 37381 36159
rect 37381 36125 37415 36159
rect 37415 36125 37424 36159
rect 37372 36116 37424 36125
rect 37556 36116 37608 36168
rect 38936 36252 38988 36304
rect 39580 36252 39632 36304
rect 40040 36252 40092 36304
rect 33784 36048 33836 36100
rect 34612 36048 34664 36100
rect 34796 36048 34848 36100
rect 34520 35980 34572 36032
rect 36084 35980 36136 36032
rect 38016 36116 38068 36168
rect 40684 36227 40736 36236
rect 40684 36193 40693 36227
rect 40693 36193 40727 36227
rect 40727 36193 40736 36227
rect 40684 36184 40736 36193
rect 38660 36159 38712 36168
rect 38660 36125 38669 36159
rect 38669 36125 38703 36159
rect 38703 36125 38712 36159
rect 38660 36116 38712 36125
rect 38936 36116 38988 36168
rect 39304 36159 39356 36168
rect 39304 36125 39313 36159
rect 39313 36125 39347 36159
rect 39347 36125 39356 36159
rect 39304 36116 39356 36125
rect 39580 36116 39632 36168
rect 38476 36048 38528 36100
rect 38568 36091 38620 36100
rect 38568 36057 38577 36091
rect 38577 36057 38611 36091
rect 38611 36057 38620 36091
rect 38568 36048 38620 36057
rect 39212 36048 39264 36100
rect 40040 36048 40092 36100
rect 40316 36091 40368 36100
rect 40316 36057 40325 36091
rect 40325 36057 40359 36091
rect 40359 36057 40368 36091
rect 40316 36048 40368 36057
rect 41420 36048 41472 36100
rect 38752 35980 38804 36032
rect 40224 35980 40276 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 3884 35776 3936 35828
rect 3240 35708 3292 35760
rect 4620 35708 4672 35760
rect 4804 35708 4856 35760
rect 4712 35683 4764 35692
rect 4712 35649 4721 35683
rect 4721 35649 4755 35683
rect 4755 35649 4764 35683
rect 4712 35640 4764 35649
rect 4988 35683 5040 35692
rect 4988 35649 4997 35683
rect 4997 35649 5031 35683
rect 5031 35649 5040 35683
rect 4988 35640 5040 35649
rect 5356 35683 5408 35692
rect 5356 35649 5365 35683
rect 5365 35649 5399 35683
rect 5399 35649 5408 35683
rect 5356 35640 5408 35649
rect 8392 35819 8444 35828
rect 8392 35785 8401 35819
rect 8401 35785 8435 35819
rect 8435 35785 8444 35819
rect 8392 35776 8444 35785
rect 10416 35776 10468 35828
rect 14096 35776 14148 35828
rect 14464 35776 14516 35828
rect 5540 35751 5592 35760
rect 5540 35717 5549 35751
rect 5549 35717 5583 35751
rect 5583 35717 5592 35751
rect 5540 35708 5592 35717
rect 6828 35708 6880 35760
rect 8760 35751 8812 35760
rect 8760 35717 8769 35751
rect 8769 35717 8803 35751
rect 8803 35717 8812 35751
rect 8760 35708 8812 35717
rect 2964 35615 3016 35624
rect 2964 35581 2973 35615
rect 2973 35581 3007 35615
rect 3007 35581 3016 35615
rect 2964 35572 3016 35581
rect 4620 35572 4672 35624
rect 7288 35683 7340 35692
rect 7288 35649 7297 35683
rect 7297 35649 7331 35683
rect 7331 35649 7340 35683
rect 7288 35640 7340 35649
rect 7380 35640 7432 35692
rect 6828 35572 6880 35624
rect 3332 35436 3384 35488
rect 5356 35504 5408 35556
rect 5448 35504 5500 35556
rect 7104 35504 7156 35556
rect 9036 35683 9088 35692
rect 9036 35649 9045 35683
rect 9045 35649 9079 35683
rect 9079 35649 9088 35683
rect 9036 35640 9088 35649
rect 9956 35640 10008 35692
rect 10416 35640 10468 35692
rect 10508 35683 10560 35692
rect 10508 35649 10517 35683
rect 10517 35649 10551 35683
rect 10551 35649 10560 35683
rect 10508 35640 10560 35649
rect 8944 35572 8996 35624
rect 10784 35683 10836 35692
rect 10784 35649 10793 35683
rect 10793 35649 10827 35683
rect 10827 35649 10836 35683
rect 10784 35640 10836 35649
rect 10876 35683 10928 35692
rect 10876 35649 10885 35683
rect 10885 35649 10919 35683
rect 10919 35649 10928 35683
rect 10876 35640 10928 35649
rect 11060 35708 11112 35760
rect 13452 35708 13504 35760
rect 13728 35708 13780 35760
rect 15016 35708 15068 35760
rect 15752 35708 15804 35760
rect 17040 35776 17092 35828
rect 22744 35776 22796 35828
rect 22928 35819 22980 35828
rect 22928 35785 22937 35819
rect 22937 35785 22971 35819
rect 22971 35785 22980 35819
rect 22928 35776 22980 35785
rect 17132 35708 17184 35760
rect 18604 35708 18656 35760
rect 21180 35708 21232 35760
rect 22560 35708 22612 35760
rect 26240 35776 26292 35828
rect 27804 35776 27856 35828
rect 28448 35819 28500 35828
rect 28448 35785 28457 35819
rect 28457 35785 28491 35819
rect 28491 35785 28500 35819
rect 28448 35776 28500 35785
rect 30472 35776 30524 35828
rect 31668 35819 31720 35828
rect 31668 35785 31677 35819
rect 31677 35785 31711 35819
rect 31711 35785 31720 35819
rect 31668 35776 31720 35785
rect 34888 35776 34940 35828
rect 35440 35776 35492 35828
rect 23480 35708 23532 35760
rect 13360 35640 13412 35692
rect 12256 35572 12308 35624
rect 12440 35572 12492 35624
rect 14096 35640 14148 35692
rect 14188 35683 14240 35692
rect 14188 35649 14197 35683
rect 14197 35649 14231 35683
rect 14231 35649 14240 35683
rect 14188 35640 14240 35649
rect 14464 35683 14516 35692
rect 14464 35649 14473 35683
rect 14473 35649 14507 35683
rect 14507 35649 14516 35683
rect 14464 35640 14516 35649
rect 17592 35640 17644 35692
rect 15108 35572 15160 35624
rect 13360 35504 13412 35556
rect 17040 35615 17092 35624
rect 17040 35581 17049 35615
rect 17049 35581 17083 35615
rect 17083 35581 17092 35615
rect 17040 35572 17092 35581
rect 4988 35436 5040 35488
rect 5540 35436 5592 35488
rect 8760 35436 8812 35488
rect 10232 35436 10284 35488
rect 10416 35436 10468 35488
rect 10600 35479 10652 35488
rect 10600 35445 10609 35479
rect 10609 35445 10643 35479
rect 10643 35445 10652 35479
rect 10600 35436 10652 35445
rect 12624 35436 12676 35488
rect 16856 35504 16908 35556
rect 19984 35640 20036 35692
rect 21548 35683 21600 35692
rect 21548 35649 21557 35683
rect 21557 35649 21591 35683
rect 21591 35649 21600 35683
rect 21548 35640 21600 35649
rect 25136 35708 25188 35760
rect 29552 35708 29604 35760
rect 31760 35751 31812 35760
rect 31760 35717 31769 35751
rect 31769 35717 31803 35751
rect 31803 35717 31812 35751
rect 31760 35708 31812 35717
rect 34520 35751 34572 35760
rect 34520 35717 34529 35751
rect 34529 35717 34563 35751
rect 34563 35717 34572 35751
rect 34520 35708 34572 35717
rect 34796 35708 34848 35760
rect 39304 35819 39356 35828
rect 39304 35785 39313 35819
rect 39313 35785 39347 35819
rect 39347 35785 39356 35819
rect 39304 35776 39356 35785
rect 18236 35572 18288 35624
rect 20904 35504 20956 35556
rect 17316 35436 17368 35488
rect 17684 35479 17736 35488
rect 17684 35445 17693 35479
rect 17693 35445 17727 35479
rect 17727 35445 17736 35479
rect 17684 35436 17736 35445
rect 20536 35479 20588 35488
rect 20536 35445 20545 35479
rect 20545 35445 20579 35479
rect 20579 35445 20588 35479
rect 20536 35436 20588 35445
rect 21640 35572 21692 35624
rect 22376 35615 22428 35624
rect 22376 35581 22385 35615
rect 22385 35581 22419 35615
rect 22419 35581 22428 35615
rect 22376 35572 22428 35581
rect 24676 35615 24728 35624
rect 24676 35581 24685 35615
rect 24685 35581 24719 35615
rect 24719 35581 24728 35615
rect 24676 35572 24728 35581
rect 25412 35572 25464 35624
rect 28908 35572 28960 35624
rect 22100 35436 22152 35488
rect 30196 35504 30248 35556
rect 31024 35572 31076 35624
rect 33324 35615 33376 35624
rect 33324 35581 33333 35615
rect 33333 35581 33367 35615
rect 33367 35581 33376 35615
rect 33324 35572 33376 35581
rect 35164 35683 35216 35692
rect 35164 35649 35173 35683
rect 35173 35649 35207 35683
rect 35207 35649 35216 35683
rect 35164 35640 35216 35649
rect 33232 35504 33284 35556
rect 34520 35572 34572 35624
rect 36084 35640 36136 35692
rect 25412 35436 25464 35488
rect 26332 35436 26384 35488
rect 29828 35479 29880 35488
rect 29828 35445 29837 35479
rect 29837 35445 29871 35479
rect 29871 35445 29880 35479
rect 29828 35436 29880 35445
rect 32404 35436 32456 35488
rect 34152 35504 34204 35556
rect 35808 35572 35860 35624
rect 38660 35708 38712 35760
rect 39212 35708 39264 35760
rect 38936 35640 38988 35692
rect 39764 35708 39816 35760
rect 41328 35819 41380 35828
rect 41328 35785 41337 35819
rect 41337 35785 41371 35819
rect 41371 35785 41380 35819
rect 41328 35776 41380 35785
rect 41420 35708 41472 35760
rect 38108 35615 38160 35624
rect 38108 35581 38117 35615
rect 38117 35581 38151 35615
rect 38151 35581 38160 35615
rect 38108 35572 38160 35581
rect 35440 35504 35492 35556
rect 38476 35572 38528 35624
rect 39580 35683 39632 35692
rect 39580 35649 39589 35683
rect 39589 35649 39623 35683
rect 39623 35649 39632 35683
rect 39580 35640 39632 35649
rect 38752 35504 38804 35556
rect 34428 35436 34480 35488
rect 34796 35436 34848 35488
rect 35348 35479 35400 35488
rect 35348 35445 35357 35479
rect 35357 35445 35391 35479
rect 35391 35445 35400 35479
rect 35348 35436 35400 35445
rect 37648 35479 37700 35488
rect 37648 35445 37657 35479
rect 37657 35445 37691 35479
rect 37691 35445 37700 35479
rect 37648 35436 37700 35445
rect 39856 35615 39908 35624
rect 39856 35581 39865 35615
rect 39865 35581 39899 35615
rect 39899 35581 39908 35615
rect 39856 35572 39908 35581
rect 41236 35572 41288 35624
rect 40040 35436 40092 35488
rect 42156 35479 42208 35488
rect 42156 35445 42165 35479
rect 42165 35445 42199 35479
rect 42199 35445 42208 35479
rect 42156 35436 42208 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 2964 35232 3016 35284
rect 4068 35232 4120 35284
rect 4896 35232 4948 35284
rect 5356 35232 5408 35284
rect 7380 35232 7432 35284
rect 7012 35164 7064 35216
rect 10508 35232 10560 35284
rect 12256 35275 12308 35284
rect 12256 35241 12265 35275
rect 12265 35241 12299 35275
rect 12299 35241 12308 35275
rect 12256 35232 12308 35241
rect 13176 35232 13228 35284
rect 13636 35232 13688 35284
rect 15568 35232 15620 35284
rect 17316 35232 17368 35284
rect 18144 35232 18196 35284
rect 18236 35232 18288 35284
rect 24676 35232 24728 35284
rect 29276 35232 29328 35284
rect 31024 35232 31076 35284
rect 34520 35232 34572 35284
rect 35348 35232 35400 35284
rect 38660 35232 38712 35284
rect 39764 35232 39816 35284
rect 39856 35232 39908 35284
rect 41420 35232 41472 35284
rect 3332 35071 3384 35080
rect 3332 35037 3341 35071
rect 3341 35037 3375 35071
rect 3375 35037 3384 35071
rect 3332 35028 3384 35037
rect 3516 35071 3568 35080
rect 3516 35037 3525 35071
rect 3525 35037 3559 35071
rect 3559 35037 3568 35071
rect 3516 35028 3568 35037
rect 3884 35028 3936 35080
rect 4068 35028 4120 35080
rect 5540 35139 5592 35148
rect 5540 35105 5549 35139
rect 5549 35105 5583 35139
rect 5583 35105 5592 35139
rect 5540 35096 5592 35105
rect 5264 35071 5316 35080
rect 5264 35037 5273 35071
rect 5273 35037 5307 35071
rect 5307 35037 5316 35071
rect 5264 35028 5316 35037
rect 6920 35028 6972 35080
rect 8944 35164 8996 35216
rect 9036 35164 9088 35216
rect 10784 35164 10836 35216
rect 4712 35003 4764 35012
rect 4712 34969 4739 35003
rect 4739 34969 4764 35003
rect 4712 34960 4764 34969
rect 4804 34960 4856 35012
rect 4988 34960 5040 35012
rect 7104 34960 7156 35012
rect 7748 34960 7800 35012
rect 10600 35028 10652 35080
rect 12440 35071 12492 35080
rect 12440 35037 12449 35071
rect 12449 35037 12483 35071
rect 12483 35037 12492 35071
rect 12440 35028 12492 35037
rect 14188 35164 14240 35216
rect 13820 35096 13872 35148
rect 16672 35164 16724 35216
rect 15936 35096 15988 35148
rect 17132 35139 17184 35148
rect 17132 35105 17141 35139
rect 17141 35105 17175 35139
rect 17175 35105 17184 35139
rect 17132 35096 17184 35105
rect 9036 34960 9088 35012
rect 4436 34892 4488 34944
rect 4528 34935 4580 34944
rect 4528 34901 4537 34935
rect 4537 34901 4571 34935
rect 4571 34901 4580 34935
rect 4528 34892 4580 34901
rect 6828 34892 6880 34944
rect 9312 34892 9364 34944
rect 10876 34892 10928 34944
rect 14648 35028 14700 35080
rect 16028 35071 16080 35080
rect 16028 35037 16037 35071
rect 16037 35037 16071 35071
rect 16071 35037 16080 35071
rect 16028 35028 16080 35037
rect 17684 35028 17736 35080
rect 18604 35028 18656 35080
rect 22100 35096 22152 35148
rect 23020 35096 23072 35148
rect 23388 35139 23440 35148
rect 23388 35105 23397 35139
rect 23397 35105 23431 35139
rect 23431 35105 23440 35139
rect 23388 35096 23440 35105
rect 24768 35096 24820 35148
rect 26332 35096 26384 35148
rect 35808 35164 35860 35216
rect 29828 35139 29880 35148
rect 29828 35105 29837 35139
rect 29837 35105 29871 35139
rect 29871 35105 29880 35139
rect 29828 35096 29880 35105
rect 31484 35096 31536 35148
rect 32128 35139 32180 35148
rect 32128 35105 32137 35139
rect 32137 35105 32171 35139
rect 32171 35105 32180 35139
rect 32128 35096 32180 35105
rect 32404 35139 32456 35148
rect 32404 35105 32413 35139
rect 32413 35105 32447 35139
rect 32447 35105 32456 35139
rect 32404 35096 32456 35105
rect 33416 35096 33468 35148
rect 35992 35139 36044 35148
rect 35992 35105 36001 35139
rect 36001 35105 36035 35139
rect 36035 35105 36044 35139
rect 35992 35096 36044 35105
rect 37096 35164 37148 35216
rect 13176 35003 13228 35012
rect 13176 34969 13185 35003
rect 13185 34969 13219 35003
rect 13219 34969 13228 35003
rect 13176 34960 13228 34969
rect 13360 35003 13412 35012
rect 13360 34969 13369 35003
rect 13369 34969 13403 35003
rect 13403 34969 13412 35003
rect 13360 34960 13412 34969
rect 13912 34960 13964 35012
rect 17224 34960 17276 35012
rect 17776 34960 17828 35012
rect 26240 35071 26292 35080
rect 26240 35037 26249 35071
rect 26249 35037 26283 35071
rect 26283 35037 26292 35071
rect 26240 35028 26292 35037
rect 14096 34892 14148 34944
rect 14464 34892 14516 34944
rect 15844 34892 15896 34944
rect 16672 34935 16724 34944
rect 16672 34901 16681 34935
rect 16681 34901 16715 34935
rect 16715 34901 16724 34935
rect 16672 34892 16724 34901
rect 19156 34892 19208 34944
rect 21364 34935 21416 34944
rect 21364 34901 21373 34935
rect 21373 34901 21407 34935
rect 21407 34901 21416 34935
rect 21364 34892 21416 34901
rect 22192 34960 22244 35012
rect 27068 34960 27120 35012
rect 27160 35003 27212 35012
rect 27160 34969 27169 35003
rect 27169 34969 27203 35003
rect 27203 34969 27212 35003
rect 27160 34960 27212 34969
rect 28816 34960 28868 35012
rect 33508 35028 33560 35080
rect 33784 35028 33836 35080
rect 29736 34960 29788 35012
rect 21916 34935 21968 34944
rect 21916 34901 21925 34935
rect 21925 34901 21959 34935
rect 21959 34901 21968 34935
rect 21916 34892 21968 34901
rect 22836 34935 22888 34944
rect 22836 34901 22845 34935
rect 22845 34901 22879 34935
rect 22879 34901 22888 34935
rect 22836 34892 22888 34901
rect 23204 34935 23256 34944
rect 23204 34901 23213 34935
rect 23213 34901 23247 34935
rect 23247 34901 23256 34935
rect 23204 34892 23256 34901
rect 25320 34935 25372 34944
rect 25320 34901 25329 34935
rect 25329 34901 25363 34935
rect 25363 34901 25372 34935
rect 25320 34892 25372 34901
rect 28724 34935 28776 34944
rect 28724 34901 28733 34935
rect 28733 34901 28767 34935
rect 28767 34901 28776 34935
rect 28724 34892 28776 34901
rect 30288 34960 30340 35012
rect 34428 34960 34480 35012
rect 37004 35071 37056 35080
rect 37004 35037 37013 35071
rect 37013 35037 37047 35071
rect 37047 35037 37056 35071
rect 37004 35028 37056 35037
rect 39580 35028 39632 35080
rect 40132 34960 40184 35012
rect 40316 35096 40368 35148
rect 40776 35028 40828 35080
rect 41328 35028 41380 35080
rect 41788 35071 41840 35080
rect 41788 35037 41797 35071
rect 41797 35037 41831 35071
rect 41831 35037 41840 35071
rect 41788 35028 41840 35037
rect 31392 34935 31444 34944
rect 31392 34901 31401 34935
rect 31401 34901 31435 34935
rect 31435 34901 31444 34935
rect 31392 34892 31444 34901
rect 34336 34892 34388 34944
rect 35348 34892 35400 34944
rect 36268 34892 36320 34944
rect 37556 34892 37608 34944
rect 39028 34935 39080 34944
rect 39028 34901 39037 34935
rect 39037 34901 39071 34935
rect 39071 34901 39080 34935
rect 39028 34892 39080 34901
rect 40592 34935 40644 34944
rect 40592 34901 40601 34935
rect 40601 34901 40635 34935
rect 40635 34901 40644 34935
rect 40592 34892 40644 34901
rect 40960 34935 41012 34944
rect 40960 34901 40969 34935
rect 40969 34901 41003 34935
rect 41003 34901 41012 34935
rect 40960 34892 41012 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 3516 34688 3568 34740
rect 4528 34620 4580 34672
rect 3240 34484 3292 34536
rect 3976 34484 4028 34536
rect 5356 34595 5408 34604
rect 5356 34561 5365 34595
rect 5365 34561 5399 34595
rect 5399 34561 5408 34595
rect 5356 34552 5408 34561
rect 6828 34552 6880 34604
rect 8300 34552 8352 34604
rect 11428 34688 11480 34740
rect 16028 34688 16080 34740
rect 17224 34731 17276 34740
rect 17224 34697 17233 34731
rect 17233 34697 17267 34731
rect 17267 34697 17276 34731
rect 17224 34688 17276 34697
rect 8944 34620 8996 34672
rect 10600 34620 10652 34672
rect 13452 34620 13504 34672
rect 15752 34620 15804 34672
rect 19156 34731 19208 34740
rect 19156 34697 19165 34731
rect 19165 34697 19199 34731
rect 19199 34697 19208 34731
rect 19156 34688 19208 34697
rect 19248 34688 19300 34740
rect 9128 34595 9180 34604
rect 9128 34561 9137 34595
rect 9137 34561 9171 34595
rect 9171 34561 9180 34595
rect 9128 34552 9180 34561
rect 9312 34595 9364 34604
rect 9312 34561 9321 34595
rect 9321 34561 9355 34595
rect 9355 34561 9364 34595
rect 9312 34552 9364 34561
rect 16396 34552 16448 34604
rect 9036 34484 9088 34536
rect 9588 34527 9640 34536
rect 9588 34493 9597 34527
rect 9597 34493 9631 34527
rect 9631 34493 9640 34527
rect 9588 34484 9640 34493
rect 11428 34484 11480 34536
rect 12900 34527 12952 34536
rect 12900 34493 12909 34527
rect 12909 34493 12943 34527
rect 12943 34493 12952 34527
rect 12900 34484 12952 34493
rect 14556 34484 14608 34536
rect 17132 34484 17184 34536
rect 18604 34595 18656 34604
rect 18604 34561 18613 34595
rect 18613 34561 18647 34595
rect 18647 34561 18656 34595
rect 18604 34552 18656 34561
rect 19340 34552 19392 34604
rect 20536 34620 20588 34672
rect 20904 34688 20956 34740
rect 22560 34688 22612 34740
rect 23480 34688 23532 34740
rect 24860 34731 24912 34740
rect 24860 34697 24869 34731
rect 24869 34697 24903 34731
rect 24903 34697 24912 34731
rect 24860 34688 24912 34697
rect 25320 34688 25372 34740
rect 27160 34688 27212 34740
rect 28724 34688 28776 34740
rect 22836 34620 22888 34672
rect 25596 34620 25648 34672
rect 29092 34663 29144 34672
rect 29092 34629 29101 34663
rect 29101 34629 29135 34663
rect 29135 34629 29144 34663
rect 29092 34620 29144 34629
rect 30288 34620 30340 34672
rect 31484 34731 31536 34740
rect 31484 34697 31493 34731
rect 31493 34697 31527 34731
rect 31527 34697 31536 34731
rect 31484 34688 31536 34697
rect 38292 34688 38344 34740
rect 5356 34416 5408 34468
rect 8576 34459 8628 34468
rect 8576 34425 8585 34459
rect 8585 34425 8619 34459
rect 8619 34425 8628 34459
rect 8576 34416 8628 34425
rect 19248 34527 19300 34536
rect 19248 34493 19257 34527
rect 19257 34493 19291 34527
rect 19291 34493 19300 34527
rect 19248 34484 19300 34493
rect 24124 34595 24176 34604
rect 24124 34561 24133 34595
rect 24133 34561 24167 34595
rect 24167 34561 24176 34595
rect 24124 34552 24176 34561
rect 22008 34484 22060 34536
rect 23664 34527 23716 34536
rect 23664 34493 23673 34527
rect 23673 34493 23707 34527
rect 23707 34493 23716 34527
rect 23664 34484 23716 34493
rect 23848 34484 23900 34536
rect 25136 34484 25188 34536
rect 25412 34484 25464 34536
rect 27988 34527 28040 34536
rect 27988 34493 27997 34527
rect 27997 34493 28031 34527
rect 28031 34493 28040 34527
rect 27988 34484 28040 34493
rect 28172 34527 28224 34536
rect 28172 34493 28181 34527
rect 28181 34493 28215 34527
rect 28215 34493 28224 34527
rect 28172 34484 28224 34493
rect 28908 34484 28960 34536
rect 29736 34527 29788 34536
rect 29736 34493 29745 34527
rect 29745 34493 29779 34527
rect 29779 34493 29788 34527
rect 29736 34484 29788 34493
rect 30012 34527 30064 34536
rect 30012 34493 30021 34527
rect 30021 34493 30055 34527
rect 30055 34493 30064 34527
rect 30012 34484 30064 34493
rect 30748 34484 30800 34536
rect 31300 34552 31352 34604
rect 32128 34595 32180 34604
rect 32128 34561 32137 34595
rect 32137 34561 32171 34595
rect 32171 34561 32180 34595
rect 32128 34552 32180 34561
rect 4804 34348 4856 34400
rect 5632 34391 5684 34400
rect 5632 34357 5641 34391
rect 5641 34357 5675 34391
rect 5675 34357 5684 34391
rect 5632 34348 5684 34357
rect 6920 34348 6972 34400
rect 9680 34348 9732 34400
rect 10048 34348 10100 34400
rect 13912 34348 13964 34400
rect 23020 34348 23072 34400
rect 31116 34416 31168 34468
rect 32772 34484 32824 34536
rect 34336 34663 34388 34672
rect 34336 34629 34345 34663
rect 34345 34629 34379 34663
rect 34379 34629 34388 34663
rect 34336 34620 34388 34629
rect 34428 34620 34480 34672
rect 34796 34620 34848 34672
rect 35532 34620 35584 34672
rect 37096 34620 37148 34672
rect 37648 34620 37700 34672
rect 40132 34731 40184 34740
rect 40132 34697 40141 34731
rect 40141 34697 40175 34731
rect 40175 34697 40184 34731
rect 40132 34688 40184 34697
rect 41144 34688 41196 34740
rect 41236 34731 41288 34740
rect 41236 34697 41245 34731
rect 41245 34697 41279 34731
rect 41279 34697 41288 34731
rect 41236 34688 41288 34697
rect 41328 34731 41380 34740
rect 41328 34697 41337 34731
rect 41337 34697 41371 34731
rect 41371 34697 41380 34731
rect 41328 34688 41380 34697
rect 39580 34620 39632 34672
rect 41696 34663 41748 34672
rect 41696 34629 41705 34663
rect 41705 34629 41739 34663
rect 41739 34629 41748 34663
rect 41696 34620 41748 34629
rect 34428 34527 34480 34536
rect 34428 34493 34437 34527
rect 34437 34493 34471 34527
rect 34471 34493 34480 34527
rect 34428 34484 34480 34493
rect 38660 34552 38712 34604
rect 39120 34595 39172 34604
rect 39120 34561 39129 34595
rect 39129 34561 39163 34595
rect 39163 34561 39172 34595
rect 39120 34552 39172 34561
rect 39212 34552 39264 34604
rect 34796 34527 34848 34536
rect 34796 34493 34805 34527
rect 34805 34493 34839 34527
rect 34839 34493 34848 34527
rect 34796 34484 34848 34493
rect 33508 34416 33560 34468
rect 35532 34484 35584 34536
rect 35624 34484 35676 34536
rect 37280 34527 37332 34536
rect 37280 34493 37289 34527
rect 37289 34493 37323 34527
rect 37323 34493 37332 34527
rect 37280 34484 37332 34493
rect 38936 34484 38988 34536
rect 41880 34595 41932 34604
rect 41880 34561 41889 34595
rect 41889 34561 41923 34595
rect 41923 34561 41932 34595
rect 41880 34552 41932 34561
rect 37004 34416 37056 34468
rect 23756 34391 23808 34400
rect 23756 34357 23765 34391
rect 23765 34357 23799 34391
rect 23799 34357 23808 34391
rect 23756 34348 23808 34357
rect 25320 34348 25372 34400
rect 33968 34391 34020 34400
rect 33968 34357 33977 34391
rect 33977 34357 34011 34391
rect 34011 34357 34020 34391
rect 33968 34348 34020 34357
rect 35532 34348 35584 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5632 34144 5684 34196
rect 8576 34144 8628 34196
rect 9680 34187 9732 34196
rect 9680 34153 9689 34187
rect 9689 34153 9723 34187
rect 9723 34153 9732 34187
rect 9680 34144 9732 34153
rect 9772 34144 9824 34196
rect 10600 34144 10652 34196
rect 11152 34144 11204 34196
rect 11428 34144 11480 34196
rect 13820 34144 13872 34196
rect 13912 34144 13964 34196
rect 16396 34187 16448 34196
rect 16396 34153 16405 34187
rect 16405 34153 16439 34187
rect 16439 34153 16448 34187
rect 16396 34144 16448 34153
rect 19248 34144 19300 34196
rect 20996 34187 21048 34196
rect 20996 34153 21005 34187
rect 21005 34153 21039 34187
rect 21039 34153 21048 34187
rect 20996 34144 21048 34153
rect 25872 34187 25924 34196
rect 25872 34153 25881 34187
rect 25881 34153 25915 34187
rect 25915 34153 25924 34187
rect 25872 34144 25924 34153
rect 27712 34144 27764 34196
rect 30196 34187 30248 34196
rect 30196 34153 30205 34187
rect 30205 34153 30239 34187
rect 30239 34153 30248 34187
rect 30196 34144 30248 34153
rect 33048 34144 33100 34196
rect 9128 34076 9180 34128
rect 5264 34008 5316 34060
rect 8300 34008 8352 34060
rect 8576 34008 8628 34060
rect 10048 34008 10100 34060
rect 5908 33983 5960 33992
rect 5908 33949 5917 33983
rect 5917 33949 5951 33983
rect 5951 33949 5960 33983
rect 5908 33940 5960 33949
rect 9772 33940 9824 33992
rect 9864 33983 9916 33992
rect 9864 33949 9873 33983
rect 9873 33949 9907 33983
rect 9907 33949 9916 33983
rect 9864 33940 9916 33949
rect 17500 34076 17552 34128
rect 10968 34008 11020 34060
rect 6920 33872 6972 33924
rect 7012 33915 7064 33924
rect 7012 33881 7021 33915
rect 7021 33881 7055 33915
rect 7055 33881 7064 33915
rect 7012 33872 7064 33881
rect 8668 33872 8720 33924
rect 11060 33940 11112 33992
rect 12900 34008 12952 34060
rect 13452 34008 13504 34060
rect 14648 34051 14700 34060
rect 14648 34017 14657 34051
rect 14657 34017 14691 34051
rect 14691 34017 14700 34051
rect 14648 34008 14700 34017
rect 16488 34008 16540 34060
rect 16672 34008 16724 34060
rect 17040 34051 17092 34060
rect 17040 34017 17049 34051
rect 17049 34017 17083 34051
rect 17083 34017 17092 34051
rect 17040 34008 17092 34017
rect 18604 34008 18656 34060
rect 33784 34187 33836 34196
rect 33784 34153 33793 34187
rect 33793 34153 33827 34187
rect 33827 34153 33836 34187
rect 33784 34144 33836 34153
rect 39212 34144 39264 34196
rect 40592 34144 40644 34196
rect 41972 34076 42024 34128
rect 26424 34051 26476 34060
rect 26424 34017 26433 34051
rect 26433 34017 26467 34051
rect 26467 34017 26476 34051
rect 26424 34008 26476 34017
rect 30840 34051 30892 34060
rect 30840 34017 30849 34051
rect 30849 34017 30883 34051
rect 30883 34017 30892 34051
rect 30840 34008 30892 34017
rect 31668 34008 31720 34060
rect 32036 34051 32088 34060
rect 32036 34017 32045 34051
rect 32045 34017 32079 34051
rect 32079 34017 32088 34051
rect 32036 34008 32088 34017
rect 33968 34008 34020 34060
rect 34796 34008 34848 34060
rect 35624 34008 35676 34060
rect 37280 34051 37332 34060
rect 37280 34017 37289 34051
rect 37289 34017 37323 34051
rect 37323 34017 37332 34051
rect 37280 34008 37332 34017
rect 39580 34008 39632 34060
rect 40684 34051 40736 34060
rect 40684 34017 40693 34051
rect 40693 34017 40727 34051
rect 40727 34017 40736 34051
rect 40684 34008 40736 34017
rect 41696 34008 41748 34060
rect 14464 33983 14516 33992
rect 14464 33949 14473 33983
rect 14473 33949 14507 33983
rect 14507 33949 14516 33983
rect 14464 33940 14516 33949
rect 14556 33940 14608 33992
rect 15660 33983 15712 33992
rect 15660 33949 15669 33983
rect 15669 33949 15703 33983
rect 15703 33949 15712 33983
rect 15660 33940 15712 33949
rect 15844 33983 15896 33992
rect 15844 33949 15853 33983
rect 15853 33949 15887 33983
rect 15887 33949 15896 33983
rect 15844 33940 15896 33949
rect 22100 33983 22152 33992
rect 22100 33949 22109 33983
rect 22109 33949 22143 33983
rect 22143 33949 22152 33983
rect 22100 33940 22152 33949
rect 23664 33940 23716 33992
rect 24400 33983 24452 33992
rect 24400 33949 24409 33983
rect 24409 33949 24443 33983
rect 24443 33949 24452 33983
rect 24400 33940 24452 33949
rect 31116 33940 31168 33992
rect 33416 33940 33468 33992
rect 38660 33940 38712 33992
rect 40960 33940 41012 33992
rect 41328 33983 41380 33992
rect 41328 33949 41337 33983
rect 41337 33949 41371 33983
rect 41371 33949 41380 33983
rect 41328 33940 41380 33949
rect 12532 33872 12584 33924
rect 19800 33872 19852 33924
rect 21456 33872 21508 33924
rect 5724 33847 5776 33856
rect 5724 33813 5733 33847
rect 5733 33813 5767 33847
rect 5767 33813 5776 33847
rect 5724 33804 5776 33813
rect 8944 33847 8996 33856
rect 8944 33813 8953 33847
rect 8953 33813 8987 33847
rect 8987 33813 8996 33847
rect 8944 33804 8996 33813
rect 10140 33804 10192 33856
rect 11336 33804 11388 33856
rect 17316 33804 17368 33856
rect 21088 33847 21140 33856
rect 21088 33813 21097 33847
rect 21097 33813 21131 33847
rect 21131 33813 21140 33847
rect 21088 33804 21140 33813
rect 23940 33872 23992 33924
rect 24768 33872 24820 33924
rect 26700 33915 26752 33924
rect 26700 33881 26709 33915
rect 26709 33881 26743 33915
rect 26743 33881 26752 33915
rect 26700 33872 26752 33881
rect 27068 33872 27120 33924
rect 28724 33872 28776 33924
rect 31576 33872 31628 33924
rect 35348 33872 35400 33924
rect 35532 33872 35584 33924
rect 37556 33915 37608 33924
rect 37556 33881 37565 33915
rect 37565 33881 37599 33915
rect 37599 33881 37608 33915
rect 37556 33872 37608 33881
rect 22376 33804 22428 33856
rect 23204 33804 23256 33856
rect 25136 33804 25188 33856
rect 26240 33847 26292 33856
rect 26240 33813 26249 33847
rect 26249 33813 26283 33847
rect 26283 33813 26292 33847
rect 26240 33804 26292 33813
rect 26332 33847 26384 33856
rect 26332 33813 26341 33847
rect 26341 33813 26375 33847
rect 26375 33813 26384 33847
rect 26332 33804 26384 33813
rect 28356 33847 28408 33856
rect 28356 33813 28365 33847
rect 28365 33813 28399 33847
rect 28399 33813 28408 33847
rect 28356 33804 28408 33813
rect 31484 33804 31536 33856
rect 36728 33847 36780 33856
rect 36728 33813 36737 33847
rect 36737 33813 36771 33847
rect 36771 33813 36780 33847
rect 36728 33804 36780 33813
rect 36820 33804 36872 33856
rect 41880 33872 41932 33924
rect 40224 33804 40276 33856
rect 40500 33847 40552 33856
rect 40500 33813 40509 33847
rect 40509 33813 40543 33847
rect 40543 33813 40552 33847
rect 40500 33804 40552 33813
rect 41236 33804 41288 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 3240 33600 3292 33652
rect 10968 33600 11020 33652
rect 12440 33600 12492 33652
rect 16580 33600 16632 33652
rect 18604 33600 18656 33652
rect 19800 33643 19852 33652
rect 19800 33609 19809 33643
rect 19809 33609 19843 33643
rect 19843 33609 19852 33643
rect 19800 33600 19852 33609
rect 21088 33600 21140 33652
rect 21916 33600 21968 33652
rect 23848 33643 23900 33652
rect 23848 33609 23857 33643
rect 23857 33609 23891 33643
rect 23891 33609 23900 33643
rect 23848 33600 23900 33609
rect 23940 33643 23992 33652
rect 23940 33609 23949 33643
rect 23949 33609 23983 33643
rect 23983 33609 23992 33643
rect 23940 33600 23992 33609
rect 24768 33643 24820 33652
rect 24768 33609 24777 33643
rect 24777 33609 24811 33643
rect 24811 33609 24820 33643
rect 24768 33600 24820 33609
rect 26792 33600 26844 33652
rect 27988 33600 28040 33652
rect 30012 33600 30064 33652
rect 31484 33643 31536 33652
rect 31484 33609 31493 33643
rect 31493 33609 31527 33643
rect 31527 33609 31536 33643
rect 31484 33600 31536 33609
rect 31576 33643 31628 33652
rect 31576 33609 31585 33643
rect 31585 33609 31619 33643
rect 31619 33609 31628 33643
rect 31576 33600 31628 33609
rect 33324 33600 33376 33652
rect 34244 33600 34296 33652
rect 34428 33600 34480 33652
rect 36268 33600 36320 33652
rect 38108 33600 38160 33652
rect 39028 33600 39080 33652
rect 41328 33643 41380 33652
rect 41328 33609 41337 33643
rect 41337 33609 41371 33643
rect 41371 33609 41380 33643
rect 41328 33600 41380 33609
rect 42156 33600 42208 33652
rect 3148 33532 3200 33584
rect 3608 33532 3660 33584
rect 1860 33464 1912 33516
rect 2136 33507 2188 33516
rect 2136 33473 2145 33507
rect 2145 33473 2179 33507
rect 2179 33473 2188 33507
rect 5264 33532 5316 33584
rect 5908 33532 5960 33584
rect 7656 33575 7708 33584
rect 7656 33541 7665 33575
rect 7665 33541 7699 33575
rect 7699 33541 7708 33575
rect 7656 33532 7708 33541
rect 8116 33532 8168 33584
rect 8300 33532 8352 33584
rect 2136 33464 2188 33473
rect 5356 33507 5408 33516
rect 5356 33473 5365 33507
rect 5365 33473 5399 33507
rect 5399 33473 5408 33507
rect 5356 33464 5408 33473
rect 5448 33507 5500 33516
rect 5448 33473 5457 33507
rect 5457 33473 5491 33507
rect 5491 33473 5500 33507
rect 5448 33464 5500 33473
rect 5540 33464 5592 33516
rect 8576 33464 8628 33516
rect 9588 33532 9640 33584
rect 13176 33532 13228 33584
rect 10600 33464 10652 33516
rect 11152 33464 11204 33516
rect 11336 33507 11388 33516
rect 11336 33473 11345 33507
rect 11345 33473 11379 33507
rect 11379 33473 11388 33507
rect 11336 33464 11388 33473
rect 12440 33464 12492 33516
rect 17224 33464 17276 33516
rect 26240 33532 26292 33584
rect 27252 33532 27304 33584
rect 31392 33532 31444 33584
rect 18236 33464 18288 33516
rect 4620 33439 4672 33448
rect 4620 33405 4629 33439
rect 4629 33405 4663 33439
rect 4663 33405 4672 33439
rect 4620 33396 4672 33405
rect 5172 33439 5224 33448
rect 5172 33405 5181 33439
rect 5181 33405 5215 33439
rect 5215 33405 5224 33439
rect 5172 33396 5224 33405
rect 5264 33439 5316 33448
rect 5264 33405 5273 33439
rect 5273 33405 5307 33439
rect 5307 33405 5316 33439
rect 5264 33396 5316 33405
rect 8668 33439 8720 33448
rect 8668 33405 8677 33439
rect 8677 33405 8711 33439
rect 8711 33405 8720 33439
rect 8668 33396 8720 33405
rect 9128 33396 9180 33448
rect 9496 33439 9548 33448
rect 9496 33405 9505 33439
rect 9505 33405 9539 33439
rect 9539 33405 9548 33439
rect 9496 33396 9548 33405
rect 11060 33371 11112 33380
rect 11060 33337 11069 33371
rect 11069 33337 11103 33371
rect 11103 33337 11112 33371
rect 11060 33328 11112 33337
rect 11428 33396 11480 33448
rect 12348 33439 12400 33448
rect 12348 33405 12357 33439
rect 12357 33405 12391 33439
rect 12391 33405 12400 33439
rect 12348 33396 12400 33405
rect 13084 33439 13136 33448
rect 13084 33405 13093 33439
rect 13093 33405 13127 33439
rect 13127 33405 13136 33439
rect 13084 33396 13136 33405
rect 12716 33328 12768 33380
rect 16764 33328 16816 33380
rect 18788 33507 18840 33516
rect 18788 33473 18833 33507
rect 18833 33473 18840 33507
rect 18788 33464 18840 33473
rect 18972 33507 19024 33516
rect 18972 33473 18981 33507
rect 18981 33473 19015 33507
rect 19015 33473 19024 33507
rect 18972 33464 19024 33473
rect 19800 33464 19852 33516
rect 21364 33464 21416 33516
rect 23204 33507 23256 33516
rect 23204 33473 23213 33507
rect 23213 33473 23247 33507
rect 23247 33473 23256 33507
rect 23204 33464 23256 33473
rect 23756 33464 23808 33516
rect 25412 33464 25464 33516
rect 26332 33464 26384 33516
rect 28264 33507 28316 33516
rect 28264 33473 28273 33507
rect 28273 33473 28307 33507
rect 28307 33473 28316 33507
rect 28264 33464 28316 33473
rect 28724 33464 28776 33516
rect 36820 33532 36872 33584
rect 20720 33396 20772 33448
rect 25228 33439 25280 33448
rect 25228 33405 25237 33439
rect 25237 33405 25271 33439
rect 25271 33405 25280 33439
rect 25228 33396 25280 33405
rect 25320 33439 25372 33448
rect 25320 33405 25329 33439
rect 25329 33405 25363 33439
rect 25363 33405 25372 33439
rect 25320 33396 25372 33405
rect 25964 33396 26016 33448
rect 26424 33396 26476 33448
rect 33048 33507 33100 33516
rect 33048 33473 33057 33507
rect 33057 33473 33091 33507
rect 33091 33473 33100 33507
rect 33048 33464 33100 33473
rect 34152 33464 34204 33516
rect 38292 33507 38344 33516
rect 38292 33473 38301 33507
rect 38301 33473 38335 33507
rect 38335 33473 38344 33507
rect 38292 33464 38344 33473
rect 38660 33464 38712 33516
rect 39580 33464 39632 33516
rect 40224 33507 40276 33516
rect 40224 33473 40258 33507
rect 40258 33473 40276 33507
rect 40224 33464 40276 33473
rect 41604 33464 41656 33516
rect 28908 33396 28960 33448
rect 20628 33328 20680 33380
rect 31668 33439 31720 33448
rect 31668 33405 31677 33439
rect 31677 33405 31711 33439
rect 31711 33405 31720 33439
rect 31668 33396 31720 33405
rect 33232 33328 33284 33380
rect 34428 33396 34480 33448
rect 36728 33396 36780 33448
rect 41972 33439 42024 33448
rect 41972 33405 41981 33439
rect 41981 33405 42015 33439
rect 42015 33405 42024 33439
rect 41972 33396 42024 33405
rect 40960 33328 41012 33380
rect 2228 33260 2280 33312
rect 2412 33303 2464 33312
rect 2412 33269 2421 33303
rect 2421 33269 2455 33303
rect 2455 33269 2464 33303
rect 2412 33260 2464 33269
rect 3332 33260 3384 33312
rect 4988 33303 5040 33312
rect 4988 33269 4997 33303
rect 4997 33269 5031 33303
rect 5031 33269 5040 33303
rect 4988 33260 5040 33269
rect 5816 33260 5868 33312
rect 8760 33303 8812 33312
rect 8760 33269 8769 33303
rect 8769 33269 8803 33303
rect 8803 33269 8812 33303
rect 8760 33260 8812 33269
rect 10692 33260 10744 33312
rect 10968 33303 11020 33312
rect 10968 33269 10977 33303
rect 10977 33269 11011 33303
rect 11011 33269 11020 33303
rect 10968 33260 11020 33269
rect 11520 33303 11572 33312
rect 11520 33269 11529 33303
rect 11529 33269 11563 33303
rect 11563 33269 11572 33303
rect 11520 33260 11572 33269
rect 13636 33303 13688 33312
rect 13636 33269 13645 33303
rect 13645 33269 13679 33303
rect 13679 33269 13688 33303
rect 13636 33260 13688 33269
rect 18144 33260 18196 33312
rect 26056 33260 26108 33312
rect 34244 33260 34296 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4620 33056 4672 33108
rect 5080 33056 5132 33108
rect 5448 33056 5500 33108
rect 6552 33056 6604 33108
rect 7012 33056 7064 33108
rect 9496 33099 9548 33108
rect 9496 33065 9505 33099
rect 9505 33065 9539 33099
rect 9539 33065 9548 33099
rect 9496 33056 9548 33065
rect 9588 33056 9640 33108
rect 4804 32988 4856 33040
rect 2780 32920 2832 32972
rect 4988 32920 5040 32972
rect 3332 32895 3384 32904
rect 3332 32861 3341 32895
rect 3341 32861 3375 32895
rect 3375 32861 3384 32895
rect 3332 32852 3384 32861
rect 2320 32784 2372 32836
rect 2872 32827 2924 32836
rect 2872 32793 2881 32827
rect 2881 32793 2915 32827
rect 2915 32793 2924 32827
rect 2872 32784 2924 32793
rect 2136 32716 2188 32768
rect 2504 32716 2556 32768
rect 4160 32827 4212 32836
rect 4160 32793 4169 32827
rect 4169 32793 4203 32827
rect 4203 32793 4212 32827
rect 4160 32784 4212 32793
rect 4712 32852 4764 32904
rect 5356 32920 5408 32972
rect 5908 32988 5960 33040
rect 8300 32920 8352 32972
rect 5632 32895 5684 32904
rect 5632 32861 5641 32895
rect 5641 32861 5675 32895
rect 5675 32861 5684 32895
rect 5632 32852 5684 32861
rect 7748 32895 7800 32904
rect 7748 32861 7757 32895
rect 7757 32861 7791 32895
rect 7791 32861 7800 32895
rect 7748 32852 7800 32861
rect 8760 32852 8812 32904
rect 10232 32920 10284 32972
rect 12348 33099 12400 33108
rect 12348 33065 12357 33099
rect 12357 33065 12391 33099
rect 12391 33065 12400 33099
rect 12348 33056 12400 33065
rect 13084 33056 13136 33108
rect 5080 32784 5132 32836
rect 5448 32784 5500 32836
rect 5908 32784 5960 32836
rect 7196 32827 7248 32836
rect 7196 32793 7205 32827
rect 7205 32793 7239 32827
rect 7239 32793 7248 32827
rect 7196 32784 7248 32793
rect 8116 32827 8168 32836
rect 8116 32793 8125 32827
rect 8125 32793 8159 32827
rect 8159 32793 8168 32827
rect 8116 32784 8168 32793
rect 8944 32784 8996 32836
rect 4436 32716 4488 32768
rect 4528 32716 4580 32768
rect 5540 32716 5592 32768
rect 9956 32895 10008 32904
rect 9956 32861 9991 32895
rect 9991 32861 10008 32895
rect 9956 32852 10008 32861
rect 10140 32895 10192 32904
rect 10140 32861 10149 32895
rect 10149 32861 10183 32895
rect 10183 32861 10192 32895
rect 10140 32852 10192 32861
rect 10692 32895 10744 32904
rect 10692 32861 10701 32895
rect 10701 32861 10735 32895
rect 10735 32861 10744 32895
rect 10692 32852 10744 32861
rect 10600 32827 10652 32836
rect 10600 32793 10609 32827
rect 10609 32793 10643 32827
rect 10643 32793 10652 32827
rect 11520 32852 11572 32904
rect 13820 32895 13872 32904
rect 13820 32861 13829 32895
rect 13829 32861 13863 32895
rect 13863 32861 13872 32895
rect 13820 32852 13872 32861
rect 10600 32784 10652 32793
rect 11336 32784 11388 32836
rect 13912 32784 13964 32836
rect 17224 33099 17276 33108
rect 17224 33065 17233 33099
rect 17233 33065 17267 33099
rect 17267 33065 17276 33099
rect 17224 33056 17276 33065
rect 18788 33056 18840 33108
rect 20904 33056 20956 33108
rect 21272 33056 21324 33108
rect 22744 33056 22796 33108
rect 23112 33056 23164 33108
rect 25228 33056 25280 33108
rect 26332 33056 26384 33108
rect 38292 33056 38344 33108
rect 15660 32988 15712 33040
rect 15476 32784 15528 32836
rect 15200 32716 15252 32768
rect 15844 32920 15896 32972
rect 16580 32920 16632 32972
rect 17040 32988 17092 33040
rect 16764 32963 16816 32972
rect 16764 32929 16773 32963
rect 16773 32929 16807 32963
rect 16807 32929 16816 32963
rect 16764 32920 16816 32929
rect 19616 32920 19668 32972
rect 17868 32852 17920 32904
rect 23020 32988 23072 33040
rect 28264 32988 28316 33040
rect 24400 32920 24452 32972
rect 19524 32784 19576 32836
rect 16028 32759 16080 32768
rect 16028 32725 16037 32759
rect 16037 32725 16071 32759
rect 16071 32725 16080 32759
rect 16028 32716 16080 32725
rect 17776 32716 17828 32768
rect 20076 32784 20128 32836
rect 21364 32784 21416 32836
rect 21456 32827 21508 32836
rect 21456 32793 21465 32827
rect 21465 32793 21499 32827
rect 21499 32793 21508 32827
rect 21456 32784 21508 32793
rect 25136 32895 25188 32904
rect 25136 32861 25145 32895
rect 25145 32861 25179 32895
rect 25179 32861 25188 32895
rect 25136 32852 25188 32861
rect 29736 32920 29788 32972
rect 33600 32920 33652 32972
rect 33968 32920 34020 32972
rect 34244 32963 34296 32972
rect 34244 32929 34253 32963
rect 34253 32929 34287 32963
rect 34287 32929 34296 32963
rect 34244 32920 34296 32929
rect 41236 33056 41288 33108
rect 27068 32852 27120 32904
rect 30656 32895 30708 32904
rect 30656 32861 30665 32895
rect 30665 32861 30699 32895
rect 30699 32861 30708 32895
rect 30656 32852 30708 32861
rect 34704 32852 34756 32904
rect 35440 32852 35492 32904
rect 37188 32852 37240 32904
rect 39672 32852 39724 32904
rect 40960 32852 41012 32904
rect 21732 32716 21784 32768
rect 25780 32784 25832 32836
rect 27436 32827 27488 32836
rect 27436 32793 27470 32827
rect 27470 32793 27488 32827
rect 27436 32784 27488 32793
rect 28080 32784 28132 32836
rect 32036 32784 32088 32836
rect 34336 32784 34388 32836
rect 34612 32784 34664 32836
rect 38108 32784 38160 32836
rect 23664 32716 23716 32768
rect 30104 32759 30156 32768
rect 30104 32725 30113 32759
rect 30113 32725 30147 32759
rect 30147 32725 30156 32759
rect 30104 32716 30156 32725
rect 32588 32759 32640 32768
rect 32588 32725 32597 32759
rect 32597 32725 32631 32759
rect 32631 32725 32640 32759
rect 32588 32716 32640 32725
rect 33692 32759 33744 32768
rect 33692 32725 33701 32759
rect 33701 32725 33735 32759
rect 33735 32725 33744 32759
rect 33692 32716 33744 32725
rect 34888 32716 34940 32768
rect 34980 32759 35032 32768
rect 34980 32725 34989 32759
rect 34989 32725 35023 32759
rect 35023 32725 35032 32759
rect 34980 32716 35032 32725
rect 38568 32759 38620 32768
rect 38568 32725 38577 32759
rect 38577 32725 38611 32759
rect 38611 32725 38620 32759
rect 38568 32716 38620 32725
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 2872 32512 2924 32564
rect 3240 32555 3292 32564
rect 3240 32521 3249 32555
rect 3249 32521 3283 32555
rect 3283 32521 3292 32555
rect 3240 32512 3292 32521
rect 4528 32512 4580 32564
rect 2412 32487 2464 32496
rect 2412 32453 2421 32487
rect 2421 32453 2455 32487
rect 2455 32453 2464 32487
rect 2412 32444 2464 32453
rect 4988 32512 5040 32564
rect 2228 32419 2280 32428
rect 2228 32385 2237 32419
rect 2237 32385 2271 32419
rect 2271 32385 2280 32419
rect 2228 32376 2280 32385
rect 2504 32419 2556 32428
rect 2504 32385 2513 32419
rect 2513 32385 2547 32419
rect 2547 32385 2556 32419
rect 2504 32376 2556 32385
rect 3148 32419 3200 32428
rect 3148 32385 3157 32419
rect 3157 32385 3191 32419
rect 3191 32385 3200 32419
rect 3148 32376 3200 32385
rect 3424 32376 3476 32428
rect 5356 32444 5408 32496
rect 5816 32512 5868 32564
rect 7196 32512 7248 32564
rect 8116 32512 8168 32564
rect 9956 32512 10008 32564
rect 21916 32512 21968 32564
rect 32128 32512 32180 32564
rect 34152 32555 34204 32564
rect 34152 32521 34161 32555
rect 34161 32521 34195 32555
rect 34195 32521 34204 32555
rect 34152 32512 34204 32521
rect 34796 32512 34848 32564
rect 34888 32512 34940 32564
rect 38660 32555 38712 32564
rect 38660 32521 38669 32555
rect 38669 32521 38703 32555
rect 38703 32521 38712 32555
rect 38660 32512 38712 32521
rect 40868 32512 40920 32564
rect 12164 32444 12216 32496
rect 16856 32487 16908 32496
rect 16856 32453 16865 32487
rect 16865 32453 16899 32487
rect 16899 32453 16908 32487
rect 16856 32444 16908 32453
rect 18144 32487 18196 32496
rect 18144 32453 18153 32487
rect 18153 32453 18187 32487
rect 18187 32453 18196 32487
rect 18144 32444 18196 32453
rect 4804 32376 4856 32428
rect 4988 32419 5040 32428
rect 4988 32385 4997 32419
rect 4997 32385 5031 32419
rect 5031 32385 5040 32419
rect 4988 32376 5040 32385
rect 5448 32419 5500 32428
rect 5448 32385 5457 32419
rect 5457 32385 5491 32419
rect 5491 32385 5500 32419
rect 5448 32376 5500 32385
rect 3700 32351 3752 32360
rect 3700 32317 3709 32351
rect 3709 32317 3743 32351
rect 3743 32317 3752 32351
rect 3700 32308 3752 32317
rect 4712 32308 4764 32360
rect 5080 32351 5132 32360
rect 5080 32317 5089 32351
rect 5089 32317 5123 32351
rect 5123 32317 5132 32351
rect 5080 32308 5132 32317
rect 6276 32376 6328 32428
rect 3332 32240 3384 32292
rect 4068 32172 4120 32224
rect 5540 32240 5592 32292
rect 4712 32215 4764 32224
rect 4712 32181 4721 32215
rect 4721 32181 4755 32215
rect 4755 32181 4764 32215
rect 4712 32172 4764 32181
rect 4988 32172 5040 32224
rect 5264 32172 5316 32224
rect 6000 32308 6052 32360
rect 6092 32308 6144 32360
rect 6460 32376 6512 32428
rect 9864 32376 9916 32428
rect 10600 32376 10652 32428
rect 13912 32419 13964 32428
rect 13912 32385 13921 32419
rect 13921 32385 13955 32419
rect 13955 32385 13964 32419
rect 13912 32376 13964 32385
rect 15568 32376 15620 32428
rect 16396 32376 16448 32428
rect 17868 32419 17920 32428
rect 17868 32385 17877 32419
rect 17877 32385 17911 32419
rect 17911 32385 17920 32419
rect 17868 32376 17920 32385
rect 8668 32308 8720 32360
rect 14464 32351 14516 32360
rect 14464 32317 14473 32351
rect 14473 32317 14507 32351
rect 14507 32317 14516 32351
rect 14464 32308 14516 32317
rect 18604 32308 18656 32360
rect 20076 32444 20128 32496
rect 20628 32487 20680 32496
rect 20628 32453 20637 32487
rect 20637 32453 20671 32487
rect 20671 32453 20680 32487
rect 20628 32444 20680 32453
rect 20812 32444 20864 32496
rect 21364 32487 21416 32496
rect 21364 32453 21373 32487
rect 21373 32453 21407 32487
rect 21407 32453 21416 32487
rect 21364 32444 21416 32453
rect 22376 32444 22428 32496
rect 23020 32444 23072 32496
rect 24032 32444 24084 32496
rect 26056 32444 26108 32496
rect 26332 32444 26384 32496
rect 20536 32419 20588 32428
rect 20536 32385 20545 32419
rect 20545 32385 20579 32419
rect 20579 32385 20588 32419
rect 20536 32376 20588 32385
rect 20720 32419 20772 32428
rect 20720 32385 20729 32419
rect 20729 32385 20763 32419
rect 20763 32385 20772 32419
rect 20720 32376 20772 32385
rect 20904 32419 20956 32428
rect 20904 32385 20913 32419
rect 20913 32385 20947 32419
rect 20947 32385 20956 32419
rect 20904 32376 20956 32385
rect 19708 32308 19760 32360
rect 21824 32376 21876 32428
rect 22744 32376 22796 32428
rect 24308 32419 24360 32428
rect 24308 32385 24317 32419
rect 24317 32385 24351 32419
rect 24351 32385 24360 32419
rect 24308 32376 24360 32385
rect 24584 32419 24636 32428
rect 24584 32385 24593 32419
rect 24593 32385 24627 32419
rect 24627 32385 24636 32419
rect 24584 32376 24636 32385
rect 25596 32419 25648 32428
rect 25596 32385 25605 32419
rect 25605 32385 25639 32419
rect 25639 32385 25648 32419
rect 25596 32376 25648 32385
rect 27160 32376 27212 32428
rect 28080 32419 28132 32428
rect 28080 32385 28089 32419
rect 28089 32385 28123 32419
rect 28123 32385 28132 32419
rect 28080 32376 28132 32385
rect 28816 32444 28868 32496
rect 29736 32444 29788 32496
rect 30104 32444 30156 32496
rect 6552 32283 6604 32292
rect 6552 32249 6561 32283
rect 6561 32249 6595 32283
rect 6595 32249 6604 32283
rect 6552 32240 6604 32249
rect 13176 32240 13228 32292
rect 9588 32172 9640 32224
rect 15108 32172 15160 32224
rect 20720 32240 20772 32292
rect 23664 32308 23716 32360
rect 26056 32308 26108 32360
rect 25780 32283 25832 32292
rect 25780 32249 25789 32283
rect 25789 32249 25823 32283
rect 25823 32249 25832 32283
rect 25780 32240 25832 32249
rect 27436 32240 27488 32292
rect 16120 32172 16172 32224
rect 22008 32172 22060 32224
rect 22560 32215 22612 32224
rect 22560 32181 22569 32215
rect 22569 32181 22603 32215
rect 22603 32181 22612 32215
rect 22560 32172 22612 32181
rect 25044 32215 25096 32224
rect 25044 32181 25053 32215
rect 25053 32181 25087 32215
rect 25087 32181 25096 32215
rect 25044 32172 25096 32181
rect 30196 32376 30248 32428
rect 31484 32376 31536 32428
rect 33324 32376 33376 32428
rect 34980 32444 35032 32496
rect 37372 32376 37424 32428
rect 39672 32419 39724 32428
rect 39672 32385 39681 32419
rect 39681 32385 39715 32419
rect 39715 32385 39724 32419
rect 39672 32376 39724 32385
rect 39948 32419 40000 32428
rect 39948 32385 39982 32419
rect 39982 32385 40000 32419
rect 39948 32376 40000 32385
rect 42156 32376 42208 32428
rect 32772 32351 32824 32360
rect 32772 32317 32781 32351
rect 32781 32317 32815 32351
rect 32815 32317 32824 32351
rect 32772 32308 32824 32317
rect 30288 32240 30340 32292
rect 37280 32351 37332 32360
rect 37280 32317 37289 32351
rect 37289 32317 37323 32351
rect 37323 32317 37332 32351
rect 37280 32308 37332 32317
rect 29184 32172 29236 32224
rect 30656 32172 30708 32224
rect 31024 32215 31076 32224
rect 31024 32181 31033 32215
rect 31033 32181 31067 32215
rect 31067 32181 31076 32215
rect 31024 32172 31076 32181
rect 34428 32172 34480 32224
rect 35532 32172 35584 32224
rect 37924 32172 37976 32224
rect 38752 32215 38804 32224
rect 38752 32181 38761 32215
rect 38761 32181 38795 32215
rect 38795 32181 38804 32215
rect 38752 32172 38804 32181
rect 41144 32215 41196 32224
rect 41144 32181 41153 32215
rect 41153 32181 41187 32215
rect 41187 32181 41196 32215
rect 41144 32172 41196 32181
rect 42064 32215 42116 32224
rect 42064 32181 42073 32215
rect 42073 32181 42107 32215
rect 42107 32181 42116 32215
rect 42064 32172 42116 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4620 32011 4672 32020
rect 4620 31977 4629 32011
rect 4629 31977 4663 32011
rect 4663 31977 4672 32011
rect 4620 31968 4672 31977
rect 3700 31900 3752 31952
rect 5172 31968 5224 32020
rect 5356 31968 5408 32020
rect 5632 32011 5684 32020
rect 5632 31977 5641 32011
rect 5641 31977 5675 32011
rect 5675 31977 5684 32011
rect 5632 31968 5684 31977
rect 7656 31968 7708 32020
rect 11520 31968 11572 32020
rect 14464 31968 14516 32020
rect 15476 32011 15528 32020
rect 15476 31977 15485 32011
rect 15485 31977 15519 32011
rect 15519 31977 15528 32011
rect 15476 31968 15528 31977
rect 15568 32011 15620 32020
rect 15568 31977 15577 32011
rect 15577 31977 15611 32011
rect 15611 31977 15620 32011
rect 15568 31968 15620 31977
rect 3332 31832 3384 31884
rect 3976 31832 4028 31884
rect 6276 31832 6328 31884
rect 2872 31764 2924 31816
rect 4804 31807 4856 31816
rect 4804 31773 4813 31807
rect 4813 31773 4847 31807
rect 4847 31773 4856 31807
rect 4804 31764 4856 31773
rect 5080 31764 5132 31816
rect 5356 31764 5408 31816
rect 6460 31764 6512 31816
rect 6644 31764 6696 31816
rect 8300 31832 8352 31884
rect 13176 31875 13228 31884
rect 13176 31841 13185 31875
rect 13185 31841 13219 31875
rect 13219 31841 13228 31875
rect 13176 31832 13228 31841
rect 13636 31832 13688 31884
rect 16396 31968 16448 32020
rect 17776 31968 17828 32020
rect 20352 31968 20404 32020
rect 20536 31968 20588 32020
rect 21456 31968 21508 32020
rect 22560 31968 22612 32020
rect 23480 31968 23532 32020
rect 24032 32011 24084 32020
rect 24032 31977 24041 32011
rect 24041 31977 24075 32011
rect 24075 31977 24084 32011
rect 24032 31968 24084 31977
rect 21548 31900 21600 31952
rect 25596 31968 25648 32020
rect 27252 32011 27304 32020
rect 27252 31977 27261 32011
rect 27261 31977 27295 32011
rect 27295 31977 27304 32011
rect 27252 31968 27304 31977
rect 28724 31943 28776 31952
rect 28724 31909 28733 31943
rect 28733 31909 28767 31943
rect 28767 31909 28776 31943
rect 28724 31900 28776 31909
rect 10508 31764 10560 31816
rect 5264 31739 5316 31748
rect 5264 31705 5273 31739
rect 5273 31705 5307 31739
rect 5307 31705 5316 31739
rect 5264 31696 5316 31705
rect 7012 31739 7064 31748
rect 7012 31705 7021 31739
rect 7021 31705 7055 31739
rect 7055 31705 7064 31739
rect 7012 31696 7064 31705
rect 9404 31739 9456 31748
rect 9404 31705 9413 31739
rect 9413 31705 9447 31739
rect 9447 31705 9456 31739
rect 9404 31696 9456 31705
rect 11612 31764 11664 31816
rect 12164 31764 12216 31816
rect 13820 31764 13872 31816
rect 16028 31807 16080 31816
rect 16028 31773 16037 31807
rect 16037 31773 16071 31807
rect 16071 31773 16080 31807
rect 16028 31764 16080 31773
rect 16120 31764 16172 31816
rect 16396 31875 16448 31884
rect 16396 31841 16405 31875
rect 16405 31841 16439 31875
rect 16439 31841 16448 31875
rect 16396 31832 16448 31841
rect 19708 31832 19760 31884
rect 20628 31832 20680 31884
rect 22376 31832 22428 31884
rect 22744 31832 22796 31884
rect 22008 31764 22060 31816
rect 14464 31696 14516 31748
rect 16580 31696 16632 31748
rect 16672 31739 16724 31748
rect 16672 31705 16681 31739
rect 16681 31705 16715 31739
rect 16715 31705 16724 31739
rect 16672 31696 16724 31705
rect 18144 31696 18196 31748
rect 18604 31696 18656 31748
rect 19340 31696 19392 31748
rect 22100 31739 22152 31748
rect 22100 31705 22109 31739
rect 22109 31705 22143 31739
rect 22143 31705 22152 31739
rect 22100 31696 22152 31705
rect 23480 31807 23532 31816
rect 23480 31773 23489 31807
rect 23489 31773 23523 31807
rect 23523 31773 23532 31807
rect 23480 31764 23532 31773
rect 23664 31807 23716 31816
rect 23664 31773 23673 31807
rect 23673 31773 23707 31807
rect 23707 31773 23716 31807
rect 23664 31764 23716 31773
rect 25780 31764 25832 31816
rect 27068 31764 27120 31816
rect 28816 31764 28868 31816
rect 24032 31696 24084 31748
rect 24860 31696 24912 31748
rect 26148 31739 26200 31748
rect 26148 31705 26182 31739
rect 26182 31705 26200 31739
rect 26148 31696 26200 31705
rect 27712 31696 27764 31748
rect 31484 31968 31536 32020
rect 33968 31968 34020 32020
rect 34428 32011 34480 32020
rect 34428 31977 34437 32011
rect 34437 31977 34471 32011
rect 34471 31977 34480 32011
rect 34428 31968 34480 31977
rect 37372 31968 37424 32020
rect 38108 32011 38160 32020
rect 38108 31977 38117 32011
rect 38117 31977 38151 32011
rect 38151 31977 38160 32011
rect 38108 31968 38160 31977
rect 39948 31968 40000 32020
rect 31208 31943 31260 31952
rect 31208 31909 31217 31943
rect 31217 31909 31251 31943
rect 31251 31909 31260 31943
rect 31208 31900 31260 31909
rect 31576 31900 31628 31952
rect 34796 31832 34848 31884
rect 38752 31900 38804 31952
rect 29000 31764 29052 31816
rect 30380 31764 30432 31816
rect 31760 31764 31812 31816
rect 32772 31764 32824 31816
rect 33692 31764 33744 31816
rect 38568 31875 38620 31884
rect 38568 31841 38577 31875
rect 38577 31841 38611 31875
rect 38611 31841 38620 31875
rect 38568 31832 38620 31841
rect 39488 31832 39540 31884
rect 41144 31900 41196 31952
rect 38936 31764 38988 31816
rect 39948 31764 40000 31816
rect 40684 31832 40736 31884
rect 40500 31764 40552 31816
rect 40776 31807 40828 31816
rect 40776 31773 40785 31807
rect 40785 31773 40819 31807
rect 40819 31773 40828 31807
rect 40776 31764 40828 31773
rect 41420 31807 41472 31816
rect 41420 31773 41429 31807
rect 41429 31773 41463 31807
rect 41463 31773 41472 31807
rect 41420 31764 41472 31773
rect 42156 31807 42208 31816
rect 42156 31773 42165 31807
rect 42165 31773 42199 31807
rect 42199 31773 42208 31807
rect 42156 31764 42208 31773
rect 29184 31696 29236 31748
rect 30288 31696 30340 31748
rect 31944 31696 31996 31748
rect 35348 31739 35400 31748
rect 35348 31705 35357 31739
rect 35357 31705 35391 31739
rect 35391 31705 35400 31739
rect 35348 31696 35400 31705
rect 3332 31671 3384 31680
rect 3332 31637 3341 31671
rect 3341 31637 3375 31671
rect 3375 31637 3384 31671
rect 3332 31628 3384 31637
rect 5172 31628 5224 31680
rect 8484 31671 8536 31680
rect 8484 31637 8493 31671
rect 8493 31637 8527 31671
rect 8527 31637 8536 31671
rect 8484 31628 8536 31637
rect 10416 31628 10468 31680
rect 10876 31671 10928 31680
rect 10876 31637 10885 31671
rect 10885 31637 10919 31671
rect 10919 31637 10928 31671
rect 10876 31628 10928 31637
rect 10968 31671 11020 31680
rect 10968 31637 10977 31671
rect 10977 31637 11011 31671
rect 11011 31637 11020 31671
rect 10968 31628 11020 31637
rect 13452 31671 13504 31680
rect 13452 31637 13461 31671
rect 13461 31637 13495 31671
rect 13495 31637 13504 31671
rect 13452 31628 13504 31637
rect 15936 31671 15988 31680
rect 15936 31637 15945 31671
rect 15945 31637 15979 31671
rect 15979 31637 15988 31671
rect 15936 31628 15988 31637
rect 17592 31628 17644 31680
rect 19524 31671 19576 31680
rect 19524 31637 19533 31671
rect 19533 31637 19567 31671
rect 19567 31637 19576 31671
rect 19524 31628 19576 31637
rect 28816 31628 28868 31680
rect 29000 31628 29052 31680
rect 33508 31628 33560 31680
rect 36820 31671 36872 31680
rect 36820 31637 36829 31671
rect 36829 31637 36863 31671
rect 36863 31637 36872 31671
rect 36820 31628 36872 31637
rect 38476 31671 38528 31680
rect 38476 31637 38485 31671
rect 38485 31637 38519 31671
rect 38519 31637 38528 31671
rect 38476 31628 38528 31637
rect 38660 31628 38712 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 4068 31424 4120 31476
rect 6184 31424 6236 31476
rect 7012 31424 7064 31476
rect 2412 31356 2464 31408
rect 5908 31356 5960 31408
rect 8668 31424 8720 31476
rect 9128 31424 9180 31476
rect 9404 31424 9456 31476
rect 14464 31467 14516 31476
rect 14464 31433 14473 31467
rect 14473 31433 14507 31467
rect 14507 31433 14516 31467
rect 14464 31424 14516 31433
rect 15936 31424 15988 31476
rect 16488 31424 16540 31476
rect 17592 31424 17644 31476
rect 8116 31356 8168 31408
rect 8208 31356 8260 31408
rect 3056 31288 3108 31340
rect 3700 31288 3752 31340
rect 8760 31356 8812 31408
rect 9588 31399 9640 31408
rect 9588 31365 9597 31399
rect 9597 31365 9631 31399
rect 9631 31365 9640 31399
rect 9588 31356 9640 31365
rect 2044 31220 2096 31272
rect 3240 31220 3292 31272
rect 4712 31220 4764 31272
rect 7840 31220 7892 31272
rect 1400 31084 1452 31136
rect 2688 31084 2740 31136
rect 2964 31084 3016 31136
rect 8484 31152 8536 31204
rect 4620 31084 4672 31136
rect 5632 31084 5684 31136
rect 9496 31331 9548 31340
rect 9496 31297 9505 31331
rect 9505 31297 9539 31331
rect 9539 31297 9548 31331
rect 9496 31288 9548 31297
rect 9128 31220 9180 31272
rect 9956 31356 10008 31408
rect 12900 31356 12952 31408
rect 15384 31356 15436 31408
rect 21548 31424 21600 31476
rect 21640 31424 21692 31476
rect 22192 31424 22244 31476
rect 23296 31424 23348 31476
rect 24860 31467 24912 31476
rect 24860 31433 24869 31467
rect 24869 31433 24903 31467
rect 24903 31433 24912 31467
rect 24860 31424 24912 31433
rect 25044 31424 25096 31476
rect 26148 31424 26200 31476
rect 30380 31467 30432 31476
rect 30380 31433 30389 31467
rect 30389 31433 30423 31467
rect 30423 31433 30432 31467
rect 30380 31424 30432 31433
rect 31024 31424 31076 31476
rect 31944 31424 31996 31476
rect 32036 31424 32088 31476
rect 32588 31467 32640 31476
rect 32588 31433 32597 31467
rect 32597 31433 32631 31467
rect 32631 31433 32640 31467
rect 32588 31424 32640 31433
rect 33324 31467 33376 31476
rect 33324 31433 33333 31467
rect 33333 31433 33367 31467
rect 33367 31433 33376 31467
rect 33324 31424 33376 31433
rect 33784 31424 33836 31476
rect 41052 31467 41104 31476
rect 41052 31433 41061 31467
rect 41061 31433 41095 31467
rect 41095 31433 41104 31467
rect 41052 31424 41104 31433
rect 19156 31356 19208 31408
rect 23388 31356 23440 31408
rect 10968 31288 11020 31340
rect 13452 31288 13504 31340
rect 10232 31263 10284 31272
rect 10232 31229 10241 31263
rect 10241 31229 10275 31263
rect 10275 31229 10284 31263
rect 10232 31220 10284 31229
rect 9772 31152 9824 31204
rect 9864 31152 9916 31204
rect 10140 31152 10192 31204
rect 10416 31263 10468 31272
rect 10416 31229 10425 31263
rect 10425 31229 10459 31263
rect 10459 31229 10468 31263
rect 10416 31220 10468 31229
rect 10876 31220 10928 31272
rect 11612 31263 11664 31272
rect 11612 31229 11621 31263
rect 11621 31229 11655 31263
rect 11655 31229 11664 31263
rect 11612 31220 11664 31229
rect 12624 31220 12676 31272
rect 12992 31152 13044 31204
rect 15476 31288 15528 31340
rect 16580 31220 16632 31272
rect 16856 31263 16908 31272
rect 16856 31229 16865 31263
rect 16865 31229 16899 31263
rect 16899 31229 16908 31263
rect 16856 31220 16908 31229
rect 18144 31288 18196 31340
rect 19616 31288 19668 31340
rect 21180 31288 21232 31340
rect 22284 31288 22336 31340
rect 24124 31288 24176 31340
rect 25228 31331 25280 31340
rect 25228 31297 25237 31331
rect 25237 31297 25271 31331
rect 25271 31297 25280 31331
rect 25228 31288 25280 31297
rect 16580 31084 16632 31136
rect 16856 31084 16908 31136
rect 19708 31220 19760 31272
rect 24216 31220 24268 31272
rect 26792 31356 26844 31408
rect 28356 31356 28408 31408
rect 27252 31288 27304 31340
rect 28816 31331 28868 31340
rect 28816 31297 28825 31331
rect 28825 31297 28859 31331
rect 28859 31297 28868 31331
rect 28816 31288 28868 31297
rect 26056 31220 26108 31272
rect 28172 31263 28224 31272
rect 28172 31229 28181 31263
rect 28181 31229 28215 31263
rect 28215 31229 28224 31263
rect 28172 31220 28224 31229
rect 29184 31356 29236 31408
rect 29460 31356 29512 31408
rect 30196 31356 30248 31408
rect 33140 31356 33192 31408
rect 37924 31356 37976 31408
rect 29552 31288 29604 31340
rect 32404 31288 32456 31340
rect 32680 31288 32732 31340
rect 34244 31288 34296 31340
rect 30288 31152 30340 31204
rect 31668 31263 31720 31272
rect 31668 31229 31677 31263
rect 31677 31229 31711 31263
rect 31711 31229 31720 31263
rect 31668 31220 31720 31229
rect 33048 31220 33100 31272
rect 33968 31263 34020 31272
rect 33968 31229 33977 31263
rect 33977 31229 34011 31263
rect 34011 31229 34020 31263
rect 33968 31220 34020 31229
rect 39672 31331 39724 31340
rect 39672 31297 39688 31331
rect 39688 31297 39722 31331
rect 39722 31297 39724 31331
rect 40408 31356 40460 31408
rect 39672 31288 39724 31297
rect 40960 31288 41012 31340
rect 17408 31127 17460 31136
rect 17408 31093 17417 31127
rect 17417 31093 17451 31127
rect 17451 31093 17460 31127
rect 17408 31084 17460 31093
rect 18236 31084 18288 31136
rect 21824 31084 21876 31136
rect 22652 31084 22704 31136
rect 24032 31084 24084 31136
rect 28264 31084 28316 31136
rect 30932 31084 30984 31136
rect 39488 31084 39540 31136
rect 40040 31084 40092 31136
rect 41236 31127 41288 31136
rect 41236 31093 41245 31127
rect 41245 31093 41279 31127
rect 41279 31093 41288 31127
rect 41236 31084 41288 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2872 30880 2924 30932
rect 4712 30880 4764 30932
rect 5172 30880 5224 30932
rect 5816 30880 5868 30932
rect 7840 30923 7892 30932
rect 7840 30889 7849 30923
rect 7849 30889 7883 30923
rect 7883 30889 7892 30923
rect 7840 30880 7892 30889
rect 8760 30880 8812 30932
rect 10232 30880 10284 30932
rect 12624 30923 12676 30932
rect 12624 30889 12633 30923
rect 12633 30889 12667 30923
rect 12667 30889 12676 30923
rect 12624 30880 12676 30889
rect 16672 30880 16724 30932
rect 2596 30812 2648 30864
rect 2044 30787 2096 30796
rect 2044 30753 2053 30787
rect 2053 30753 2087 30787
rect 2087 30753 2096 30787
rect 2044 30744 2096 30753
rect 2964 30744 3016 30796
rect 3056 30787 3108 30796
rect 3056 30753 3065 30787
rect 3065 30753 3099 30787
rect 3099 30753 3108 30787
rect 3056 30744 3108 30753
rect 3424 30744 3476 30796
rect 5448 30812 5500 30864
rect 5724 30812 5776 30864
rect 4804 30744 4856 30796
rect 1584 30651 1636 30660
rect 1584 30617 1593 30651
rect 1593 30617 1627 30651
rect 1627 30617 1636 30651
rect 1584 30608 1636 30617
rect 3240 30719 3292 30728
rect 3240 30685 3249 30719
rect 3249 30685 3283 30719
rect 3283 30685 3292 30719
rect 3240 30676 3292 30685
rect 1860 30608 1912 30660
rect 2412 30651 2464 30660
rect 2412 30617 2421 30651
rect 2421 30617 2455 30651
rect 2455 30617 2464 30651
rect 2412 30608 2464 30617
rect 2964 30608 3016 30660
rect 3884 30608 3936 30660
rect 3332 30540 3384 30592
rect 4620 30676 4672 30728
rect 6644 30744 6696 30796
rect 13360 30744 13412 30796
rect 5172 30676 5224 30728
rect 5724 30676 5776 30728
rect 5816 30719 5868 30728
rect 5816 30685 5825 30719
rect 5825 30685 5859 30719
rect 5859 30685 5868 30719
rect 5816 30676 5868 30685
rect 6184 30719 6236 30728
rect 6184 30685 6193 30719
rect 6193 30685 6227 30719
rect 6227 30685 6236 30719
rect 6184 30676 6236 30685
rect 8484 30719 8536 30728
rect 4712 30608 4764 30660
rect 8484 30685 8493 30719
rect 8493 30685 8527 30719
rect 8527 30685 8536 30719
rect 8484 30676 8536 30685
rect 8760 30719 8812 30728
rect 8760 30685 8769 30719
rect 8769 30685 8803 30719
rect 8803 30685 8812 30719
rect 8760 30676 8812 30685
rect 12992 30719 13044 30728
rect 12992 30685 13001 30719
rect 13001 30685 13035 30719
rect 13035 30685 13044 30719
rect 12992 30676 13044 30685
rect 13452 30719 13504 30728
rect 13452 30685 13461 30719
rect 13461 30685 13495 30719
rect 13495 30685 13504 30719
rect 13452 30676 13504 30685
rect 13544 30676 13596 30728
rect 17224 30719 17276 30728
rect 17224 30685 17233 30719
rect 17233 30685 17267 30719
rect 17267 30685 17276 30719
rect 17224 30676 17276 30685
rect 17500 30787 17552 30796
rect 17500 30753 17509 30787
rect 17509 30753 17543 30787
rect 17543 30753 17552 30787
rect 19892 30880 19944 30932
rect 21548 30880 21600 30932
rect 22100 30923 22152 30932
rect 22100 30889 22109 30923
rect 22109 30889 22143 30923
rect 22143 30889 22152 30923
rect 22100 30880 22152 30889
rect 24584 30880 24636 30932
rect 18880 30812 18932 30864
rect 19708 30812 19760 30864
rect 17500 30744 17552 30753
rect 17868 30676 17920 30728
rect 19432 30744 19484 30796
rect 20260 30812 20312 30864
rect 19892 30787 19944 30796
rect 19892 30753 19901 30787
rect 19901 30753 19935 30787
rect 19935 30753 19944 30787
rect 19892 30744 19944 30753
rect 19984 30744 20036 30796
rect 22192 30812 22244 30864
rect 23664 30812 23716 30864
rect 27712 30923 27764 30932
rect 27712 30889 27721 30923
rect 27721 30889 27755 30923
rect 27755 30889 27764 30923
rect 27712 30880 27764 30889
rect 28172 30880 28224 30932
rect 29552 30923 29604 30932
rect 29552 30889 29561 30923
rect 29561 30889 29595 30923
rect 29595 30889 29604 30923
rect 29552 30880 29604 30889
rect 31668 30880 31720 30932
rect 35348 30880 35400 30932
rect 38844 30880 38896 30932
rect 39488 30880 39540 30932
rect 41420 30880 41472 30932
rect 41788 30880 41840 30932
rect 8208 30608 8260 30660
rect 5816 30540 5868 30592
rect 6552 30540 6604 30592
rect 8668 30583 8720 30592
rect 8668 30549 8677 30583
rect 8677 30549 8711 30583
rect 8711 30549 8720 30583
rect 8668 30540 8720 30549
rect 9220 30651 9272 30660
rect 9220 30617 9229 30651
rect 9229 30617 9263 30651
rect 9263 30617 9272 30651
rect 9220 30608 9272 30617
rect 10508 30608 10560 30660
rect 10968 30608 11020 30660
rect 18052 30608 18104 30660
rect 18788 30676 18840 30728
rect 19064 30676 19116 30728
rect 19616 30676 19668 30728
rect 19708 30676 19760 30728
rect 20628 30744 20680 30796
rect 19892 30608 19944 30660
rect 20444 30719 20496 30728
rect 20444 30685 20453 30719
rect 20453 30685 20487 30719
rect 20487 30685 20496 30719
rect 20444 30676 20496 30685
rect 20536 30719 20588 30728
rect 20536 30685 20550 30719
rect 20550 30685 20584 30719
rect 20584 30685 20588 30719
rect 20536 30676 20588 30685
rect 10140 30540 10192 30592
rect 13176 30540 13228 30592
rect 15200 30540 15252 30592
rect 17592 30540 17644 30592
rect 18420 30540 18472 30592
rect 19156 30540 19208 30592
rect 19524 30540 19576 30592
rect 21088 30676 21140 30728
rect 22008 30676 22060 30728
rect 21824 30651 21876 30660
rect 21824 30617 21833 30651
rect 21833 30617 21867 30651
rect 21867 30617 21876 30651
rect 21824 30608 21876 30617
rect 22468 30608 22520 30660
rect 23388 30676 23440 30728
rect 25688 30744 25740 30796
rect 25780 30787 25832 30796
rect 25780 30753 25789 30787
rect 25789 30753 25823 30787
rect 25823 30753 25832 30787
rect 25780 30744 25832 30753
rect 28264 30787 28316 30796
rect 28264 30753 28273 30787
rect 28273 30753 28307 30787
rect 28307 30753 28316 30787
rect 28264 30744 28316 30753
rect 28724 30744 28776 30796
rect 30288 30744 30340 30796
rect 30932 30787 30984 30796
rect 30932 30753 30941 30787
rect 30941 30753 30975 30787
rect 30975 30753 30984 30787
rect 30932 30744 30984 30753
rect 31208 30744 31260 30796
rect 31760 30744 31812 30796
rect 23572 30719 23624 30728
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 25320 30676 25372 30728
rect 33416 30676 33468 30728
rect 22008 30540 22060 30592
rect 22376 30540 22428 30592
rect 28632 30608 28684 30660
rect 30104 30608 30156 30660
rect 32312 30651 32364 30660
rect 32312 30617 32321 30651
rect 32321 30617 32355 30651
rect 32355 30617 32364 30651
rect 32312 30608 32364 30617
rect 26240 30540 26292 30592
rect 26792 30540 26844 30592
rect 33140 30540 33192 30592
rect 35716 30787 35768 30796
rect 35716 30753 35725 30787
rect 35725 30753 35759 30787
rect 35759 30753 35768 30787
rect 35716 30744 35768 30753
rect 35072 30676 35124 30728
rect 35532 30719 35584 30728
rect 35532 30685 35541 30719
rect 35541 30685 35575 30719
rect 35575 30685 35584 30719
rect 35532 30676 35584 30685
rect 35348 30608 35400 30660
rect 36820 30676 36872 30728
rect 37740 30676 37792 30728
rect 37924 30676 37976 30728
rect 40684 30744 40736 30796
rect 40132 30719 40184 30728
rect 40132 30685 40141 30719
rect 40141 30685 40175 30719
rect 40175 30685 40184 30719
rect 40132 30676 40184 30685
rect 40408 30719 40460 30728
rect 40408 30685 40417 30719
rect 40417 30685 40451 30719
rect 40451 30685 40460 30719
rect 40408 30676 40460 30685
rect 38200 30608 38252 30660
rect 38292 30608 38344 30660
rect 39856 30540 39908 30592
rect 40316 30583 40368 30592
rect 40316 30549 40325 30583
rect 40325 30549 40359 30583
rect 40359 30549 40368 30583
rect 40316 30540 40368 30549
rect 40684 30651 40736 30660
rect 40684 30617 40693 30651
rect 40693 30617 40727 30651
rect 40727 30617 40736 30651
rect 40684 30608 40736 30617
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 2412 30379 2464 30388
rect 2412 30345 2421 30379
rect 2421 30345 2455 30379
rect 2455 30345 2464 30379
rect 2412 30336 2464 30345
rect 1860 30268 1912 30320
rect 2596 30243 2648 30252
rect 2596 30209 2605 30243
rect 2605 30209 2639 30243
rect 2639 30209 2648 30243
rect 2596 30200 2648 30209
rect 4068 30336 4120 30388
rect 5816 30379 5868 30388
rect 5816 30345 5825 30379
rect 5825 30345 5859 30379
rect 5859 30345 5868 30379
rect 5816 30336 5868 30345
rect 9220 30336 9272 30388
rect 16488 30379 16540 30388
rect 16488 30345 16497 30379
rect 16497 30345 16531 30379
rect 16531 30345 16540 30379
rect 16488 30336 16540 30345
rect 3240 30311 3292 30320
rect 3240 30277 3249 30311
rect 3249 30277 3283 30311
rect 3283 30277 3292 30311
rect 3240 30268 3292 30277
rect 4160 30268 4212 30320
rect 4620 30311 4672 30320
rect 4620 30277 4629 30311
rect 4629 30277 4663 30311
rect 4663 30277 4672 30311
rect 4620 30268 4672 30277
rect 5448 30311 5500 30320
rect 5448 30277 5457 30311
rect 5457 30277 5491 30311
rect 5491 30277 5500 30311
rect 5448 30268 5500 30277
rect 8668 30268 8720 30320
rect 1584 30132 1636 30184
rect 2504 30132 2556 30184
rect 3608 30132 3660 30184
rect 5264 30200 5316 30252
rect 6552 30243 6604 30252
rect 6552 30209 6561 30243
rect 6561 30209 6595 30243
rect 6595 30209 6604 30243
rect 6552 30200 6604 30209
rect 6828 30243 6880 30252
rect 6828 30209 6837 30243
rect 6837 30209 6871 30243
rect 6871 30209 6880 30243
rect 6828 30200 6880 30209
rect 9036 30243 9088 30252
rect 9036 30209 9045 30243
rect 9045 30209 9079 30243
rect 9079 30209 9088 30243
rect 9036 30200 9088 30209
rect 9220 30243 9272 30252
rect 9220 30209 9229 30243
rect 9229 30209 9263 30243
rect 9263 30209 9272 30243
rect 9220 30200 9272 30209
rect 5540 30132 5592 30184
rect 5632 30175 5684 30184
rect 5632 30141 5641 30175
rect 5641 30141 5675 30175
rect 5675 30141 5684 30175
rect 5632 30132 5684 30141
rect 5724 30175 5776 30184
rect 5724 30141 5733 30175
rect 5733 30141 5767 30175
rect 5767 30141 5776 30175
rect 5724 30132 5776 30141
rect 6000 30175 6052 30184
rect 6000 30141 6009 30175
rect 6009 30141 6043 30175
rect 6043 30141 6052 30175
rect 6000 30132 6052 30141
rect 6184 30132 6236 30184
rect 6276 30132 6328 30184
rect 10232 30200 10284 30252
rect 11612 30243 11664 30252
rect 11612 30209 11621 30243
rect 11621 30209 11655 30243
rect 11655 30209 11664 30243
rect 11612 30200 11664 30209
rect 12992 30200 13044 30252
rect 13544 30243 13596 30252
rect 13544 30209 13553 30243
rect 13553 30209 13587 30243
rect 13587 30209 13596 30243
rect 13544 30200 13596 30209
rect 13912 30200 13964 30252
rect 14924 30268 14976 30320
rect 16672 30268 16724 30320
rect 17224 30336 17276 30388
rect 19432 30336 19484 30388
rect 19616 30336 19668 30388
rect 19984 30336 20036 30388
rect 13084 30132 13136 30184
rect 13820 30132 13872 30184
rect 17592 30243 17644 30252
rect 17592 30209 17601 30243
rect 17601 30209 17635 30243
rect 17635 30209 17644 30243
rect 17592 30200 17644 30209
rect 17684 30243 17736 30252
rect 17684 30209 17693 30243
rect 17693 30209 17727 30243
rect 17727 30209 17736 30243
rect 17684 30200 17736 30209
rect 17868 30200 17920 30252
rect 16304 30132 16356 30184
rect 17316 30132 17368 30184
rect 19156 30243 19208 30252
rect 19156 30209 19165 30243
rect 19165 30209 19199 30243
rect 19199 30209 19208 30243
rect 19156 30200 19208 30209
rect 19064 30132 19116 30184
rect 19892 30243 19944 30252
rect 19892 30209 19901 30243
rect 19901 30209 19935 30243
rect 19935 30209 19944 30243
rect 19892 30200 19944 30209
rect 20628 30336 20680 30388
rect 21088 30336 21140 30388
rect 20444 30268 20496 30320
rect 21824 30268 21876 30320
rect 20536 30200 20588 30252
rect 21272 30243 21324 30252
rect 21272 30209 21281 30243
rect 21281 30209 21315 30243
rect 21315 30209 21324 30243
rect 21272 30200 21324 30209
rect 20168 30132 20220 30184
rect 2596 30064 2648 30116
rect 3240 30064 3292 30116
rect 4620 30064 4672 30116
rect 5172 30064 5224 30116
rect 5448 30064 5500 30116
rect 3884 30039 3936 30048
rect 3884 30005 3893 30039
rect 3893 30005 3927 30039
rect 3927 30005 3936 30039
rect 3884 29996 3936 30005
rect 5816 29996 5868 30048
rect 5908 29996 5960 30048
rect 6460 29996 6512 30048
rect 17040 30064 17092 30116
rect 18696 30107 18748 30116
rect 18696 30073 18705 30107
rect 18705 30073 18739 30107
rect 18739 30073 18748 30107
rect 18696 30064 18748 30073
rect 19800 30107 19852 30116
rect 19800 30073 19809 30107
rect 19809 30073 19843 30107
rect 19843 30073 19852 30107
rect 19800 30064 19852 30073
rect 20812 30064 20864 30116
rect 21640 30243 21692 30252
rect 21640 30209 21649 30243
rect 21649 30209 21683 30243
rect 21683 30209 21692 30243
rect 21640 30200 21692 30209
rect 22008 30243 22060 30252
rect 22008 30209 22012 30243
rect 22012 30209 22046 30243
rect 22046 30209 22060 30243
rect 22008 30200 22060 30209
rect 22192 30243 22244 30252
rect 22192 30209 22201 30243
rect 22201 30209 22235 30243
rect 22235 30209 22244 30243
rect 22192 30200 22244 30209
rect 23020 30336 23072 30388
rect 25688 30336 25740 30388
rect 27804 30336 27856 30388
rect 32312 30336 32364 30388
rect 35072 30379 35124 30388
rect 35072 30345 35081 30379
rect 35081 30345 35115 30379
rect 35115 30345 35124 30379
rect 35072 30336 35124 30345
rect 35440 30336 35492 30388
rect 26148 30268 26200 30320
rect 26240 30311 26292 30320
rect 26240 30277 26249 30311
rect 26249 30277 26283 30311
rect 26283 30277 26292 30311
rect 26240 30268 26292 30277
rect 34704 30311 34756 30320
rect 34704 30277 34731 30311
rect 34731 30277 34756 30311
rect 34704 30268 34756 30277
rect 22468 30243 22520 30252
rect 22468 30209 22477 30243
rect 22477 30209 22511 30243
rect 22511 30209 22520 30243
rect 22468 30200 22520 30209
rect 21548 30175 21600 30184
rect 21548 30141 21557 30175
rect 21557 30141 21591 30175
rect 21591 30141 21600 30175
rect 21548 30132 21600 30141
rect 14004 30039 14056 30048
rect 14004 30005 14013 30039
rect 14013 30005 14047 30039
rect 14047 30005 14056 30039
rect 14004 29996 14056 30005
rect 15384 29996 15436 30048
rect 16764 29996 16816 30048
rect 17132 29996 17184 30048
rect 18236 29996 18288 30048
rect 18328 30039 18380 30048
rect 18328 30005 18337 30039
rect 18337 30005 18371 30039
rect 18371 30005 18380 30039
rect 18328 29996 18380 30005
rect 18420 29996 18472 30048
rect 21180 29996 21232 30048
rect 23296 30132 23348 30184
rect 24584 30132 24636 30184
rect 26516 30243 26568 30252
rect 26516 30209 26525 30243
rect 26525 30209 26559 30243
rect 26559 30209 26568 30243
rect 26516 30200 26568 30209
rect 26792 30243 26844 30252
rect 26792 30209 26801 30243
rect 26801 30209 26835 30243
rect 26835 30209 26844 30243
rect 26792 30200 26844 30209
rect 31760 30200 31812 30252
rect 22468 29996 22520 30048
rect 23204 29996 23256 30048
rect 24492 29996 24544 30048
rect 24676 29996 24728 30048
rect 26608 30132 26660 30184
rect 32956 30200 33008 30252
rect 33140 30200 33192 30252
rect 34336 30200 34388 30252
rect 33692 30132 33744 30184
rect 34612 30132 34664 30184
rect 26056 30064 26108 30116
rect 30472 30064 30524 30116
rect 33968 30064 34020 30116
rect 36360 30336 36412 30388
rect 37556 30336 37608 30388
rect 38200 30379 38252 30388
rect 38200 30345 38209 30379
rect 38209 30345 38243 30379
rect 38243 30345 38252 30379
rect 38200 30336 38252 30345
rect 40040 30336 40092 30388
rect 40500 30379 40552 30388
rect 40500 30345 40509 30379
rect 40509 30345 40543 30379
rect 40543 30345 40552 30379
rect 40500 30336 40552 30345
rect 40960 30379 41012 30388
rect 40960 30345 40969 30379
rect 40969 30345 41003 30379
rect 41003 30345 41012 30379
rect 40960 30336 41012 30345
rect 41236 30336 41288 30388
rect 36728 30268 36780 30320
rect 35992 30243 36044 30252
rect 35992 30209 36037 30243
rect 36037 30209 36044 30243
rect 35992 30200 36044 30209
rect 36176 30243 36228 30252
rect 36176 30209 36185 30243
rect 36185 30209 36219 30243
rect 36219 30209 36228 30243
rect 36176 30200 36228 30209
rect 36268 30243 36320 30252
rect 36268 30209 36277 30243
rect 36277 30209 36311 30243
rect 36311 30209 36320 30243
rect 36268 30200 36320 30209
rect 36452 30243 36504 30252
rect 36452 30209 36461 30243
rect 36461 30209 36495 30243
rect 36495 30209 36504 30243
rect 36452 30200 36504 30209
rect 36544 30243 36596 30252
rect 36544 30209 36553 30243
rect 36553 30209 36587 30243
rect 36587 30209 36596 30243
rect 36544 30200 36596 30209
rect 36636 30243 36688 30252
rect 36636 30209 36645 30243
rect 36645 30209 36679 30243
rect 36679 30209 36688 30243
rect 36636 30200 36688 30209
rect 35808 30132 35860 30184
rect 37372 30200 37424 30252
rect 37924 30268 37976 30320
rect 37556 30243 37608 30252
rect 37556 30209 37565 30243
rect 37565 30209 37599 30243
rect 37599 30209 37608 30243
rect 37556 30200 37608 30209
rect 37832 30200 37884 30252
rect 38660 30268 38712 30320
rect 38752 30268 38804 30320
rect 39120 30311 39172 30320
rect 39120 30277 39129 30311
rect 39129 30277 39163 30311
rect 39163 30277 39172 30311
rect 39120 30268 39172 30277
rect 39948 30268 40000 30320
rect 38384 30200 38436 30252
rect 39764 30200 39816 30252
rect 38660 30175 38712 30184
rect 38660 30141 38669 30175
rect 38669 30141 38703 30175
rect 38703 30141 38712 30175
rect 38660 30132 38712 30141
rect 38936 30132 38988 30184
rect 39028 30132 39080 30184
rect 41788 30243 41840 30252
rect 41788 30209 41797 30243
rect 41797 30209 41831 30243
rect 41831 30209 41840 30243
rect 41788 30200 41840 30209
rect 40408 30132 40460 30184
rect 40592 30132 40644 30184
rect 26148 29996 26200 30048
rect 34428 29996 34480 30048
rect 34796 29996 34848 30048
rect 35624 29996 35676 30048
rect 35900 29996 35952 30048
rect 36268 29996 36320 30048
rect 36544 29996 36596 30048
rect 40040 29996 40092 30048
rect 41972 30039 42024 30048
rect 41972 30005 41981 30039
rect 41981 30005 42015 30039
rect 42015 30005 42024 30039
rect 41972 29996 42024 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3424 29724 3476 29776
rect 3608 29724 3660 29776
rect 5632 29792 5684 29844
rect 9036 29792 9088 29844
rect 13084 29835 13136 29844
rect 13084 29801 13093 29835
rect 13093 29801 13127 29835
rect 13127 29801 13136 29835
rect 13084 29792 13136 29801
rect 16304 29835 16356 29844
rect 16304 29801 16313 29835
rect 16313 29801 16347 29835
rect 16347 29801 16356 29835
rect 16304 29792 16356 29801
rect 4436 29656 4488 29708
rect 5724 29724 5776 29776
rect 6092 29724 6144 29776
rect 6552 29724 6604 29776
rect 1768 29588 1820 29640
rect 2872 29588 2924 29640
rect 3056 29631 3108 29640
rect 3056 29597 3065 29631
rect 3065 29597 3099 29631
rect 3099 29597 3108 29631
rect 3056 29588 3108 29597
rect 3700 29588 3752 29640
rect 3792 29588 3844 29640
rect 3976 29631 4028 29640
rect 3976 29597 3985 29631
rect 3985 29597 4019 29631
rect 4019 29597 4028 29631
rect 3976 29588 4028 29597
rect 1952 29520 2004 29572
rect 2412 29495 2464 29504
rect 2412 29461 2421 29495
rect 2421 29461 2455 29495
rect 2455 29461 2464 29495
rect 2412 29452 2464 29461
rect 2872 29495 2924 29504
rect 2872 29461 2881 29495
rect 2881 29461 2915 29495
rect 2915 29461 2924 29495
rect 2872 29452 2924 29461
rect 3148 29563 3200 29572
rect 3148 29529 3157 29563
rect 3157 29529 3191 29563
rect 3191 29529 3200 29563
rect 3148 29520 3200 29529
rect 3884 29520 3936 29572
rect 4344 29588 4396 29640
rect 4804 29520 4856 29572
rect 5448 29588 5500 29640
rect 5632 29631 5684 29640
rect 5632 29597 5641 29631
rect 5641 29597 5675 29631
rect 5675 29597 5684 29631
rect 5632 29588 5684 29597
rect 5908 29699 5960 29708
rect 5908 29665 5917 29699
rect 5917 29665 5951 29699
rect 5951 29665 5960 29699
rect 5908 29656 5960 29665
rect 6460 29656 6512 29708
rect 6644 29699 6696 29708
rect 6644 29665 6653 29699
rect 6653 29665 6687 29699
rect 6687 29665 6696 29699
rect 6644 29656 6696 29665
rect 5816 29588 5868 29640
rect 10968 29724 11020 29776
rect 13544 29724 13596 29776
rect 10232 29656 10284 29708
rect 11612 29656 11664 29708
rect 14004 29656 14056 29708
rect 3608 29452 3660 29504
rect 3792 29495 3844 29504
rect 3792 29461 3801 29495
rect 3801 29461 3835 29495
rect 3835 29461 3844 29495
rect 3792 29452 3844 29461
rect 3976 29452 4028 29504
rect 5724 29452 5776 29504
rect 8208 29452 8260 29504
rect 13268 29631 13320 29640
rect 13268 29597 13277 29631
rect 13277 29597 13311 29631
rect 13311 29597 13320 29631
rect 13268 29588 13320 29597
rect 15200 29631 15252 29640
rect 15200 29597 15209 29631
rect 15209 29597 15243 29631
rect 15243 29597 15252 29631
rect 15200 29588 15252 29597
rect 17592 29792 17644 29844
rect 19156 29792 19208 29844
rect 19708 29835 19760 29844
rect 19708 29801 19717 29835
rect 19717 29801 19751 29835
rect 19751 29801 19760 29835
rect 19708 29792 19760 29801
rect 21180 29835 21232 29844
rect 21180 29801 21210 29835
rect 21210 29801 21232 29835
rect 18328 29724 18380 29776
rect 21180 29792 21232 29801
rect 21824 29792 21876 29844
rect 22468 29792 22520 29844
rect 16764 29699 16816 29708
rect 16764 29665 16773 29699
rect 16773 29665 16807 29699
rect 16807 29665 16816 29699
rect 16764 29656 16816 29665
rect 16856 29656 16908 29708
rect 18236 29656 18288 29708
rect 10416 29520 10468 29572
rect 11796 29520 11848 29572
rect 12992 29520 13044 29572
rect 13544 29452 13596 29504
rect 13912 29520 13964 29572
rect 16948 29631 17000 29640
rect 16948 29597 16957 29631
rect 16957 29597 16991 29631
rect 16991 29597 17000 29631
rect 16948 29588 17000 29597
rect 17408 29588 17460 29640
rect 17868 29588 17920 29640
rect 17960 29520 18012 29572
rect 14740 29452 14792 29504
rect 16212 29452 16264 29504
rect 17224 29452 17276 29504
rect 17592 29452 17644 29504
rect 17776 29495 17828 29504
rect 17776 29461 17785 29495
rect 17785 29461 17819 29495
rect 17819 29461 17828 29495
rect 17776 29452 17828 29461
rect 18420 29588 18472 29640
rect 18604 29588 18656 29640
rect 19800 29656 19852 29708
rect 23848 29724 23900 29776
rect 24584 29792 24636 29844
rect 25228 29724 25280 29776
rect 26516 29792 26568 29844
rect 26608 29792 26660 29844
rect 32588 29792 32640 29844
rect 32956 29835 33008 29844
rect 32956 29801 32965 29835
rect 32965 29801 32999 29835
rect 32999 29801 33008 29835
rect 32956 29792 33008 29801
rect 19524 29588 19576 29640
rect 20076 29588 20128 29640
rect 18696 29563 18748 29572
rect 18696 29529 18705 29563
rect 18705 29529 18739 29563
rect 18739 29529 18748 29563
rect 18696 29520 18748 29529
rect 20260 29631 20312 29640
rect 20260 29597 20269 29631
rect 20269 29597 20303 29631
rect 20303 29597 20312 29631
rect 20260 29588 20312 29597
rect 20720 29588 20772 29640
rect 23020 29588 23072 29640
rect 23204 29588 23256 29640
rect 23480 29631 23532 29640
rect 23480 29597 23487 29631
rect 23487 29597 23532 29631
rect 23480 29588 23532 29597
rect 23664 29631 23716 29640
rect 23664 29597 23673 29631
rect 23673 29597 23707 29631
rect 23707 29597 23716 29631
rect 23664 29588 23716 29597
rect 23756 29631 23808 29640
rect 23756 29597 23770 29631
rect 23770 29597 23804 29631
rect 23804 29597 23808 29631
rect 23756 29588 23808 29597
rect 19616 29452 19668 29504
rect 21364 29452 21416 29504
rect 24492 29699 24544 29708
rect 24492 29665 24501 29699
rect 24501 29665 24535 29699
rect 24535 29665 24544 29699
rect 24492 29656 24544 29665
rect 24584 29656 24636 29708
rect 31484 29724 31536 29776
rect 31668 29724 31720 29776
rect 31760 29724 31812 29776
rect 33140 29792 33192 29844
rect 33692 29835 33744 29844
rect 33692 29801 33701 29835
rect 33701 29801 33735 29835
rect 33735 29801 33744 29835
rect 33692 29792 33744 29801
rect 34152 29792 34204 29844
rect 34612 29792 34664 29844
rect 26608 29699 26660 29708
rect 26608 29665 26617 29699
rect 26617 29665 26651 29699
rect 26651 29665 26660 29699
rect 26608 29656 26660 29665
rect 24124 29588 24176 29640
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 24768 29588 24820 29597
rect 25596 29631 25648 29640
rect 25596 29597 25605 29631
rect 25605 29597 25639 29631
rect 25639 29597 25648 29631
rect 25596 29588 25648 29597
rect 25780 29588 25832 29640
rect 26516 29588 26568 29640
rect 26792 29588 26844 29640
rect 27896 29656 27948 29708
rect 30472 29699 30524 29708
rect 30472 29665 30481 29699
rect 30481 29665 30515 29699
rect 30515 29665 30524 29699
rect 30472 29656 30524 29665
rect 34244 29767 34296 29776
rect 34244 29733 34253 29767
rect 34253 29733 34287 29767
rect 34287 29733 34296 29767
rect 34244 29724 34296 29733
rect 32772 29699 32824 29708
rect 32772 29665 32781 29699
rect 32781 29665 32815 29699
rect 32815 29665 32824 29699
rect 32772 29656 32824 29665
rect 21824 29452 21876 29504
rect 22100 29452 22152 29504
rect 25320 29520 25372 29572
rect 27344 29631 27396 29640
rect 27344 29597 27353 29631
rect 27353 29597 27387 29631
rect 27387 29597 27396 29631
rect 27344 29588 27396 29597
rect 27436 29631 27488 29640
rect 27436 29597 27445 29631
rect 27445 29597 27479 29631
rect 27479 29597 27488 29631
rect 27436 29588 27488 29597
rect 27620 29631 27672 29640
rect 27620 29597 27629 29631
rect 27629 29597 27663 29631
rect 27663 29597 27672 29631
rect 27620 29588 27672 29597
rect 28540 29588 28592 29640
rect 29736 29631 29788 29640
rect 29736 29597 29745 29631
rect 29745 29597 29779 29631
rect 29779 29597 29788 29631
rect 29736 29588 29788 29597
rect 29828 29631 29880 29640
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 30104 29631 30156 29640
rect 30104 29597 30113 29631
rect 30113 29597 30147 29631
rect 30147 29597 30156 29631
rect 30104 29588 30156 29597
rect 30380 29588 30432 29640
rect 31024 29588 31076 29640
rect 31116 29631 31168 29640
rect 31116 29597 31125 29631
rect 31125 29597 31159 29631
rect 31159 29597 31168 29631
rect 31116 29588 31168 29597
rect 27252 29520 27304 29572
rect 25504 29452 25556 29504
rect 25872 29495 25924 29504
rect 25872 29461 25881 29495
rect 25881 29461 25915 29495
rect 25915 29461 25924 29495
rect 25872 29452 25924 29461
rect 26516 29452 26568 29504
rect 29000 29520 29052 29572
rect 34428 29656 34480 29708
rect 34980 29699 35032 29708
rect 34980 29665 34989 29699
rect 34989 29665 35023 29699
rect 35023 29665 35032 29699
rect 34980 29656 35032 29665
rect 33048 29520 33100 29572
rect 30564 29452 30616 29504
rect 31300 29452 31352 29504
rect 32404 29452 32456 29504
rect 32864 29452 32916 29504
rect 33416 29631 33468 29640
rect 33416 29597 33461 29631
rect 33461 29597 33468 29631
rect 33416 29588 33468 29597
rect 33600 29631 33652 29640
rect 33600 29597 33609 29631
rect 33609 29597 33643 29631
rect 33643 29597 33652 29631
rect 33600 29588 33652 29597
rect 35992 29792 36044 29844
rect 36084 29792 36136 29844
rect 35532 29724 35584 29776
rect 33876 29563 33928 29572
rect 33876 29529 33885 29563
rect 33885 29529 33919 29563
rect 33919 29529 33928 29563
rect 33876 29520 33928 29529
rect 34060 29520 34112 29572
rect 35440 29631 35492 29640
rect 35440 29597 35449 29631
rect 35449 29597 35483 29631
rect 35483 29597 35492 29631
rect 35440 29588 35492 29597
rect 35624 29588 35676 29640
rect 34796 29520 34848 29572
rect 33416 29452 33468 29504
rect 35900 29588 35952 29640
rect 36360 29588 36412 29640
rect 36820 29656 36872 29708
rect 36728 29631 36780 29640
rect 36728 29597 36738 29631
rect 36738 29597 36772 29631
rect 36772 29597 36780 29631
rect 38660 29792 38712 29844
rect 40684 29792 40736 29844
rect 42156 29835 42208 29844
rect 42156 29801 42165 29835
rect 42165 29801 42199 29835
rect 42199 29801 42208 29835
rect 42156 29792 42208 29801
rect 40132 29724 40184 29776
rect 38016 29656 38068 29708
rect 38476 29656 38528 29708
rect 39488 29699 39540 29708
rect 39488 29665 39497 29699
rect 39497 29665 39531 29699
rect 39531 29665 39540 29699
rect 39488 29656 39540 29665
rect 40316 29656 40368 29708
rect 36728 29588 36780 29597
rect 37096 29588 37148 29640
rect 37832 29588 37884 29640
rect 39856 29631 39908 29640
rect 39856 29597 39865 29631
rect 39865 29597 39899 29631
rect 39899 29597 39908 29631
rect 39856 29588 39908 29597
rect 40040 29588 40092 29640
rect 40408 29631 40460 29640
rect 40408 29597 40417 29631
rect 40417 29597 40451 29631
rect 40451 29597 40460 29631
rect 40408 29588 40460 29597
rect 35532 29452 35584 29504
rect 35716 29452 35768 29504
rect 36176 29452 36228 29504
rect 37372 29520 37424 29572
rect 40776 29520 40828 29572
rect 41696 29520 41748 29572
rect 38568 29452 38620 29504
rect 40500 29452 40552 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 1952 29155 2004 29164
rect 1952 29121 1961 29155
rect 1961 29121 1995 29155
rect 1995 29121 2004 29155
rect 1952 29112 2004 29121
rect 3792 29248 3844 29300
rect 4712 29248 4764 29300
rect 5540 29291 5592 29300
rect 5540 29257 5549 29291
rect 5549 29257 5583 29291
rect 5583 29257 5592 29291
rect 5540 29248 5592 29257
rect 5724 29248 5776 29300
rect 2412 29223 2464 29232
rect 2412 29189 2421 29223
rect 2421 29189 2455 29223
rect 2455 29189 2464 29223
rect 2412 29180 2464 29189
rect 3056 29180 3108 29232
rect 3148 29180 3200 29232
rect 4436 29223 4488 29232
rect 4436 29189 4445 29223
rect 4445 29189 4479 29223
rect 4479 29189 4488 29223
rect 4436 29180 4488 29189
rect 3608 29112 3660 29164
rect 4160 29155 4212 29164
rect 4160 29121 4169 29155
rect 4169 29121 4203 29155
rect 4203 29121 4212 29155
rect 4160 29112 4212 29121
rect 4712 29044 4764 29096
rect 3424 28976 3476 29028
rect 3976 28976 4028 29028
rect 5172 29155 5224 29164
rect 5172 29121 5181 29155
rect 5181 29121 5215 29155
rect 5215 29121 5224 29155
rect 5172 29112 5224 29121
rect 5172 28976 5224 29028
rect 5724 29155 5776 29164
rect 5724 29121 5733 29155
rect 5733 29121 5767 29155
rect 5767 29121 5776 29155
rect 5724 29112 5776 29121
rect 5816 29155 5868 29164
rect 5816 29121 5825 29155
rect 5825 29121 5859 29155
rect 5859 29121 5868 29155
rect 5816 29112 5868 29121
rect 6460 29248 6512 29300
rect 11796 29248 11848 29300
rect 13360 29248 13412 29300
rect 16488 29248 16540 29300
rect 17408 29291 17460 29300
rect 17408 29257 17417 29291
rect 17417 29257 17451 29291
rect 17451 29257 17460 29291
rect 17408 29248 17460 29257
rect 17592 29248 17644 29300
rect 18236 29248 18288 29300
rect 18972 29248 19024 29300
rect 19249 29248 19301 29300
rect 21364 29248 21416 29300
rect 24768 29248 24820 29300
rect 25228 29248 25280 29300
rect 6276 29112 6328 29164
rect 8208 29112 8260 29164
rect 17132 29180 17184 29232
rect 6552 29044 6604 29096
rect 9496 29087 9548 29096
rect 9496 29053 9505 29087
rect 9505 29053 9539 29087
rect 9539 29053 9548 29087
rect 9496 29044 9548 29053
rect 9772 29087 9824 29096
rect 9772 29053 9781 29087
rect 9781 29053 9815 29087
rect 9815 29053 9824 29087
rect 9772 29044 9824 29053
rect 10968 29044 11020 29096
rect 5724 28976 5776 29028
rect 13452 29155 13504 29164
rect 13452 29121 13461 29155
rect 13461 29121 13495 29155
rect 13495 29121 13504 29155
rect 13452 29112 13504 29121
rect 13544 29155 13596 29164
rect 13544 29121 13553 29155
rect 13553 29121 13587 29155
rect 13587 29121 13596 29155
rect 13544 29112 13596 29121
rect 11244 29019 11296 29028
rect 11244 28985 11253 29019
rect 11253 28985 11287 29019
rect 11287 28985 11296 29019
rect 11244 28976 11296 28985
rect 12532 29044 12584 29096
rect 13268 29044 13320 29096
rect 17040 29112 17092 29164
rect 17776 29180 17828 29232
rect 16856 29044 16908 29096
rect 17132 29044 17184 29096
rect 13544 28976 13596 29028
rect 17316 28976 17368 29028
rect 17684 28976 17736 29028
rect 17960 29112 18012 29164
rect 18696 29180 18748 29232
rect 17868 29087 17920 29096
rect 17868 29053 17877 29087
rect 17877 29053 17911 29087
rect 17911 29053 17920 29087
rect 17868 29044 17920 29053
rect 19432 29112 19484 29164
rect 19616 29155 19668 29164
rect 19616 29121 19625 29155
rect 19625 29121 19659 29155
rect 19659 29121 19668 29155
rect 19616 29112 19668 29121
rect 19800 29155 19852 29164
rect 19800 29121 19809 29155
rect 19809 29121 19843 29155
rect 19843 29121 19852 29155
rect 19800 29112 19852 29121
rect 20996 29112 21048 29164
rect 21824 29155 21876 29164
rect 18696 28976 18748 29028
rect 19064 29044 19116 29096
rect 19524 29087 19576 29096
rect 19524 29053 19533 29087
rect 19533 29053 19567 29087
rect 19567 29053 19576 29087
rect 19524 29044 19576 29053
rect 20260 29044 20312 29096
rect 21824 29121 21833 29155
rect 21833 29121 21867 29155
rect 21867 29121 21876 29155
rect 21824 29112 21876 29121
rect 22008 29155 22060 29164
rect 22008 29121 22030 29155
rect 22030 29121 22060 29155
rect 22008 29112 22060 29121
rect 22100 29155 22152 29164
rect 22100 29121 22109 29155
rect 22109 29121 22143 29155
rect 22143 29121 22152 29155
rect 22100 29112 22152 29121
rect 22468 29180 22520 29232
rect 22744 29180 22796 29232
rect 23388 29180 23440 29232
rect 23572 29180 23624 29232
rect 24400 29180 24452 29232
rect 25872 29180 25924 29232
rect 19616 28976 19668 29028
rect 2044 28951 2096 28960
rect 2044 28917 2053 28951
rect 2053 28917 2087 28951
rect 2087 28917 2096 28951
rect 2044 28908 2096 28917
rect 4344 28908 4396 28960
rect 5080 28908 5132 28960
rect 5632 28908 5684 28960
rect 12900 28908 12952 28960
rect 12992 28908 13044 28960
rect 17776 28908 17828 28960
rect 18328 28908 18380 28960
rect 21456 28908 21508 28960
rect 22376 28908 22428 28960
rect 22560 29044 22612 29096
rect 23112 29155 23164 29164
rect 23112 29121 23121 29155
rect 23121 29121 23155 29155
rect 23155 29121 23164 29155
rect 23112 29112 23164 29121
rect 23020 29044 23072 29096
rect 23296 29112 23348 29164
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 24308 29155 24360 29164
rect 24308 29121 24317 29155
rect 24317 29121 24351 29155
rect 24351 29121 24360 29155
rect 24308 29112 24360 29121
rect 25228 29155 25280 29164
rect 25228 29121 25237 29155
rect 25237 29121 25271 29155
rect 25271 29121 25280 29155
rect 25228 29112 25280 29121
rect 25780 29112 25832 29164
rect 26608 29223 26660 29232
rect 26608 29189 26617 29223
rect 26617 29189 26651 29223
rect 26651 29189 26660 29223
rect 26608 29180 26660 29189
rect 26792 29248 26844 29300
rect 27436 29248 27488 29300
rect 27160 29180 27212 29232
rect 27804 29223 27856 29232
rect 27804 29189 27813 29223
rect 27813 29189 27847 29223
rect 27847 29189 27856 29223
rect 27804 29180 27856 29189
rect 27896 29223 27948 29232
rect 27896 29189 27905 29223
rect 27905 29189 27939 29223
rect 27939 29189 27948 29223
rect 27896 29180 27948 29189
rect 25596 29044 25648 29096
rect 27344 29112 27396 29164
rect 28080 29112 28132 29164
rect 29184 29248 29236 29300
rect 31024 29248 31076 29300
rect 32036 29248 32088 29300
rect 28540 29223 28592 29232
rect 28540 29189 28549 29223
rect 28549 29189 28583 29223
rect 28583 29189 28592 29223
rect 28540 29180 28592 29189
rect 28632 29180 28684 29232
rect 26608 29044 26660 29096
rect 26792 29044 26844 29096
rect 30104 29155 30156 29164
rect 30104 29121 30113 29155
rect 30113 29121 30147 29155
rect 30147 29121 30156 29155
rect 30104 29112 30156 29121
rect 30380 29180 30432 29232
rect 30656 29180 30708 29232
rect 32864 29248 32916 29300
rect 33048 29291 33100 29300
rect 33048 29257 33057 29291
rect 33057 29257 33091 29291
rect 33091 29257 33100 29291
rect 33048 29248 33100 29257
rect 33232 29248 33284 29300
rect 36360 29248 36412 29300
rect 36912 29248 36964 29300
rect 30564 29155 30616 29164
rect 30564 29121 30573 29155
rect 30573 29121 30607 29155
rect 30607 29121 30616 29155
rect 30564 29112 30616 29121
rect 31024 29155 31076 29164
rect 31024 29121 31033 29155
rect 31033 29121 31067 29155
rect 31067 29121 31076 29155
rect 31024 29112 31076 29121
rect 31116 29155 31168 29164
rect 31116 29121 31125 29155
rect 31125 29121 31159 29155
rect 31159 29121 31168 29155
rect 31116 29112 31168 29121
rect 31300 29112 31352 29164
rect 32220 29155 32272 29164
rect 32220 29121 32230 29155
rect 32230 29121 32264 29155
rect 32264 29121 32272 29155
rect 32220 29112 32272 29121
rect 23664 28976 23716 29028
rect 24584 28976 24636 29028
rect 31484 29087 31536 29096
rect 31484 29053 31493 29087
rect 31493 29053 31527 29087
rect 31527 29053 31536 29087
rect 31484 29044 31536 29053
rect 33048 29112 33100 29164
rect 33140 29112 33192 29164
rect 34060 29180 34112 29232
rect 34336 29180 34388 29232
rect 28172 29019 28224 29028
rect 28172 28985 28181 29019
rect 28181 28985 28215 29019
rect 28215 28985 28224 29019
rect 28172 28976 28224 28985
rect 29736 28976 29788 29028
rect 23296 28908 23348 28960
rect 25044 28951 25096 28960
rect 25044 28917 25053 28951
rect 25053 28917 25087 28951
rect 25087 28917 25096 28951
rect 25044 28908 25096 28917
rect 26424 28951 26476 28960
rect 26424 28917 26433 28951
rect 26433 28917 26467 28951
rect 26467 28917 26476 28951
rect 26424 28908 26476 28917
rect 27068 28908 27120 28960
rect 30380 28908 30432 28960
rect 33416 29044 33468 29096
rect 33600 28976 33652 29028
rect 33876 29155 33928 29164
rect 33876 29121 33885 29155
rect 33885 29121 33919 29155
rect 33919 29121 33928 29155
rect 33876 29112 33928 29121
rect 34888 29112 34940 29164
rect 34428 29044 34480 29096
rect 35532 29112 35584 29164
rect 35900 29112 35952 29164
rect 36820 29180 36872 29232
rect 36176 29155 36228 29164
rect 36176 29121 36185 29155
rect 36185 29121 36219 29155
rect 36219 29121 36228 29155
rect 36176 29112 36228 29121
rect 39948 29180 40000 29232
rect 35624 29044 35676 29096
rect 41880 29155 41932 29164
rect 36452 29044 36504 29096
rect 36820 29044 36872 29096
rect 37924 29044 37976 29096
rect 41880 29121 41889 29155
rect 41889 29121 41923 29155
rect 41923 29121 41932 29155
rect 41880 29112 41932 29121
rect 40132 29044 40184 29096
rect 40408 29044 40460 29096
rect 34152 29019 34204 29028
rect 34152 28985 34161 29019
rect 34161 28985 34195 29019
rect 34195 28985 34204 29019
rect 34152 28976 34204 28985
rect 34244 29019 34296 29028
rect 34244 28985 34253 29019
rect 34253 28985 34287 29019
rect 34287 28985 34296 29019
rect 34244 28976 34296 28985
rect 35256 28976 35308 29028
rect 35808 28976 35860 29028
rect 35992 28976 36044 29028
rect 36912 28976 36964 29028
rect 39028 29019 39080 29028
rect 39028 28985 39037 29019
rect 39037 28985 39071 29019
rect 39071 28985 39080 29019
rect 39028 28976 39080 28985
rect 39856 28976 39908 29028
rect 34796 28908 34848 28960
rect 40684 28976 40736 29028
rect 42064 29019 42116 29028
rect 42064 28985 42073 29019
rect 42073 28985 42107 29019
rect 42107 28985 42116 29019
rect 42064 28976 42116 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 3608 28704 3660 28756
rect 4804 28704 4856 28756
rect 3056 28636 3108 28688
rect 3700 28636 3752 28688
rect 5356 28704 5408 28756
rect 6000 28704 6052 28756
rect 6828 28704 6880 28756
rect 7472 28704 7524 28756
rect 10876 28704 10928 28756
rect 13544 28704 13596 28756
rect 13912 28747 13964 28756
rect 13912 28713 13921 28747
rect 13921 28713 13955 28747
rect 13955 28713 13964 28747
rect 13912 28704 13964 28713
rect 17960 28704 18012 28756
rect 18604 28704 18656 28756
rect 19248 28747 19300 28756
rect 19248 28713 19257 28747
rect 19257 28713 19291 28747
rect 19291 28713 19300 28747
rect 19248 28704 19300 28713
rect 21272 28747 21324 28756
rect 21272 28713 21281 28747
rect 21281 28713 21315 28747
rect 21315 28713 21324 28747
rect 21272 28704 21324 28713
rect 21364 28704 21416 28756
rect 21824 28704 21876 28756
rect 22560 28747 22612 28756
rect 22560 28713 22569 28747
rect 22569 28713 22603 28747
rect 22603 28713 22612 28747
rect 22560 28704 22612 28713
rect 23112 28704 23164 28756
rect 23664 28747 23716 28756
rect 23664 28713 23673 28747
rect 23673 28713 23707 28747
rect 23707 28713 23716 28747
rect 23664 28704 23716 28713
rect 25780 28704 25832 28756
rect 26148 28704 26200 28756
rect 29276 28704 29328 28756
rect 29828 28704 29880 28756
rect 30656 28747 30708 28756
rect 30656 28713 30665 28747
rect 30665 28713 30699 28747
rect 30699 28713 30708 28747
rect 30656 28704 30708 28713
rect 30748 28704 30800 28756
rect 31024 28747 31076 28756
rect 31024 28713 31033 28747
rect 31033 28713 31067 28747
rect 31067 28713 31076 28747
rect 31024 28704 31076 28713
rect 34336 28704 34388 28756
rect 34796 28704 34848 28756
rect 36176 28704 36228 28756
rect 41880 28704 41932 28756
rect 1400 28611 1452 28620
rect 1400 28577 1409 28611
rect 1409 28577 1443 28611
rect 1443 28577 1452 28611
rect 1400 28568 1452 28577
rect 2044 28568 2096 28620
rect 3424 28568 3476 28620
rect 2780 28500 2832 28552
rect 4160 28543 4212 28552
rect 4160 28509 4169 28543
rect 4169 28509 4203 28543
rect 4203 28509 4212 28543
rect 4160 28500 4212 28509
rect 5080 28636 5132 28688
rect 5540 28636 5592 28688
rect 11980 28636 12032 28688
rect 4804 28568 4856 28620
rect 4620 28500 4672 28552
rect 3608 28364 3660 28416
rect 4804 28432 4856 28484
rect 5172 28543 5224 28552
rect 5172 28509 5181 28543
rect 5181 28509 5215 28543
rect 5215 28509 5224 28543
rect 5172 28500 5224 28509
rect 5540 28500 5592 28552
rect 9496 28568 9548 28620
rect 12716 28679 12768 28688
rect 12716 28645 12725 28679
rect 12725 28645 12759 28679
rect 12759 28645 12768 28679
rect 12716 28636 12768 28645
rect 14648 28636 14700 28688
rect 6276 28543 6328 28552
rect 6276 28509 6285 28543
rect 6285 28509 6319 28543
rect 6319 28509 6328 28543
rect 6276 28500 6328 28509
rect 7656 28543 7708 28552
rect 7656 28509 7665 28543
rect 7665 28509 7699 28543
rect 7699 28509 7708 28543
rect 7656 28500 7708 28509
rect 11520 28543 11572 28552
rect 11520 28509 11529 28543
rect 11529 28509 11563 28543
rect 11563 28509 11572 28543
rect 11520 28500 11572 28509
rect 12808 28500 12860 28552
rect 4620 28364 4672 28416
rect 5356 28432 5408 28484
rect 10968 28432 11020 28484
rect 11612 28432 11664 28484
rect 12348 28475 12400 28484
rect 12348 28441 12357 28475
rect 12357 28441 12391 28475
rect 12391 28441 12400 28475
rect 12348 28432 12400 28441
rect 12900 28475 12952 28484
rect 12900 28441 12909 28475
rect 12909 28441 12943 28475
rect 12943 28441 12952 28475
rect 12900 28432 12952 28441
rect 11520 28364 11572 28416
rect 12624 28364 12676 28416
rect 14556 28543 14608 28552
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 14924 28611 14976 28620
rect 14924 28577 14933 28611
rect 14933 28577 14967 28611
rect 14967 28577 14976 28611
rect 14924 28568 14976 28577
rect 18236 28636 18288 28688
rect 18788 28636 18840 28688
rect 15568 28568 15620 28620
rect 16672 28568 16724 28620
rect 18512 28568 18564 28620
rect 17132 28500 17184 28552
rect 17408 28500 17460 28552
rect 18144 28500 18196 28552
rect 18236 28543 18288 28552
rect 18236 28509 18245 28543
rect 18245 28509 18279 28543
rect 18279 28509 18288 28543
rect 18236 28500 18288 28509
rect 18972 28500 19024 28552
rect 19064 28543 19116 28552
rect 19064 28509 19073 28543
rect 19073 28509 19107 28543
rect 19107 28509 19116 28543
rect 19064 28500 19116 28509
rect 14464 28407 14516 28416
rect 14464 28373 14473 28407
rect 14473 28373 14507 28407
rect 14507 28373 14516 28407
rect 14464 28364 14516 28373
rect 14832 28364 14884 28416
rect 15200 28475 15252 28484
rect 15200 28441 15209 28475
rect 15209 28441 15243 28475
rect 15243 28441 15252 28475
rect 15200 28432 15252 28441
rect 16856 28432 16908 28484
rect 18052 28432 18104 28484
rect 20168 28636 20220 28688
rect 22008 28636 22060 28688
rect 19432 28543 19484 28552
rect 19432 28509 19441 28543
rect 19441 28509 19475 28543
rect 19475 28509 19484 28543
rect 19432 28500 19484 28509
rect 20812 28500 20864 28552
rect 22192 28568 22244 28620
rect 19616 28475 19668 28484
rect 19616 28441 19625 28475
rect 19625 28441 19659 28475
rect 19659 28441 19668 28475
rect 19616 28432 19668 28441
rect 22376 28500 22428 28552
rect 23480 28636 23532 28688
rect 24308 28636 24360 28688
rect 24400 28636 24452 28688
rect 26056 28636 26108 28688
rect 26424 28636 26476 28688
rect 24124 28568 24176 28620
rect 26884 28568 26936 28620
rect 30564 28636 30616 28688
rect 31208 28679 31260 28688
rect 31208 28645 31217 28679
rect 31217 28645 31251 28679
rect 31251 28645 31260 28679
rect 31208 28636 31260 28645
rect 32036 28636 32088 28688
rect 34704 28636 34756 28688
rect 35532 28636 35584 28688
rect 28724 28568 28776 28620
rect 21456 28475 21508 28484
rect 21456 28441 21465 28475
rect 21465 28441 21499 28475
rect 21499 28441 21508 28475
rect 21456 28432 21508 28441
rect 21548 28432 21600 28484
rect 22192 28432 22244 28484
rect 23020 28543 23072 28552
rect 23020 28509 23029 28543
rect 23029 28509 23063 28543
rect 23063 28509 23072 28543
rect 23020 28500 23072 28509
rect 23112 28500 23164 28552
rect 23296 28543 23348 28552
rect 23296 28509 23305 28543
rect 23305 28509 23339 28543
rect 23339 28509 23348 28543
rect 23296 28500 23348 28509
rect 23388 28543 23440 28552
rect 23388 28509 23397 28543
rect 23397 28509 23431 28543
rect 23431 28509 23440 28543
rect 23388 28500 23440 28509
rect 30104 28568 30156 28620
rect 30748 28611 30800 28620
rect 25688 28500 25740 28552
rect 25964 28500 26016 28552
rect 26516 28543 26568 28552
rect 26516 28509 26525 28543
rect 26525 28509 26559 28543
rect 26559 28509 26568 28543
rect 26516 28500 26568 28509
rect 27068 28543 27120 28552
rect 27068 28509 27077 28543
rect 27077 28509 27111 28543
rect 27111 28509 27120 28543
rect 27068 28500 27120 28509
rect 24308 28432 24360 28484
rect 26332 28432 26384 28484
rect 27620 28500 27672 28552
rect 27712 28500 27764 28552
rect 26056 28407 26108 28416
rect 26056 28373 26065 28407
rect 26065 28373 26099 28407
rect 26099 28373 26108 28407
rect 26056 28364 26108 28373
rect 26516 28364 26568 28416
rect 27528 28432 27580 28484
rect 26792 28364 26844 28416
rect 28816 28364 28868 28416
rect 29644 28543 29696 28552
rect 29644 28509 29654 28543
rect 29654 28509 29688 28543
rect 29688 28509 29696 28543
rect 29644 28500 29696 28509
rect 29920 28543 29972 28552
rect 29920 28509 29929 28543
rect 29929 28509 29963 28543
rect 29963 28509 29972 28543
rect 29920 28500 29972 28509
rect 30012 28543 30064 28552
rect 30012 28509 30026 28543
rect 30026 28509 30060 28543
rect 30060 28509 30064 28543
rect 30012 28500 30064 28509
rect 30288 28543 30340 28552
rect 30288 28509 30297 28543
rect 30297 28509 30331 28543
rect 30331 28509 30340 28543
rect 30288 28500 30340 28509
rect 30472 28543 30524 28552
rect 30472 28509 30481 28543
rect 30481 28509 30515 28543
rect 30515 28509 30524 28543
rect 30472 28500 30524 28509
rect 30748 28577 30763 28611
rect 30763 28577 30797 28611
rect 30797 28577 30800 28611
rect 30748 28568 30800 28577
rect 31116 28568 31168 28620
rect 34060 28611 34112 28620
rect 34060 28577 34069 28611
rect 34069 28577 34103 28611
rect 34103 28577 34112 28611
rect 34060 28568 34112 28577
rect 30656 28432 30708 28484
rect 30932 28432 30984 28484
rect 31852 28543 31904 28552
rect 31852 28509 31861 28543
rect 31861 28509 31895 28543
rect 31895 28509 31904 28543
rect 31852 28500 31904 28509
rect 32036 28543 32088 28552
rect 32036 28509 32045 28543
rect 32045 28509 32079 28543
rect 32079 28509 32088 28543
rect 32036 28500 32088 28509
rect 34428 28568 34480 28620
rect 34152 28432 34204 28484
rect 34612 28432 34664 28484
rect 35716 28543 35768 28552
rect 35716 28509 35725 28543
rect 35725 28509 35759 28543
rect 35759 28509 35768 28543
rect 35716 28500 35768 28509
rect 37924 28611 37976 28620
rect 37924 28577 37933 28611
rect 37933 28577 37967 28611
rect 37967 28577 37976 28611
rect 37924 28568 37976 28577
rect 40684 28611 40736 28620
rect 40684 28577 40693 28611
rect 40693 28577 40727 28611
rect 40727 28577 40736 28611
rect 40684 28568 40736 28577
rect 35900 28543 35952 28552
rect 35900 28509 35909 28543
rect 35909 28509 35943 28543
rect 35943 28509 35952 28543
rect 35900 28500 35952 28509
rect 36544 28500 36596 28552
rect 37648 28543 37700 28552
rect 37648 28509 37657 28543
rect 37657 28509 37691 28543
rect 37691 28509 37700 28543
rect 37648 28500 37700 28509
rect 40132 28500 40184 28552
rect 37832 28475 37884 28484
rect 37832 28441 37841 28475
rect 37841 28441 37875 28475
rect 37875 28441 37884 28475
rect 37832 28432 37884 28441
rect 30564 28364 30616 28416
rect 32312 28364 32364 28416
rect 35348 28407 35400 28416
rect 35348 28373 35357 28407
rect 35357 28373 35391 28407
rect 35391 28373 35400 28407
rect 35348 28364 35400 28373
rect 39948 28432 40000 28484
rect 41696 28432 41748 28484
rect 38844 28364 38896 28416
rect 41512 28364 41564 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 3608 28160 3660 28212
rect 4160 28160 4212 28212
rect 4804 28160 4856 28212
rect 5080 28160 5132 28212
rect 5356 28160 5408 28212
rect 2780 28092 2832 28144
rect 3516 28092 3568 28144
rect 5632 28160 5684 28212
rect 9772 28160 9824 28212
rect 10876 28203 10928 28212
rect 10876 28169 10885 28203
rect 10885 28169 10919 28203
rect 10919 28169 10928 28203
rect 10876 28160 10928 28169
rect 11244 28160 11296 28212
rect 11520 28203 11572 28212
rect 11520 28169 11529 28203
rect 11529 28169 11563 28203
rect 11563 28169 11572 28203
rect 11520 28160 11572 28169
rect 11980 28203 12032 28212
rect 11980 28169 11989 28203
rect 11989 28169 12023 28203
rect 12023 28169 12032 28203
rect 11980 28160 12032 28169
rect 13728 28160 13780 28212
rect 4804 28024 4856 28076
rect 5724 28092 5776 28144
rect 6092 28092 6144 28144
rect 6552 28024 6604 28076
rect 8300 28024 8352 28076
rect 9496 28092 9548 28144
rect 9680 28024 9732 28076
rect 1400 27956 1452 28008
rect 2872 27956 2924 28008
rect 4712 27956 4764 28008
rect 12532 28135 12584 28144
rect 12532 28101 12541 28135
rect 12541 28101 12575 28135
rect 12575 28101 12584 28135
rect 12532 28092 12584 28101
rect 14740 28160 14792 28212
rect 14464 28092 14516 28144
rect 15200 28160 15252 28212
rect 17960 28160 18012 28212
rect 18328 28160 18380 28212
rect 19524 28160 19576 28212
rect 23664 28160 23716 28212
rect 28448 28160 28500 28212
rect 11152 28024 11204 28076
rect 12440 28067 12492 28076
rect 12440 28033 12449 28067
rect 12449 28033 12483 28067
rect 12483 28033 12492 28067
rect 12440 28024 12492 28033
rect 12624 28067 12676 28076
rect 12624 28033 12633 28067
rect 12633 28033 12667 28067
rect 12667 28033 12676 28067
rect 12624 28024 12676 28033
rect 5172 27888 5224 27940
rect 5540 27888 5592 27940
rect 12072 27999 12124 28008
rect 12072 27965 12081 27999
rect 12081 27965 12115 27999
rect 12115 27965 12124 27999
rect 12072 27956 12124 27965
rect 12348 27956 12400 28008
rect 848 27820 900 27872
rect 4988 27863 5040 27872
rect 4988 27829 4997 27863
rect 4997 27829 5031 27863
rect 5031 27829 5040 27863
rect 4988 27820 5040 27829
rect 5080 27820 5132 27872
rect 5816 27820 5868 27872
rect 6184 27820 6236 27872
rect 7656 27820 7708 27872
rect 9036 27863 9088 27872
rect 9036 27829 9045 27863
rect 9045 27829 9079 27863
rect 9079 27829 9088 27863
rect 9036 27820 9088 27829
rect 10876 27820 10928 27872
rect 11612 27820 11664 27872
rect 14464 27956 14516 28008
rect 17132 28092 17184 28144
rect 15016 28024 15068 28076
rect 15108 27956 15160 28008
rect 18236 28024 18288 28076
rect 18512 28024 18564 28076
rect 16856 27956 16908 28008
rect 18420 27956 18472 28008
rect 19156 28024 19208 28076
rect 20076 28067 20128 28076
rect 20076 28033 20085 28067
rect 20085 28033 20119 28067
rect 20119 28033 20128 28067
rect 20076 28024 20128 28033
rect 21640 28024 21692 28076
rect 23572 28067 23624 28076
rect 23572 28033 23581 28067
rect 23581 28033 23615 28067
rect 23615 28033 23624 28067
rect 23572 28024 23624 28033
rect 23756 28067 23808 28076
rect 23756 28033 23765 28067
rect 23765 28033 23799 28067
rect 23799 28033 23808 28067
rect 23756 28024 23808 28033
rect 25044 28092 25096 28144
rect 26424 28092 26476 28144
rect 27436 28092 27488 28144
rect 28724 28160 28776 28212
rect 30104 28160 30156 28212
rect 30472 28160 30524 28212
rect 19064 27956 19116 28008
rect 25228 28024 25280 28076
rect 25320 28024 25372 28076
rect 14004 27820 14056 27872
rect 14832 27863 14884 27872
rect 14832 27829 14841 27863
rect 14841 27829 14875 27863
rect 14875 27829 14884 27863
rect 14832 27820 14884 27829
rect 15108 27820 15160 27872
rect 15384 27820 15436 27872
rect 16488 27820 16540 27872
rect 18696 27888 18748 27940
rect 23664 27888 23716 27940
rect 25504 27956 25556 28008
rect 25780 28067 25832 28076
rect 25780 28033 25789 28067
rect 25789 28033 25823 28067
rect 25823 28033 25832 28067
rect 25780 28024 25832 28033
rect 26608 28024 26660 28076
rect 27712 28067 27764 28076
rect 27712 28033 27721 28067
rect 27721 28033 27755 28067
rect 27755 28033 27764 28067
rect 27712 28024 27764 28033
rect 27804 28067 27856 28076
rect 27804 28033 27814 28067
rect 27814 28033 27848 28067
rect 27848 28033 27856 28067
rect 27804 28024 27856 28033
rect 19524 27820 19576 27872
rect 21732 27820 21784 27872
rect 22008 27820 22060 27872
rect 24492 27820 24544 27872
rect 24952 27820 25004 27872
rect 25688 27956 25740 28008
rect 27252 27888 27304 27940
rect 26516 27820 26568 27872
rect 28172 28067 28224 28076
rect 28172 28033 28186 28067
rect 28186 28033 28220 28067
rect 28220 28033 28224 28067
rect 28172 28024 28224 28033
rect 28448 28067 28500 28076
rect 28448 28033 28457 28067
rect 28457 28033 28491 28067
rect 28491 28033 28500 28067
rect 28448 28024 28500 28033
rect 28540 27956 28592 28008
rect 29552 28092 29604 28144
rect 29460 28024 29512 28076
rect 29920 28092 29972 28144
rect 33140 28160 33192 28212
rect 33876 28160 33928 28212
rect 37740 28203 37792 28212
rect 37740 28169 37749 28203
rect 37749 28169 37783 28203
rect 37783 28169 37792 28203
rect 37740 28160 37792 28169
rect 37832 28160 37884 28212
rect 39028 28160 39080 28212
rect 39764 28203 39816 28212
rect 39764 28169 39773 28203
rect 39773 28169 39807 28203
rect 39807 28169 39816 28203
rect 39764 28160 39816 28169
rect 30380 28067 30432 28076
rect 30380 28033 30389 28067
rect 30389 28033 30423 28067
rect 30423 28033 30432 28067
rect 30380 28024 30432 28033
rect 31116 28092 31168 28144
rect 29644 27956 29696 28008
rect 30012 27956 30064 28008
rect 30840 28067 30892 28076
rect 30840 28033 30849 28067
rect 30849 28033 30883 28067
rect 30883 28033 30892 28067
rect 30840 28024 30892 28033
rect 31208 28024 31260 28076
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 32772 28092 32824 28144
rect 31852 27956 31904 28008
rect 33600 28024 33652 28076
rect 33876 28024 33928 28076
rect 34336 28092 34388 28144
rect 34428 28135 34480 28144
rect 34428 28101 34437 28135
rect 34437 28101 34471 28135
rect 34471 28101 34480 28135
rect 34428 28092 34480 28101
rect 37372 28092 37424 28144
rect 39396 28092 39448 28144
rect 33508 27956 33560 28008
rect 34704 27956 34756 28008
rect 37556 27999 37608 28008
rect 37556 27965 37565 27999
rect 37565 27965 37599 27999
rect 37599 27965 37608 27999
rect 37556 27956 37608 27965
rect 38016 28024 38068 28076
rect 38476 28067 38528 28076
rect 38476 28033 38485 28067
rect 38485 28033 38519 28067
rect 38519 28033 38528 28067
rect 38476 28024 38528 28033
rect 38660 28067 38712 28076
rect 38660 28033 38669 28067
rect 38669 28033 38703 28067
rect 38703 28033 38712 28067
rect 38660 28024 38712 28033
rect 38844 28067 38896 28076
rect 38844 28033 38853 28067
rect 38853 28033 38887 28067
rect 38887 28033 38896 28067
rect 38844 28024 38896 28033
rect 39028 28067 39080 28076
rect 39028 28033 39037 28067
rect 39037 28033 39071 28067
rect 39071 28033 39080 28067
rect 39028 28024 39080 28033
rect 40040 28024 40092 28076
rect 28632 27888 28684 27940
rect 29092 27888 29144 27940
rect 30196 27888 30248 27940
rect 41512 28067 41564 28076
rect 41512 28033 41521 28067
rect 41521 28033 41555 28067
rect 41555 28033 41564 28067
rect 41512 28024 41564 28033
rect 41880 28067 41932 28076
rect 41880 28033 41889 28067
rect 41889 28033 41923 28067
rect 41923 28033 41932 28067
rect 41880 28024 41932 28033
rect 41696 27931 41748 27940
rect 41696 27897 41705 27931
rect 41705 27897 41739 27931
rect 41739 27897 41748 27931
rect 41696 27888 41748 27897
rect 30104 27863 30156 27872
rect 30104 27829 30113 27863
rect 30113 27829 30147 27863
rect 30147 27829 30156 27863
rect 30104 27820 30156 27829
rect 32128 27863 32180 27872
rect 32128 27829 32137 27863
rect 32137 27829 32171 27863
rect 32171 27829 32180 27863
rect 32128 27820 32180 27829
rect 32588 27863 32640 27872
rect 32588 27829 32597 27863
rect 32597 27829 32631 27863
rect 32631 27829 32640 27863
rect 33784 27863 33836 27872
rect 32588 27820 32640 27829
rect 33784 27829 33793 27863
rect 33793 27829 33827 27863
rect 33827 27829 33836 27863
rect 33784 27820 33836 27829
rect 34520 27820 34572 27872
rect 34612 27863 34664 27872
rect 34612 27829 34621 27863
rect 34621 27829 34655 27863
rect 34655 27829 34664 27863
rect 34612 27820 34664 27829
rect 35164 27820 35216 27872
rect 35532 27820 35584 27872
rect 38200 27863 38252 27872
rect 38200 27829 38209 27863
rect 38209 27829 38243 27863
rect 38243 27829 38252 27863
rect 38200 27820 38252 27829
rect 39396 27820 39448 27872
rect 40408 27820 40460 27872
rect 40592 27863 40644 27872
rect 40592 27829 40601 27863
rect 40601 27829 40635 27863
rect 40635 27829 40644 27863
rect 40592 27820 40644 27829
rect 42064 27863 42116 27872
rect 42064 27829 42073 27863
rect 42073 27829 42107 27863
rect 42107 27829 42116 27863
rect 42064 27820 42116 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4160 27616 4212 27668
rect 4988 27616 5040 27668
rect 4620 27591 4672 27600
rect 4620 27557 4629 27591
rect 4629 27557 4663 27591
rect 4663 27557 4672 27591
rect 4620 27548 4672 27557
rect 5724 27616 5776 27668
rect 10968 27616 11020 27668
rect 3608 27412 3660 27464
rect 8300 27548 8352 27600
rect 9680 27548 9732 27600
rect 6644 27480 6696 27532
rect 2780 27344 2832 27396
rect 4528 27344 4580 27396
rect 7104 27455 7156 27464
rect 7104 27421 7113 27455
rect 7113 27421 7147 27455
rect 7147 27421 7156 27455
rect 7104 27412 7156 27421
rect 8024 27480 8076 27532
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 9036 27523 9088 27532
rect 9036 27489 9045 27523
rect 9045 27489 9079 27523
rect 9079 27489 9088 27523
rect 9036 27480 9088 27489
rect 10876 27523 10928 27532
rect 10876 27489 10885 27523
rect 10885 27489 10919 27523
rect 10919 27489 10928 27523
rect 10876 27480 10928 27489
rect 14464 27591 14516 27600
rect 14464 27557 14473 27591
rect 14473 27557 14507 27591
rect 14507 27557 14516 27591
rect 14464 27548 14516 27557
rect 18236 27616 18288 27668
rect 15200 27548 15252 27600
rect 15292 27591 15344 27600
rect 15292 27557 15301 27591
rect 15301 27557 15335 27591
rect 15335 27557 15344 27591
rect 15292 27548 15344 27557
rect 16856 27548 16908 27600
rect 5172 27344 5224 27396
rect 5356 27344 5408 27396
rect 5724 27344 5776 27396
rect 8116 27387 8168 27396
rect 8116 27353 8125 27387
rect 8125 27353 8159 27387
rect 8159 27353 8168 27387
rect 8116 27344 8168 27353
rect 4804 27276 4856 27328
rect 6920 27276 6972 27328
rect 7932 27276 7984 27328
rect 9404 27412 9456 27464
rect 13912 27480 13964 27532
rect 14924 27480 14976 27532
rect 12716 27455 12768 27464
rect 12716 27421 12725 27455
rect 12725 27421 12759 27455
rect 12759 27421 12768 27455
rect 12716 27412 12768 27421
rect 14648 27455 14700 27464
rect 14648 27421 14657 27455
rect 14657 27421 14691 27455
rect 14691 27421 14700 27455
rect 14648 27412 14700 27421
rect 11060 27344 11112 27396
rect 11152 27387 11204 27396
rect 11152 27353 11161 27387
rect 11161 27353 11195 27387
rect 11195 27353 11204 27387
rect 11152 27344 11204 27353
rect 13360 27344 13412 27396
rect 15016 27455 15068 27464
rect 15016 27421 15025 27455
rect 15025 27421 15059 27455
rect 15059 27421 15068 27455
rect 15016 27412 15068 27421
rect 17868 27548 17920 27600
rect 18880 27616 18932 27668
rect 19432 27616 19484 27668
rect 22376 27616 22428 27668
rect 23112 27616 23164 27668
rect 24492 27616 24544 27668
rect 25228 27616 25280 27668
rect 18420 27548 18472 27600
rect 14832 27344 14884 27396
rect 14924 27387 14976 27396
rect 14924 27353 14933 27387
rect 14933 27353 14967 27387
rect 14967 27353 14976 27387
rect 14924 27344 14976 27353
rect 15568 27344 15620 27396
rect 15660 27387 15712 27396
rect 15660 27353 15669 27387
rect 15669 27353 15703 27387
rect 15703 27353 15712 27387
rect 15660 27344 15712 27353
rect 9312 27276 9364 27328
rect 10140 27276 10192 27328
rect 11980 27276 12032 27328
rect 14372 27276 14424 27328
rect 14464 27276 14516 27328
rect 15108 27319 15160 27328
rect 15108 27285 15117 27319
rect 15117 27285 15151 27319
rect 15151 27285 15160 27319
rect 15108 27276 15160 27285
rect 17040 27344 17092 27396
rect 17132 27276 17184 27328
rect 17408 27276 17460 27328
rect 17960 27412 18012 27464
rect 18236 27480 18288 27532
rect 19156 27480 19208 27532
rect 20076 27548 20128 27600
rect 22008 27591 22060 27600
rect 22008 27557 22017 27591
rect 22017 27557 22051 27591
rect 22051 27557 22060 27591
rect 22008 27548 22060 27557
rect 27252 27616 27304 27668
rect 27620 27616 27672 27668
rect 30840 27616 30892 27668
rect 32128 27616 32180 27668
rect 27160 27548 27212 27600
rect 17776 27387 17828 27396
rect 17776 27353 17785 27387
rect 17785 27353 17819 27387
rect 17819 27353 17828 27387
rect 17776 27344 17828 27353
rect 17960 27319 18012 27328
rect 17960 27285 17969 27319
rect 17969 27285 18003 27319
rect 18003 27285 18012 27319
rect 17960 27276 18012 27285
rect 18144 27319 18196 27328
rect 18144 27285 18153 27319
rect 18153 27285 18187 27319
rect 18187 27285 18196 27319
rect 18144 27276 18196 27285
rect 20536 27455 20588 27464
rect 20536 27421 20545 27455
rect 20545 27421 20579 27455
rect 20579 27421 20588 27455
rect 20536 27412 20588 27421
rect 21640 27480 21692 27532
rect 23020 27523 23072 27532
rect 18328 27276 18380 27328
rect 20076 27344 20128 27396
rect 20444 27344 20496 27396
rect 21824 27455 21876 27464
rect 21824 27421 21833 27455
rect 21833 27421 21867 27455
rect 21867 27421 21876 27455
rect 21824 27412 21876 27421
rect 22100 27455 22152 27464
rect 22100 27421 22109 27455
rect 22109 27421 22143 27455
rect 22143 27421 22152 27455
rect 23020 27489 23029 27523
rect 23029 27489 23063 27523
rect 23063 27489 23072 27523
rect 23020 27480 23072 27489
rect 23848 27480 23900 27532
rect 24400 27523 24452 27532
rect 24400 27489 24409 27523
rect 24409 27489 24443 27523
rect 24443 27489 24452 27523
rect 24400 27480 24452 27489
rect 24676 27480 24728 27532
rect 22100 27412 22152 27421
rect 26516 27455 26568 27464
rect 26516 27421 26525 27455
rect 26525 27421 26559 27455
rect 26559 27421 26568 27455
rect 27528 27480 27580 27532
rect 29184 27548 29236 27600
rect 30656 27548 30708 27600
rect 33600 27616 33652 27668
rect 28632 27480 28684 27532
rect 26516 27412 26568 27421
rect 28816 27455 28868 27464
rect 28816 27421 28825 27455
rect 28825 27421 28859 27455
rect 28859 27421 28868 27455
rect 28816 27412 28868 27421
rect 29276 27480 29328 27532
rect 29920 27480 29972 27532
rect 31668 27523 31720 27532
rect 31668 27489 31677 27523
rect 31677 27489 31711 27523
rect 31711 27489 31720 27523
rect 31668 27480 31720 27489
rect 33508 27591 33560 27600
rect 33508 27557 33517 27591
rect 33517 27557 33551 27591
rect 33551 27557 33560 27591
rect 33508 27548 33560 27557
rect 33784 27616 33836 27668
rect 35532 27616 35584 27668
rect 35992 27616 36044 27668
rect 37740 27659 37792 27668
rect 37740 27625 37749 27659
rect 37749 27625 37783 27659
rect 37783 27625 37792 27659
rect 37740 27616 37792 27625
rect 40592 27616 40644 27668
rect 41880 27659 41932 27668
rect 41880 27625 41889 27659
rect 41889 27625 41923 27659
rect 41923 27625 41932 27659
rect 41880 27616 41932 27625
rect 33876 27548 33928 27600
rect 33968 27548 34020 27600
rect 34152 27548 34204 27600
rect 29184 27455 29236 27464
rect 29184 27421 29193 27455
rect 29193 27421 29227 27455
rect 29227 27421 29236 27455
rect 29184 27412 29236 27421
rect 30656 27455 30708 27464
rect 30656 27421 30665 27455
rect 30665 27421 30699 27455
rect 30699 27421 30708 27455
rect 30656 27412 30708 27421
rect 30840 27412 30892 27464
rect 30932 27455 30984 27464
rect 30932 27421 30941 27455
rect 30941 27421 30975 27455
rect 30975 27421 30984 27455
rect 30932 27412 30984 27421
rect 33048 27412 33100 27464
rect 33232 27412 33284 27464
rect 33784 27455 33836 27464
rect 33784 27421 33793 27455
rect 33793 27421 33827 27455
rect 33827 27421 33836 27455
rect 33784 27412 33836 27421
rect 34336 27480 34388 27532
rect 34612 27480 34664 27532
rect 35348 27548 35400 27600
rect 35532 27480 35584 27532
rect 22560 27344 22612 27396
rect 22836 27387 22888 27396
rect 22836 27353 22845 27387
rect 22845 27353 22879 27387
rect 22879 27353 22888 27387
rect 22836 27344 22888 27353
rect 26240 27344 26292 27396
rect 18512 27319 18564 27328
rect 18512 27285 18521 27319
rect 18521 27285 18555 27319
rect 18555 27285 18564 27319
rect 18512 27276 18564 27285
rect 18604 27276 18656 27328
rect 19064 27276 19116 27328
rect 23020 27276 23072 27328
rect 31024 27344 31076 27396
rect 31484 27387 31536 27396
rect 31484 27353 31493 27387
rect 31493 27353 31527 27387
rect 31527 27353 31536 27387
rect 31484 27344 31536 27353
rect 30380 27276 30432 27328
rect 31208 27319 31260 27328
rect 31208 27285 31217 27319
rect 31217 27285 31251 27319
rect 31251 27285 31260 27319
rect 31208 27276 31260 27285
rect 33876 27276 33928 27328
rect 34428 27455 34480 27464
rect 34428 27421 34437 27455
rect 34437 27421 34471 27455
rect 34471 27421 34480 27455
rect 34428 27412 34480 27421
rect 35256 27412 35308 27464
rect 37280 27548 37332 27600
rect 38384 27548 38436 27600
rect 40040 27548 40092 27600
rect 38660 27480 38712 27532
rect 35532 27344 35584 27396
rect 34060 27276 34112 27328
rect 34704 27319 34756 27328
rect 34704 27285 34713 27319
rect 34713 27285 34747 27319
rect 34747 27285 34756 27319
rect 34704 27276 34756 27285
rect 35992 27455 36044 27464
rect 35992 27421 36001 27455
rect 36001 27421 36035 27455
rect 36035 27421 36044 27455
rect 35992 27412 36044 27421
rect 39304 27455 39356 27464
rect 39304 27421 39313 27455
rect 39313 27421 39347 27455
rect 39347 27421 39356 27455
rect 39304 27412 39356 27421
rect 40132 27455 40184 27464
rect 40132 27421 40141 27455
rect 40141 27421 40175 27455
rect 40175 27421 40184 27455
rect 40132 27412 40184 27421
rect 39028 27344 39080 27396
rect 39396 27387 39448 27396
rect 39396 27353 39405 27387
rect 39405 27353 39439 27387
rect 39439 27353 39448 27387
rect 39396 27344 39448 27353
rect 39488 27387 39540 27396
rect 39488 27353 39497 27387
rect 39497 27353 39531 27387
rect 39531 27353 39540 27387
rect 39488 27344 39540 27353
rect 39856 27344 39908 27396
rect 39948 27344 40000 27396
rect 36636 27276 36688 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 4620 27072 4672 27124
rect 4896 27072 4948 27124
rect 5448 27115 5500 27124
rect 5448 27081 5457 27115
rect 5457 27081 5491 27115
rect 5491 27081 5500 27115
rect 5448 27072 5500 27081
rect 5724 27072 5776 27124
rect 4160 26979 4212 26988
rect 4160 26945 4169 26979
rect 4169 26945 4203 26979
rect 4203 26945 4212 26979
rect 4160 26936 4212 26945
rect 9036 27004 9088 27056
rect 9312 27115 9364 27124
rect 9312 27081 9321 27115
rect 9321 27081 9355 27115
rect 9355 27081 9364 27115
rect 9312 27072 9364 27081
rect 11152 27072 11204 27124
rect 11980 27115 12032 27124
rect 11980 27081 11989 27115
rect 11989 27081 12023 27115
rect 12023 27081 12032 27115
rect 11980 27072 12032 27081
rect 15016 27115 15068 27124
rect 15016 27081 15025 27115
rect 15025 27081 15059 27115
rect 15059 27081 15068 27115
rect 15016 27072 15068 27081
rect 15660 27072 15712 27124
rect 16304 27115 16356 27124
rect 16304 27081 16313 27115
rect 16313 27081 16347 27115
rect 16347 27081 16356 27115
rect 16304 27072 16356 27081
rect 16764 27072 16816 27124
rect 16948 27072 17000 27124
rect 18328 27072 18380 27124
rect 19432 27072 19484 27124
rect 19524 27072 19576 27124
rect 12716 27004 12768 27056
rect 14556 27004 14608 27056
rect 15936 27004 15988 27056
rect 17868 27004 17920 27056
rect 18880 27004 18932 27056
rect 20628 27072 20680 27124
rect 21824 27072 21876 27124
rect 23020 27115 23072 27124
rect 23020 27081 23029 27115
rect 23029 27081 23063 27115
rect 23063 27081 23072 27115
rect 23020 27072 23072 27081
rect 25228 27072 25280 27124
rect 27160 27072 27212 27124
rect 29184 27072 29236 27124
rect 29644 27072 29696 27124
rect 32128 27072 32180 27124
rect 34428 27072 34480 27124
rect 2780 26868 2832 26920
rect 3424 26800 3476 26852
rect 4712 26800 4764 26852
rect 4988 26979 5040 26988
rect 4988 26945 4997 26979
rect 4997 26945 5031 26979
rect 5031 26945 5040 26979
rect 4988 26936 5040 26945
rect 6552 26936 6604 26988
rect 9496 26936 9548 26988
rect 10692 26936 10744 26988
rect 10876 26936 10928 26988
rect 5632 26868 5684 26920
rect 5540 26800 5592 26852
rect 5724 26800 5776 26852
rect 2872 26732 2924 26784
rect 4528 26732 4580 26784
rect 4988 26732 5040 26784
rect 5448 26732 5500 26784
rect 8668 26732 8720 26784
rect 9404 26775 9456 26784
rect 9404 26741 9413 26775
rect 9413 26741 9447 26775
rect 9447 26741 9456 26775
rect 9404 26732 9456 26741
rect 10140 26732 10192 26784
rect 16304 26936 16356 26988
rect 16856 26936 16908 26988
rect 17776 26979 17828 26988
rect 17776 26945 17785 26979
rect 17785 26945 17819 26979
rect 17819 26945 17828 26979
rect 17776 26936 17828 26945
rect 17960 26979 18012 26988
rect 17960 26945 17969 26979
rect 17969 26945 18003 26979
rect 18003 26945 18012 26979
rect 17960 26936 18012 26945
rect 18144 26936 18196 26988
rect 18420 26979 18472 26988
rect 18420 26945 18429 26979
rect 18429 26945 18463 26979
rect 18463 26945 18472 26979
rect 18972 26979 19024 26988
rect 18420 26936 18472 26945
rect 18972 26945 18981 26979
rect 18981 26945 19015 26979
rect 19015 26945 19024 26979
rect 18972 26936 19024 26945
rect 19156 26936 19208 26988
rect 19892 26979 19944 26988
rect 19892 26945 19901 26979
rect 19901 26945 19935 26979
rect 19935 26945 19944 26979
rect 20536 27004 20588 27056
rect 19892 26936 19944 26945
rect 12072 26911 12124 26920
rect 12072 26877 12081 26911
rect 12081 26877 12115 26911
rect 12115 26877 12124 26911
rect 12072 26868 12124 26877
rect 15384 26868 15436 26920
rect 16672 26911 16724 26920
rect 16672 26877 16681 26911
rect 16681 26877 16715 26911
rect 16715 26877 16724 26911
rect 16672 26868 16724 26877
rect 12624 26800 12676 26852
rect 15752 26800 15804 26852
rect 16948 26868 17000 26920
rect 14832 26732 14884 26784
rect 15292 26732 15344 26784
rect 15844 26732 15896 26784
rect 16948 26732 17000 26784
rect 17316 26868 17368 26920
rect 18328 26868 18380 26920
rect 26700 27004 26752 27056
rect 23480 26936 23532 26988
rect 24400 26936 24452 26988
rect 25504 26936 25556 26988
rect 17500 26800 17552 26852
rect 18604 26800 18656 26852
rect 17684 26732 17736 26784
rect 17776 26732 17828 26784
rect 18696 26732 18748 26784
rect 20260 26800 20312 26852
rect 20720 26868 20772 26920
rect 21180 26868 21232 26920
rect 22560 26868 22612 26920
rect 23112 26868 23164 26920
rect 20444 26800 20496 26852
rect 20812 26800 20864 26852
rect 22100 26800 22152 26852
rect 25320 26911 25372 26920
rect 25320 26877 25329 26911
rect 25329 26877 25363 26911
rect 25363 26877 25372 26911
rect 25320 26868 25372 26877
rect 25412 26868 25464 26920
rect 25780 26868 25832 26920
rect 26424 26979 26476 26988
rect 26424 26945 26433 26979
rect 26433 26945 26467 26979
rect 26467 26945 26476 26979
rect 26424 26936 26476 26945
rect 26516 26979 26568 26988
rect 26516 26945 26525 26979
rect 26525 26945 26559 26979
rect 26559 26945 26568 26979
rect 26516 26936 26568 26945
rect 27896 26868 27948 26920
rect 29736 27004 29788 27056
rect 30656 27004 30708 27056
rect 33876 27004 33928 27056
rect 34520 27004 34572 27056
rect 28356 26936 28408 26988
rect 22468 26732 22520 26784
rect 22928 26732 22980 26784
rect 23112 26732 23164 26784
rect 24216 26732 24268 26784
rect 25596 26732 25648 26784
rect 26700 26775 26752 26784
rect 26700 26741 26709 26775
rect 26709 26741 26743 26775
rect 26743 26741 26752 26775
rect 26700 26732 26752 26741
rect 27804 26800 27856 26852
rect 28908 26979 28960 26988
rect 28908 26945 28917 26979
rect 28917 26945 28951 26979
rect 28951 26945 28960 26979
rect 28908 26936 28960 26945
rect 29000 26979 29052 26988
rect 29000 26945 29009 26979
rect 29009 26945 29043 26979
rect 29043 26945 29052 26979
rect 29000 26936 29052 26945
rect 28816 26868 28868 26920
rect 29920 26979 29972 26988
rect 29920 26945 29929 26979
rect 29929 26945 29963 26979
rect 29963 26945 29972 26979
rect 29920 26936 29972 26945
rect 35808 27072 35860 27124
rect 35532 27047 35584 27056
rect 35532 27013 35541 27047
rect 35541 27013 35575 27047
rect 35575 27013 35584 27047
rect 35532 27004 35584 27013
rect 32772 26868 32824 26920
rect 33600 26868 33652 26920
rect 34060 26868 34112 26920
rect 34520 26868 34572 26920
rect 35624 26979 35676 26988
rect 35624 26945 35633 26979
rect 35633 26945 35667 26979
rect 35667 26945 35676 26979
rect 35624 26936 35676 26945
rect 36268 27072 36320 27124
rect 36636 27115 36688 27124
rect 36636 27081 36645 27115
rect 36645 27081 36679 27115
rect 36679 27081 36688 27115
rect 36636 27072 36688 27081
rect 37740 27072 37792 27124
rect 40040 27115 40092 27124
rect 40040 27081 40049 27115
rect 40049 27081 40083 27115
rect 40083 27081 40092 27115
rect 40040 27072 40092 27081
rect 40868 27072 40920 27124
rect 41604 27072 41656 27124
rect 36176 26979 36228 26988
rect 36176 26945 36183 26979
rect 36183 26945 36228 26979
rect 36176 26936 36228 26945
rect 36544 27004 36596 27056
rect 38384 27047 38436 27056
rect 38384 27013 38393 27047
rect 38393 27013 38427 27047
rect 38427 27013 38436 27047
rect 38384 27004 38436 27013
rect 38568 27004 38620 27056
rect 36360 26979 36412 26988
rect 36360 26945 36369 26979
rect 36369 26945 36403 26979
rect 36403 26945 36412 26979
rect 36360 26936 36412 26945
rect 36452 26979 36504 26988
rect 36452 26945 36466 26979
rect 36466 26945 36500 26979
rect 36500 26945 36504 26979
rect 36452 26936 36504 26945
rect 40592 26979 40644 26988
rect 40592 26945 40601 26979
rect 40601 26945 40635 26979
rect 40635 26945 40644 26979
rect 40592 26936 40644 26945
rect 40776 26979 40828 26988
rect 40776 26945 40785 26979
rect 40785 26945 40819 26979
rect 40819 26945 40828 26979
rect 40776 26936 40828 26945
rect 41052 26936 41104 26988
rect 35256 26843 35308 26852
rect 35256 26809 35265 26843
rect 35265 26809 35299 26843
rect 35299 26809 35308 26843
rect 35256 26800 35308 26809
rect 28724 26732 28776 26784
rect 30012 26732 30064 26784
rect 30196 26775 30248 26784
rect 30196 26741 30226 26775
rect 30226 26741 30248 26775
rect 30196 26732 30248 26741
rect 30656 26732 30708 26784
rect 31208 26732 31260 26784
rect 31668 26775 31720 26784
rect 31668 26741 31677 26775
rect 31677 26741 31711 26775
rect 31711 26741 31720 26775
rect 31668 26732 31720 26741
rect 34612 26732 34664 26784
rect 36728 26868 36780 26920
rect 35716 26800 35768 26852
rect 37556 26800 37608 26852
rect 41236 26800 41288 26852
rect 36084 26732 36136 26784
rect 39212 26732 39264 26784
rect 40684 26732 40736 26784
rect 42064 26775 42116 26784
rect 42064 26741 42073 26775
rect 42073 26741 42107 26775
rect 42107 26741 42116 26775
rect 42064 26732 42116 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3424 26528 3476 26580
rect 4436 26571 4488 26580
rect 4436 26537 4445 26571
rect 4445 26537 4479 26571
rect 4479 26537 4488 26571
rect 4436 26528 4488 26537
rect 4712 26528 4764 26580
rect 5356 26528 5408 26580
rect 8484 26528 8536 26580
rect 9220 26528 9272 26580
rect 9496 26571 9548 26580
rect 9496 26537 9505 26571
rect 9505 26537 9539 26571
rect 9539 26537 9548 26571
rect 9496 26528 9548 26537
rect 9588 26528 9640 26580
rect 11336 26528 11388 26580
rect 12164 26528 12216 26580
rect 12992 26528 13044 26580
rect 14924 26528 14976 26580
rect 7932 26503 7984 26512
rect 7932 26469 7941 26503
rect 7941 26469 7975 26503
rect 7975 26469 7984 26503
rect 7932 26460 7984 26469
rect 10232 26460 10284 26512
rect 16304 26528 16356 26580
rect 17960 26528 18012 26580
rect 20444 26528 20496 26580
rect 2780 26392 2832 26444
rect 3516 26367 3568 26376
rect 3516 26333 3525 26367
rect 3525 26333 3559 26367
rect 3559 26333 3568 26367
rect 3516 26324 3568 26333
rect 3976 26324 4028 26376
rect 2964 26256 3016 26308
rect 4896 26324 4948 26376
rect 5080 26367 5132 26376
rect 5080 26333 5084 26367
rect 5084 26333 5118 26367
rect 5118 26333 5132 26367
rect 5080 26324 5132 26333
rect 7012 26392 7064 26444
rect 4804 26256 4856 26308
rect 5540 26367 5592 26376
rect 5540 26333 5549 26367
rect 5549 26333 5583 26367
rect 5583 26333 5592 26367
rect 5540 26324 5592 26333
rect 5724 26367 5776 26376
rect 5724 26333 5733 26367
rect 5733 26333 5767 26367
rect 5767 26333 5776 26367
rect 5724 26324 5776 26333
rect 6000 26324 6052 26376
rect 6184 26367 6236 26376
rect 6184 26333 6193 26367
rect 6193 26333 6227 26367
rect 6227 26333 6236 26367
rect 6184 26324 6236 26333
rect 6644 26367 6696 26376
rect 6644 26333 6653 26367
rect 6653 26333 6687 26367
rect 6687 26333 6696 26367
rect 6644 26324 6696 26333
rect 6920 26367 6972 26376
rect 6920 26333 6929 26367
rect 6929 26333 6963 26367
rect 6963 26333 6972 26367
rect 6920 26324 6972 26333
rect 7196 26324 7248 26376
rect 8300 26324 8352 26376
rect 8484 26367 8536 26376
rect 8484 26333 8493 26367
rect 8493 26333 8527 26367
rect 8527 26333 8536 26367
rect 8484 26324 8536 26333
rect 8944 26367 8996 26376
rect 8944 26333 8953 26367
rect 8953 26333 8987 26367
rect 8987 26333 8996 26367
rect 8944 26324 8996 26333
rect 9220 26367 9272 26376
rect 9220 26333 9229 26367
rect 9229 26333 9263 26367
rect 9263 26333 9272 26367
rect 9220 26324 9272 26333
rect 10140 26392 10192 26444
rect 10692 26392 10744 26444
rect 9588 26367 9640 26376
rect 9588 26333 9597 26367
rect 9597 26333 9631 26367
rect 9631 26333 9640 26367
rect 9588 26324 9640 26333
rect 13176 26392 13228 26444
rect 17408 26460 17460 26512
rect 18328 26460 18380 26512
rect 18972 26460 19024 26512
rect 13912 26435 13964 26444
rect 13912 26401 13921 26435
rect 13921 26401 13955 26435
rect 13955 26401 13964 26435
rect 13912 26392 13964 26401
rect 14924 26392 14976 26444
rect 15476 26435 15528 26444
rect 15476 26401 15485 26435
rect 15485 26401 15519 26435
rect 15519 26401 15528 26435
rect 15476 26392 15528 26401
rect 16396 26392 16448 26444
rect 16856 26392 16908 26444
rect 18144 26392 18196 26444
rect 18236 26435 18288 26444
rect 18236 26401 18245 26435
rect 18245 26401 18279 26435
rect 18279 26401 18288 26435
rect 18236 26392 18288 26401
rect 15660 26324 15712 26376
rect 15752 26367 15804 26376
rect 15752 26333 15761 26367
rect 15761 26333 15795 26367
rect 15795 26333 15804 26367
rect 15752 26324 15804 26333
rect 15844 26367 15896 26376
rect 15844 26333 15853 26367
rect 15853 26333 15887 26367
rect 15887 26333 15896 26367
rect 15844 26324 15896 26333
rect 4160 26188 4212 26240
rect 4528 26188 4580 26240
rect 5448 26188 5500 26240
rect 10692 26188 10744 26240
rect 13176 26256 13228 26308
rect 13728 26256 13780 26308
rect 16028 26324 16080 26376
rect 16120 26299 16172 26308
rect 16120 26265 16129 26299
rect 16129 26265 16163 26299
rect 16163 26265 16172 26299
rect 16120 26256 16172 26265
rect 16304 26367 16356 26376
rect 16304 26333 16318 26367
rect 16318 26333 16352 26367
rect 16352 26333 16356 26367
rect 16304 26324 16356 26333
rect 17040 26324 17092 26376
rect 17224 26367 17276 26376
rect 17224 26333 17233 26367
rect 17233 26333 17267 26367
rect 17267 26333 17276 26367
rect 17224 26324 17276 26333
rect 17408 26367 17460 26376
rect 17408 26333 17417 26367
rect 17417 26333 17451 26367
rect 17451 26333 17460 26367
rect 17408 26324 17460 26333
rect 17776 26299 17828 26308
rect 17776 26265 17794 26299
rect 17794 26265 17828 26299
rect 17776 26256 17828 26265
rect 17960 26367 18012 26376
rect 17960 26333 17969 26367
rect 17969 26333 18003 26367
rect 18003 26333 18012 26367
rect 17960 26324 18012 26333
rect 18420 26324 18472 26376
rect 18512 26367 18564 26376
rect 18512 26333 18521 26367
rect 18521 26333 18555 26367
rect 18555 26333 18564 26367
rect 18512 26324 18564 26333
rect 20260 26392 20312 26444
rect 20628 26392 20680 26444
rect 19892 26256 19944 26308
rect 20536 26299 20588 26308
rect 20536 26265 20570 26299
rect 20570 26265 20588 26299
rect 20536 26256 20588 26265
rect 11520 26188 11572 26240
rect 11980 26188 12032 26240
rect 14556 26188 14608 26240
rect 15752 26188 15804 26240
rect 17592 26231 17644 26240
rect 17592 26197 17601 26231
rect 17601 26197 17635 26231
rect 17635 26197 17644 26231
rect 17592 26188 17644 26197
rect 17868 26188 17920 26240
rect 19524 26188 19576 26240
rect 21548 26324 21600 26376
rect 22284 26324 22336 26376
rect 22560 26528 22612 26580
rect 23388 26460 23440 26512
rect 23112 26435 23164 26444
rect 23112 26401 23121 26435
rect 23121 26401 23155 26435
rect 23155 26401 23164 26435
rect 23112 26392 23164 26401
rect 23572 26435 23624 26444
rect 23572 26401 23581 26435
rect 23581 26401 23615 26435
rect 23615 26401 23624 26435
rect 23572 26392 23624 26401
rect 23848 26460 23900 26512
rect 23388 26324 23440 26376
rect 23756 26324 23808 26376
rect 24400 26392 24452 26444
rect 27896 26460 27948 26512
rect 28908 26460 28960 26512
rect 30196 26528 30248 26580
rect 31300 26528 31352 26580
rect 31484 26528 31536 26580
rect 32956 26528 33008 26580
rect 33140 26528 33192 26580
rect 33692 26528 33744 26580
rect 33876 26528 33928 26580
rect 34152 26571 34204 26580
rect 34152 26537 34161 26571
rect 34161 26537 34195 26571
rect 34195 26537 34204 26571
rect 34152 26528 34204 26537
rect 34244 26528 34296 26580
rect 31760 26460 31812 26512
rect 31944 26503 31996 26512
rect 31944 26469 31953 26503
rect 31953 26469 31987 26503
rect 31987 26469 31996 26503
rect 31944 26460 31996 26469
rect 32128 26460 32180 26512
rect 29092 26392 29144 26444
rect 29276 26392 29328 26444
rect 30840 26392 30892 26444
rect 24216 26324 24268 26376
rect 26240 26324 26292 26376
rect 29736 26324 29788 26376
rect 30288 26367 30340 26376
rect 30288 26333 30297 26367
rect 30297 26333 30331 26367
rect 30331 26333 30340 26367
rect 30288 26324 30340 26333
rect 30380 26367 30432 26376
rect 30380 26333 30389 26367
rect 30389 26333 30423 26367
rect 30423 26333 30432 26367
rect 30380 26324 30432 26333
rect 30748 26324 30800 26376
rect 21272 26231 21324 26240
rect 21272 26197 21281 26231
rect 21281 26197 21315 26231
rect 21315 26197 21324 26231
rect 21272 26188 21324 26197
rect 21456 26231 21508 26240
rect 21456 26197 21465 26231
rect 21465 26197 21499 26231
rect 21499 26197 21508 26231
rect 21456 26188 21508 26197
rect 22100 26231 22152 26240
rect 22100 26197 22109 26231
rect 22109 26197 22143 26231
rect 22143 26197 22152 26231
rect 22100 26188 22152 26197
rect 22192 26188 22244 26240
rect 24860 26256 24912 26308
rect 22560 26188 22612 26240
rect 23572 26231 23624 26240
rect 23572 26197 23581 26231
rect 23581 26197 23615 26231
rect 23615 26197 23624 26231
rect 23572 26188 23624 26197
rect 25504 26188 25556 26240
rect 31024 26324 31076 26376
rect 31484 26367 31536 26376
rect 31484 26333 31491 26367
rect 31491 26333 31536 26367
rect 31484 26324 31536 26333
rect 32680 26392 32732 26444
rect 33784 26392 33836 26444
rect 40040 26528 40092 26580
rect 31760 26367 31812 26376
rect 31760 26333 31774 26367
rect 31774 26333 31808 26367
rect 31808 26333 31812 26367
rect 31760 26324 31812 26333
rect 33600 26367 33652 26376
rect 33600 26333 33609 26367
rect 33609 26333 33643 26367
rect 33643 26333 33652 26367
rect 33600 26324 33652 26333
rect 35716 26392 35768 26444
rect 37096 26460 37148 26512
rect 39304 26460 39356 26512
rect 32772 26256 32824 26308
rect 33784 26299 33836 26308
rect 33784 26265 33793 26299
rect 33793 26265 33827 26299
rect 33827 26265 33836 26299
rect 33784 26256 33836 26265
rect 31668 26188 31720 26240
rect 33232 26188 33284 26240
rect 34428 26324 34480 26376
rect 34612 26256 34664 26308
rect 34796 26256 34848 26308
rect 36084 26367 36136 26376
rect 36084 26333 36093 26367
rect 36093 26333 36127 26367
rect 36127 26333 36136 26367
rect 36084 26324 36136 26333
rect 36360 26367 36412 26376
rect 36360 26333 36369 26367
rect 36369 26333 36403 26367
rect 36403 26333 36412 26367
rect 36360 26324 36412 26333
rect 36452 26367 36504 26376
rect 36452 26333 36461 26367
rect 36461 26333 36495 26367
rect 36495 26333 36504 26367
rect 36452 26324 36504 26333
rect 36728 26367 36780 26376
rect 36728 26333 36737 26367
rect 36737 26333 36771 26367
rect 36771 26333 36780 26367
rect 36728 26324 36780 26333
rect 36820 26324 36872 26376
rect 37004 26367 37056 26376
rect 37004 26333 37013 26367
rect 37013 26333 37047 26367
rect 37047 26333 37056 26367
rect 37004 26324 37056 26333
rect 40132 26392 40184 26444
rect 40684 26435 40736 26444
rect 40684 26401 40693 26435
rect 40693 26401 40727 26435
rect 40727 26401 40736 26435
rect 40684 26392 40736 26401
rect 41052 26392 41104 26444
rect 36268 26299 36320 26308
rect 36268 26265 36277 26299
rect 36277 26265 36311 26299
rect 36311 26265 36320 26299
rect 36268 26256 36320 26265
rect 36452 26188 36504 26240
rect 37188 26256 37240 26308
rect 38292 26367 38344 26376
rect 38292 26333 38301 26367
rect 38301 26333 38335 26367
rect 38335 26333 38344 26367
rect 38292 26324 38344 26333
rect 39028 26367 39080 26376
rect 39028 26333 39037 26367
rect 39037 26333 39071 26367
rect 39071 26333 39080 26367
rect 39028 26324 39080 26333
rect 37556 26188 37608 26240
rect 39120 26256 39172 26308
rect 39580 26256 39632 26308
rect 39948 26256 40000 26308
rect 39488 26188 39540 26240
rect 40224 26188 40276 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 848 25984 900 26036
rect 4712 25984 4764 26036
rect 5724 25984 5776 26036
rect 6092 25984 6144 26036
rect 7104 26027 7156 26036
rect 7104 25993 7113 26027
rect 7113 25993 7147 26027
rect 7147 25993 7156 26027
rect 7104 25984 7156 25993
rect 8300 26027 8352 26036
rect 8300 25993 8309 26027
rect 8309 25993 8343 26027
rect 8343 25993 8352 26027
rect 8300 25984 8352 25993
rect 2688 25891 2740 25900
rect 2688 25857 2697 25891
rect 2697 25857 2731 25891
rect 2731 25857 2740 25891
rect 2688 25848 2740 25857
rect 2780 25848 2832 25900
rect 3792 25848 3844 25900
rect 3608 25780 3660 25832
rect 3976 25891 4028 25900
rect 3976 25857 3986 25891
rect 3986 25857 4020 25891
rect 4020 25857 4028 25891
rect 3976 25848 4028 25857
rect 4436 25848 4488 25900
rect 4712 25848 4764 25900
rect 5356 25848 5408 25900
rect 5816 25891 5868 25900
rect 5816 25857 5825 25891
rect 5825 25857 5859 25891
rect 5859 25857 5868 25891
rect 5816 25848 5868 25857
rect 6000 25848 6052 25900
rect 6092 25891 6144 25900
rect 6092 25857 6101 25891
rect 6101 25857 6135 25891
rect 6135 25857 6144 25891
rect 6092 25848 6144 25857
rect 4620 25780 4672 25832
rect 4804 25780 4856 25832
rect 4528 25712 4580 25764
rect 5632 25755 5684 25764
rect 5632 25721 5641 25755
rect 5641 25721 5675 25755
rect 5675 25721 5684 25755
rect 5632 25712 5684 25721
rect 5908 25712 5960 25764
rect 4712 25644 4764 25696
rect 5724 25687 5776 25696
rect 5724 25653 5733 25687
rect 5733 25653 5767 25687
rect 5767 25653 5776 25687
rect 5724 25644 5776 25653
rect 6368 25644 6420 25696
rect 8668 25959 8720 25968
rect 8668 25925 8677 25959
rect 8677 25925 8711 25959
rect 8711 25925 8720 25959
rect 8668 25916 8720 25925
rect 8944 26027 8996 26036
rect 8944 25993 8953 26027
rect 8953 25993 8987 26027
rect 8987 25993 8996 26027
rect 8944 25984 8996 25993
rect 9588 25984 9640 26036
rect 11520 26027 11572 26036
rect 11520 25993 11529 26027
rect 11529 25993 11563 26027
rect 11563 25993 11572 26027
rect 11520 25984 11572 25993
rect 12164 25984 12216 26036
rect 14740 26027 14792 26036
rect 14740 25993 14749 26027
rect 14749 25993 14783 26027
rect 14783 25993 14792 26027
rect 14740 25984 14792 25993
rect 14924 26027 14976 26036
rect 14924 25993 14933 26027
rect 14933 25993 14967 26027
rect 14967 25993 14976 26027
rect 14924 25984 14976 25993
rect 16304 25984 16356 26036
rect 16488 25984 16540 26036
rect 18236 25984 18288 26036
rect 10232 25916 10284 25968
rect 10692 25916 10744 25968
rect 15568 25916 15620 25968
rect 16396 25916 16448 25968
rect 7288 25891 7340 25900
rect 7288 25857 7297 25891
rect 7297 25857 7331 25891
rect 7331 25857 7340 25891
rect 7288 25848 7340 25857
rect 7380 25891 7432 25900
rect 7380 25857 7389 25891
rect 7389 25857 7423 25891
rect 7423 25857 7432 25891
rect 7380 25848 7432 25857
rect 7656 25891 7708 25900
rect 7656 25857 7665 25891
rect 7665 25857 7699 25891
rect 7699 25857 7708 25891
rect 7656 25848 7708 25857
rect 7932 25891 7984 25900
rect 7932 25857 7941 25891
rect 7941 25857 7975 25891
rect 7975 25857 7984 25891
rect 7932 25848 7984 25857
rect 8024 25780 8076 25832
rect 8392 25891 8444 25900
rect 8392 25857 8401 25891
rect 8401 25857 8435 25891
rect 8435 25857 8444 25891
rect 8392 25848 8444 25857
rect 8576 25891 8628 25900
rect 8576 25857 8585 25891
rect 8585 25857 8619 25891
rect 8619 25857 8628 25891
rect 8576 25848 8628 25857
rect 8852 25848 8904 25900
rect 10784 25891 10836 25900
rect 10784 25857 10793 25891
rect 10793 25857 10827 25891
rect 10827 25857 10836 25891
rect 10784 25848 10836 25857
rect 12440 25848 12492 25900
rect 12808 25848 12860 25900
rect 14372 25891 14424 25900
rect 14372 25857 14381 25891
rect 14381 25857 14415 25891
rect 14415 25857 14424 25891
rect 14372 25848 14424 25857
rect 14556 25891 14608 25900
rect 14556 25857 14569 25891
rect 14569 25857 14608 25891
rect 14556 25848 14608 25857
rect 14832 25891 14884 25900
rect 14832 25857 14841 25891
rect 14841 25857 14875 25891
rect 14875 25857 14884 25891
rect 14832 25848 14884 25857
rect 15016 25891 15068 25900
rect 15016 25857 15025 25891
rect 15025 25857 15059 25891
rect 15059 25857 15068 25891
rect 15016 25848 15068 25857
rect 12164 25823 12216 25832
rect 12164 25789 12173 25823
rect 12173 25789 12207 25823
rect 12207 25789 12216 25823
rect 12164 25780 12216 25789
rect 14924 25780 14976 25832
rect 15292 25848 15344 25900
rect 15476 25891 15528 25900
rect 15476 25857 15485 25891
rect 15485 25857 15519 25891
rect 15519 25857 15528 25891
rect 15476 25848 15528 25857
rect 16028 25780 16080 25832
rect 17960 25848 18012 25900
rect 19432 25848 19484 25900
rect 20444 25916 20496 25968
rect 17040 25780 17092 25832
rect 19524 25780 19576 25832
rect 20168 25848 20220 25900
rect 20536 25848 20588 25900
rect 21180 25916 21232 25968
rect 21824 25984 21876 26036
rect 21456 25959 21508 25968
rect 21456 25925 21465 25959
rect 21465 25925 21499 25959
rect 21499 25925 21508 25959
rect 21456 25916 21508 25925
rect 22100 25916 22152 25968
rect 20260 25823 20312 25832
rect 20260 25789 20269 25823
rect 20269 25789 20303 25823
rect 20303 25789 20312 25823
rect 20260 25780 20312 25789
rect 7104 25712 7156 25764
rect 8576 25712 8628 25764
rect 15108 25712 15160 25764
rect 11980 25644 12032 25696
rect 12716 25644 12768 25696
rect 14832 25644 14884 25696
rect 15476 25644 15528 25696
rect 15844 25644 15896 25696
rect 16396 25644 16448 25696
rect 17868 25712 17920 25764
rect 18328 25712 18380 25764
rect 21364 25891 21416 25900
rect 21364 25857 21373 25891
rect 21373 25857 21407 25891
rect 21407 25857 21416 25891
rect 21364 25848 21416 25857
rect 22008 25891 22060 25900
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 22560 25891 22612 25900
rect 22560 25857 22593 25891
rect 22593 25857 22612 25891
rect 22560 25848 22612 25857
rect 22284 25712 22336 25764
rect 21640 25644 21692 25696
rect 22008 25644 22060 25696
rect 24860 25984 24912 26036
rect 29460 25984 29512 26036
rect 29644 25984 29696 26036
rect 31668 25984 31720 26036
rect 32680 25984 32732 26036
rect 32772 25984 32824 26036
rect 33784 25984 33836 26036
rect 36268 25984 36320 26036
rect 39028 26027 39080 26036
rect 39028 25993 39037 26027
rect 39037 25993 39071 26027
rect 39071 25993 39080 26027
rect 39028 25984 39080 25993
rect 25228 25916 25280 25968
rect 23848 25891 23900 25900
rect 23848 25857 23857 25891
rect 23857 25857 23891 25891
rect 23891 25857 23900 25891
rect 23848 25848 23900 25857
rect 24952 25848 25004 25900
rect 25504 25848 25556 25900
rect 23664 25780 23716 25832
rect 27620 25823 27672 25832
rect 27620 25789 27629 25823
rect 27629 25789 27663 25823
rect 27663 25789 27672 25823
rect 27620 25780 27672 25789
rect 27896 25823 27948 25832
rect 27896 25789 27905 25823
rect 27905 25789 27939 25823
rect 27939 25789 27948 25823
rect 27896 25780 27948 25789
rect 28448 25780 28500 25832
rect 31392 25916 31444 25968
rect 37556 25959 37608 25968
rect 37556 25925 37565 25959
rect 37565 25925 37599 25959
rect 37599 25925 37608 25959
rect 37556 25916 37608 25925
rect 39120 25916 39172 25968
rect 39304 25959 39356 25968
rect 39304 25925 39313 25959
rect 39313 25925 39347 25959
rect 39347 25925 39356 25959
rect 39304 25916 39356 25925
rect 40040 25984 40092 26036
rect 40316 25984 40368 26036
rect 40592 25984 40644 26036
rect 42064 26027 42116 26036
rect 42064 25993 42073 26027
rect 42073 25993 42107 26027
rect 42107 25993 42116 26027
rect 42064 25984 42116 25993
rect 40776 25959 40828 25968
rect 39212 25848 39264 25900
rect 40040 25891 40092 25900
rect 40040 25857 40049 25891
rect 40049 25857 40083 25891
rect 40083 25857 40092 25891
rect 40040 25848 40092 25857
rect 40132 25891 40184 25900
rect 40132 25857 40141 25891
rect 40141 25857 40175 25891
rect 40175 25857 40184 25891
rect 40132 25848 40184 25857
rect 40224 25891 40276 25900
rect 40224 25857 40233 25891
rect 40233 25857 40267 25891
rect 40267 25857 40276 25891
rect 40224 25848 40276 25857
rect 40500 25848 40552 25900
rect 40776 25925 40789 25959
rect 40789 25925 40823 25959
rect 40823 25925 40828 25959
rect 40776 25916 40828 25925
rect 40868 25891 40920 25900
rect 40868 25857 40877 25891
rect 40877 25857 40911 25891
rect 40911 25857 40920 25891
rect 40868 25848 40920 25857
rect 41052 25891 41104 25900
rect 41052 25857 41061 25891
rect 41061 25857 41095 25891
rect 41095 25857 41104 25891
rect 41052 25848 41104 25857
rect 41880 25891 41932 25900
rect 41880 25857 41889 25891
rect 41889 25857 41923 25891
rect 41923 25857 41932 25891
rect 41880 25848 41932 25857
rect 32128 25780 32180 25832
rect 37280 25823 37332 25832
rect 37280 25789 37289 25823
rect 37289 25789 37323 25823
rect 37323 25789 37332 25823
rect 37280 25780 37332 25789
rect 39396 25780 39448 25832
rect 40776 25780 40828 25832
rect 23296 25712 23348 25764
rect 23020 25687 23072 25696
rect 23020 25653 23029 25687
rect 23029 25653 23063 25687
rect 23063 25653 23072 25687
rect 23020 25644 23072 25653
rect 23756 25687 23808 25696
rect 23756 25653 23765 25687
rect 23765 25653 23799 25687
rect 23799 25653 23808 25687
rect 23756 25644 23808 25653
rect 25044 25644 25096 25696
rect 28908 25644 28960 25696
rect 30564 25644 30616 25696
rect 32864 25687 32916 25696
rect 32864 25653 32873 25687
rect 32873 25653 32907 25687
rect 32907 25653 32916 25687
rect 32864 25644 32916 25653
rect 33784 25644 33836 25696
rect 39120 25687 39172 25696
rect 39120 25653 39129 25687
rect 39129 25653 39163 25687
rect 39163 25653 39172 25687
rect 39120 25644 39172 25653
rect 40224 25712 40276 25764
rect 40868 25712 40920 25764
rect 40960 25644 41012 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 14832 25440 14884 25492
rect 14924 25440 14976 25492
rect 4436 25372 4488 25424
rect 5448 25372 5500 25424
rect 5816 25372 5868 25424
rect 17776 25440 17828 25492
rect 18144 25483 18196 25492
rect 18144 25449 18153 25483
rect 18153 25449 18187 25483
rect 18187 25449 18196 25483
rect 18144 25440 18196 25449
rect 21180 25440 21232 25492
rect 22100 25440 22152 25492
rect 23388 25440 23440 25492
rect 24952 25483 25004 25492
rect 24952 25449 24961 25483
rect 24961 25449 24995 25483
rect 24995 25449 25004 25483
rect 24952 25440 25004 25449
rect 2872 25347 2924 25356
rect 2872 25313 2881 25347
rect 2881 25313 2915 25347
rect 2915 25313 2924 25347
rect 2872 25304 2924 25313
rect 3516 25304 3568 25356
rect 6092 25304 6144 25356
rect 15108 25347 15160 25356
rect 15108 25313 15117 25347
rect 15117 25313 15151 25347
rect 15151 25313 15160 25347
rect 15108 25304 15160 25313
rect 4528 25236 4580 25288
rect 7564 25236 7616 25288
rect 2964 25168 3016 25220
rect 7748 25236 7800 25288
rect 13452 25279 13504 25288
rect 13452 25245 13461 25279
rect 13461 25245 13495 25279
rect 13495 25245 13504 25279
rect 13452 25236 13504 25245
rect 15016 25279 15068 25288
rect 15016 25245 15025 25279
rect 15025 25245 15059 25279
rect 15059 25245 15068 25279
rect 15016 25236 15068 25245
rect 20812 25372 20864 25424
rect 15844 25347 15896 25356
rect 15844 25313 15853 25347
rect 15853 25313 15887 25347
rect 15887 25313 15896 25347
rect 15844 25304 15896 25313
rect 8300 25168 8352 25220
rect 11428 25168 11480 25220
rect 14372 25211 14424 25220
rect 14372 25177 14381 25211
rect 14381 25177 14415 25211
rect 14415 25177 14424 25211
rect 14372 25168 14424 25177
rect 14556 25211 14608 25220
rect 14556 25177 14565 25211
rect 14565 25177 14599 25211
rect 14599 25177 14608 25211
rect 14556 25168 14608 25177
rect 1400 25143 1452 25152
rect 1400 25109 1409 25143
rect 1409 25109 1443 25143
rect 1443 25109 1452 25143
rect 1400 25100 1452 25109
rect 5724 25100 5776 25152
rect 6460 25100 6512 25152
rect 7840 25143 7892 25152
rect 7840 25109 7849 25143
rect 7849 25109 7883 25143
rect 7883 25109 7892 25143
rect 7840 25100 7892 25109
rect 13636 25100 13688 25152
rect 14924 25100 14976 25152
rect 15568 25279 15620 25288
rect 15568 25245 15577 25279
rect 15577 25245 15611 25279
rect 15611 25245 15620 25279
rect 15568 25236 15620 25245
rect 18328 25304 18380 25356
rect 18236 25279 18288 25288
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 20904 25236 20956 25288
rect 21088 25236 21140 25288
rect 21640 25279 21692 25288
rect 21640 25245 21649 25279
rect 21649 25245 21683 25279
rect 21683 25245 21692 25279
rect 21640 25236 21692 25245
rect 23020 25304 23072 25356
rect 17132 25168 17184 25220
rect 17868 25211 17920 25220
rect 17868 25177 17877 25211
rect 17877 25177 17911 25211
rect 17911 25177 17920 25211
rect 17868 25168 17920 25177
rect 17960 25168 18012 25220
rect 22100 25236 22152 25288
rect 22284 25279 22336 25288
rect 22284 25245 22293 25279
rect 22293 25245 22327 25279
rect 22327 25245 22336 25279
rect 23572 25304 23624 25356
rect 22284 25236 22336 25245
rect 16764 25100 16816 25152
rect 18420 25143 18472 25152
rect 18420 25109 18429 25143
rect 18429 25109 18463 25143
rect 18463 25109 18472 25143
rect 18420 25100 18472 25109
rect 20444 25100 20496 25152
rect 22100 25143 22152 25152
rect 22100 25109 22109 25143
rect 22109 25109 22143 25143
rect 22143 25109 22152 25143
rect 22100 25100 22152 25109
rect 22284 25100 22336 25152
rect 23020 25143 23072 25152
rect 23020 25109 23029 25143
rect 23029 25109 23063 25143
rect 23063 25109 23072 25143
rect 23020 25100 23072 25109
rect 23296 25279 23348 25288
rect 23296 25245 23305 25279
rect 23305 25245 23339 25279
rect 23339 25245 23348 25279
rect 23296 25236 23348 25245
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 23940 25236 23992 25288
rect 24584 25236 24636 25288
rect 26240 25440 26292 25492
rect 27896 25440 27948 25492
rect 25504 25372 25556 25424
rect 26700 25372 26752 25424
rect 29276 25372 29328 25424
rect 25412 25236 25464 25288
rect 28908 25304 28960 25356
rect 29092 25304 29144 25356
rect 30472 25372 30524 25424
rect 26976 25279 27028 25288
rect 26976 25245 26985 25279
rect 26985 25245 27019 25279
rect 27019 25245 27028 25279
rect 26976 25236 27028 25245
rect 27160 25279 27212 25288
rect 27160 25245 27169 25279
rect 27169 25245 27203 25279
rect 27203 25245 27212 25279
rect 27160 25236 27212 25245
rect 30288 25279 30340 25288
rect 30288 25245 30297 25279
rect 30297 25245 30331 25279
rect 30331 25245 30340 25279
rect 30288 25236 30340 25245
rect 30748 25236 30800 25288
rect 30932 25236 30984 25288
rect 34520 25347 34572 25356
rect 34520 25313 34529 25347
rect 34529 25313 34563 25347
rect 34563 25313 34572 25347
rect 34520 25304 34572 25313
rect 34796 25304 34848 25356
rect 32588 25236 32640 25288
rect 35256 25236 35308 25288
rect 36176 25304 36228 25356
rect 36452 25304 36504 25356
rect 35992 25279 36044 25288
rect 35992 25245 36001 25279
rect 36001 25245 36035 25279
rect 36035 25245 36044 25279
rect 35992 25236 36044 25245
rect 36544 25236 36596 25288
rect 37280 25372 37332 25424
rect 23388 25211 23440 25220
rect 23388 25177 23397 25211
rect 23397 25177 23431 25211
rect 23431 25177 23440 25211
rect 23388 25168 23440 25177
rect 23572 25168 23624 25220
rect 25320 25211 25372 25220
rect 25320 25177 25329 25211
rect 25329 25177 25363 25211
rect 25363 25177 25372 25211
rect 25320 25168 25372 25177
rect 25872 25168 25924 25220
rect 32496 25211 32548 25220
rect 32496 25177 32505 25211
rect 32505 25177 32539 25211
rect 32539 25177 32548 25211
rect 32496 25168 32548 25177
rect 33784 25168 33836 25220
rect 34244 25211 34296 25220
rect 34244 25177 34253 25211
rect 34253 25177 34287 25211
rect 34287 25177 34296 25211
rect 34244 25168 34296 25177
rect 34520 25168 34572 25220
rect 27436 25100 27488 25152
rect 28540 25143 28592 25152
rect 28540 25109 28549 25143
rect 28549 25109 28583 25143
rect 28583 25109 28592 25143
rect 28540 25100 28592 25109
rect 28632 25143 28684 25152
rect 28632 25109 28641 25143
rect 28641 25109 28675 25143
rect 28675 25109 28684 25143
rect 28632 25100 28684 25109
rect 29092 25100 29144 25152
rect 29736 25143 29788 25152
rect 29736 25109 29745 25143
rect 29745 25109 29779 25143
rect 29779 25109 29788 25143
rect 29736 25100 29788 25109
rect 30656 25143 30708 25152
rect 30656 25109 30665 25143
rect 30665 25109 30699 25143
rect 30699 25109 30708 25143
rect 30656 25100 30708 25109
rect 30840 25100 30892 25152
rect 31576 25100 31628 25152
rect 35348 25100 35400 25152
rect 35900 25211 35952 25220
rect 35900 25177 35909 25211
rect 35909 25177 35943 25211
rect 35943 25177 35952 25211
rect 35900 25168 35952 25177
rect 36268 25168 36320 25220
rect 38568 25100 38620 25152
rect 41788 25440 41840 25492
rect 40592 25236 40644 25288
rect 40500 25211 40552 25220
rect 40500 25177 40509 25211
rect 40509 25177 40543 25211
rect 40543 25177 40552 25211
rect 40500 25168 40552 25177
rect 40960 25168 41012 25220
rect 40776 25100 40828 25152
rect 41512 25143 41564 25152
rect 41512 25109 41521 25143
rect 41521 25109 41555 25143
rect 41555 25109 41564 25143
rect 41512 25100 41564 25109
rect 41604 25100 41656 25152
rect 41972 25168 42024 25220
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 2688 24760 2740 24812
rect 4712 24896 4764 24948
rect 7288 24896 7340 24948
rect 7932 24896 7984 24948
rect 8116 24896 8168 24948
rect 8392 24896 8444 24948
rect 13636 24896 13688 24948
rect 16120 24896 16172 24948
rect 17224 24896 17276 24948
rect 3884 24803 3936 24812
rect 3884 24769 3893 24803
rect 3893 24769 3927 24803
rect 3927 24769 3936 24803
rect 3884 24760 3936 24769
rect 4436 24803 4488 24812
rect 4436 24769 4445 24803
rect 4445 24769 4479 24803
rect 4479 24769 4488 24803
rect 4436 24760 4488 24769
rect 4528 24803 4580 24812
rect 4528 24769 4537 24803
rect 4537 24769 4571 24803
rect 4571 24769 4580 24803
rect 4528 24760 4580 24769
rect 4620 24803 4672 24812
rect 4620 24769 4629 24803
rect 4629 24769 4663 24803
rect 4663 24769 4672 24803
rect 4620 24760 4672 24769
rect 1308 24624 1360 24676
rect 2504 24556 2556 24608
rect 3976 24556 4028 24608
rect 5356 24828 5408 24880
rect 7380 24828 7432 24880
rect 5080 24803 5132 24812
rect 5080 24769 5089 24803
rect 5089 24769 5123 24803
rect 5123 24769 5132 24803
rect 5080 24760 5132 24769
rect 5264 24803 5316 24812
rect 5264 24769 5273 24803
rect 5273 24769 5307 24803
rect 5307 24769 5316 24803
rect 5264 24760 5316 24769
rect 6184 24760 6236 24812
rect 6092 24735 6144 24744
rect 6092 24701 6101 24735
rect 6101 24701 6135 24735
rect 6135 24701 6144 24735
rect 6092 24692 6144 24701
rect 6920 24760 6972 24812
rect 7104 24735 7156 24744
rect 7104 24701 7113 24735
rect 7113 24701 7147 24735
rect 7147 24701 7156 24735
rect 7104 24692 7156 24701
rect 7472 24735 7524 24744
rect 7472 24701 7481 24735
rect 7481 24701 7515 24735
rect 7515 24701 7524 24735
rect 7472 24692 7524 24701
rect 7564 24692 7616 24744
rect 8208 24760 8260 24812
rect 8300 24760 8352 24812
rect 9036 24803 9088 24812
rect 9036 24769 9045 24803
rect 9045 24769 9079 24803
rect 9079 24769 9088 24803
rect 9036 24760 9088 24769
rect 9220 24803 9272 24812
rect 9220 24769 9229 24803
rect 9229 24769 9263 24803
rect 9263 24769 9272 24803
rect 9220 24760 9272 24769
rect 9588 24828 9640 24880
rect 9496 24760 9548 24812
rect 6828 24624 6880 24676
rect 7748 24624 7800 24676
rect 8392 24735 8444 24744
rect 8392 24701 8401 24735
rect 8401 24701 8435 24735
rect 8435 24701 8444 24735
rect 8392 24692 8444 24701
rect 8852 24692 8904 24744
rect 10324 24692 10376 24744
rect 11336 24692 11388 24744
rect 12072 24735 12124 24744
rect 12072 24701 12081 24735
rect 12081 24701 12115 24735
rect 12115 24701 12124 24735
rect 12072 24692 12124 24701
rect 12716 24803 12768 24812
rect 12716 24769 12725 24803
rect 12725 24769 12759 24803
rect 12759 24769 12768 24803
rect 12716 24760 12768 24769
rect 13820 24760 13872 24812
rect 14372 24803 14424 24812
rect 14372 24769 14381 24803
rect 14381 24769 14415 24803
rect 14415 24769 14424 24803
rect 14372 24760 14424 24769
rect 15016 24828 15068 24880
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 14924 24803 14976 24812
rect 14924 24769 14933 24803
rect 14933 24769 14967 24803
rect 14967 24769 14976 24803
rect 14924 24760 14976 24769
rect 15660 24803 15712 24812
rect 15660 24769 15669 24803
rect 15669 24769 15703 24803
rect 15703 24769 15712 24803
rect 15660 24760 15712 24769
rect 17592 24828 17644 24880
rect 15936 24803 15988 24812
rect 15936 24769 15945 24803
rect 15945 24769 15979 24803
rect 15979 24769 15988 24803
rect 15936 24760 15988 24769
rect 18420 24760 18472 24812
rect 19340 24896 19392 24948
rect 19616 24896 19668 24948
rect 21364 24896 21416 24948
rect 22192 24939 22244 24948
rect 22192 24905 22201 24939
rect 22201 24905 22235 24939
rect 22235 24905 22244 24939
rect 22192 24896 22244 24905
rect 22376 24896 22428 24948
rect 25320 24896 25372 24948
rect 21272 24828 21324 24880
rect 9588 24624 9640 24676
rect 12808 24624 12860 24676
rect 7012 24556 7064 24608
rect 7196 24556 7248 24608
rect 7932 24556 7984 24608
rect 10232 24599 10284 24608
rect 10232 24565 10241 24599
rect 10241 24565 10275 24599
rect 10275 24565 10284 24599
rect 10232 24556 10284 24565
rect 12532 24599 12584 24608
rect 12532 24565 12541 24599
rect 12541 24565 12575 24599
rect 12575 24565 12584 24599
rect 12532 24556 12584 24565
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 13084 24599 13136 24608
rect 13084 24565 13093 24599
rect 13093 24565 13127 24599
rect 13127 24565 13136 24599
rect 13084 24556 13136 24565
rect 13176 24599 13228 24608
rect 13176 24565 13185 24599
rect 13185 24565 13219 24599
rect 13219 24565 13228 24599
rect 13176 24556 13228 24565
rect 18144 24735 18196 24744
rect 18144 24701 18153 24735
rect 18153 24701 18187 24735
rect 18187 24701 18196 24735
rect 18144 24692 18196 24701
rect 19524 24692 19576 24744
rect 15476 24624 15528 24676
rect 15660 24624 15712 24676
rect 20168 24760 20220 24812
rect 22284 24803 22336 24812
rect 22284 24769 22293 24803
rect 22293 24769 22327 24803
rect 22327 24769 22336 24803
rect 22284 24760 22336 24769
rect 23112 24760 23164 24812
rect 23388 24828 23440 24880
rect 25688 24871 25740 24880
rect 25688 24837 25697 24871
rect 25697 24837 25731 24871
rect 25731 24837 25740 24871
rect 25688 24828 25740 24837
rect 25872 24871 25924 24880
rect 24676 24760 24728 24812
rect 25228 24760 25280 24812
rect 25872 24837 25897 24871
rect 25897 24837 25924 24871
rect 25872 24828 25924 24837
rect 26056 24828 26108 24880
rect 26332 24803 26384 24812
rect 25044 24735 25096 24744
rect 25044 24701 25053 24735
rect 25053 24701 25087 24735
rect 25087 24701 25096 24735
rect 25044 24692 25096 24701
rect 25504 24735 25556 24744
rect 25504 24701 25513 24735
rect 25513 24701 25547 24735
rect 25547 24701 25556 24735
rect 25504 24692 25556 24701
rect 18328 24624 18380 24676
rect 20076 24624 20128 24676
rect 22744 24667 22796 24676
rect 22744 24633 22753 24667
rect 22753 24633 22787 24667
rect 22787 24633 22796 24667
rect 22744 24624 22796 24633
rect 24860 24667 24912 24676
rect 24860 24633 24869 24667
rect 24869 24633 24903 24667
rect 24903 24633 24912 24667
rect 24860 24624 24912 24633
rect 14004 24599 14056 24608
rect 14004 24565 14013 24599
rect 14013 24565 14047 24599
rect 14047 24565 14056 24599
rect 14004 24556 14056 24565
rect 14188 24599 14240 24608
rect 14188 24565 14197 24599
rect 14197 24565 14231 24599
rect 14231 24565 14240 24599
rect 14188 24556 14240 24565
rect 15384 24556 15436 24608
rect 15936 24556 15988 24608
rect 17040 24599 17092 24608
rect 17040 24565 17049 24599
rect 17049 24565 17083 24599
rect 17083 24565 17092 24599
rect 17040 24556 17092 24565
rect 18604 24599 18656 24608
rect 18604 24565 18613 24599
rect 18613 24565 18647 24599
rect 18647 24565 18656 24599
rect 18604 24556 18656 24565
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 25320 24556 25372 24608
rect 25688 24692 25740 24744
rect 26332 24769 26341 24803
rect 26341 24769 26375 24803
rect 26375 24769 26384 24803
rect 26332 24760 26384 24769
rect 28632 24896 28684 24948
rect 27436 24871 27488 24880
rect 27436 24837 27445 24871
rect 27445 24837 27479 24871
rect 27479 24837 27488 24871
rect 27436 24828 27488 24837
rect 27804 24828 27856 24880
rect 27528 24803 27580 24812
rect 27528 24769 27537 24803
rect 27537 24769 27571 24803
rect 27571 24769 27580 24803
rect 27528 24760 27580 24769
rect 27712 24760 27764 24812
rect 28816 24828 28868 24880
rect 27988 24803 28040 24812
rect 27988 24769 27997 24803
rect 27997 24769 28031 24803
rect 28031 24769 28040 24803
rect 27988 24760 28040 24769
rect 26516 24692 26568 24744
rect 28632 24803 28684 24812
rect 28632 24769 28641 24803
rect 28641 24769 28675 24803
rect 28675 24769 28684 24803
rect 28632 24760 28684 24769
rect 30288 24896 30340 24948
rect 31852 24939 31904 24948
rect 31852 24905 31861 24939
rect 31861 24905 31895 24939
rect 31895 24905 31904 24939
rect 31852 24896 31904 24905
rect 32680 24896 32732 24948
rect 33048 24896 33100 24948
rect 34244 24896 34296 24948
rect 35256 24896 35308 24948
rect 26056 24599 26108 24608
rect 26056 24565 26065 24599
rect 26065 24565 26099 24599
rect 26099 24565 26108 24599
rect 26056 24556 26108 24565
rect 26240 24624 26292 24676
rect 26700 24556 26752 24608
rect 27160 24624 27212 24676
rect 27252 24624 27304 24676
rect 28172 24667 28224 24676
rect 28172 24633 28181 24667
rect 28181 24633 28215 24667
rect 28215 24633 28224 24667
rect 28172 24624 28224 24633
rect 27712 24556 27764 24608
rect 27804 24599 27856 24608
rect 27804 24565 27813 24599
rect 27813 24565 27847 24599
rect 27847 24565 27856 24599
rect 27804 24556 27856 24565
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 29276 24760 29328 24812
rect 29644 24871 29696 24880
rect 29644 24837 29653 24871
rect 29653 24837 29687 24871
rect 29687 24837 29696 24871
rect 29644 24828 29696 24837
rect 31392 24828 31444 24880
rect 32588 24828 32640 24880
rect 40500 24896 40552 24948
rect 40868 24896 40920 24948
rect 29828 24803 29880 24812
rect 29828 24769 29837 24803
rect 29837 24769 29871 24803
rect 29871 24769 29880 24803
rect 29828 24760 29880 24769
rect 29552 24692 29604 24744
rect 28908 24624 28960 24676
rect 30380 24735 30432 24744
rect 30380 24701 30389 24735
rect 30389 24701 30423 24735
rect 30423 24701 30432 24735
rect 30380 24692 30432 24701
rect 32588 24692 32640 24744
rect 32772 24803 32824 24812
rect 32772 24769 32782 24803
rect 32782 24769 32816 24803
rect 32816 24769 32824 24803
rect 32772 24760 32824 24769
rect 32956 24803 33008 24812
rect 32956 24769 32965 24803
rect 32965 24769 32999 24803
rect 32999 24769 33008 24803
rect 32956 24760 33008 24769
rect 33692 24803 33744 24812
rect 33692 24769 33701 24803
rect 33701 24769 33735 24803
rect 33735 24769 33744 24803
rect 33692 24760 33744 24769
rect 35164 24760 35216 24812
rect 35348 24803 35400 24812
rect 35348 24769 35357 24803
rect 35357 24769 35391 24803
rect 35391 24769 35400 24803
rect 35348 24760 35400 24769
rect 35624 24803 35676 24812
rect 35440 24769 35449 24802
rect 35449 24769 35483 24802
rect 35483 24769 35492 24802
rect 35440 24750 35492 24769
rect 35624 24769 35641 24803
rect 35641 24769 35676 24803
rect 35624 24760 35676 24769
rect 36268 24828 36320 24880
rect 36544 24828 36596 24880
rect 29828 24556 29880 24608
rect 30932 24556 30984 24608
rect 33140 24624 33192 24676
rect 31484 24556 31536 24608
rect 34520 24692 34572 24744
rect 33692 24624 33744 24676
rect 36176 24692 36228 24744
rect 36452 24735 36504 24744
rect 36452 24701 36461 24735
rect 36461 24701 36495 24735
rect 36495 24701 36504 24735
rect 36452 24692 36504 24701
rect 36636 24624 36688 24676
rect 37004 24828 37056 24880
rect 37280 24828 37332 24880
rect 39120 24871 39172 24880
rect 39120 24837 39129 24871
rect 39129 24837 39163 24871
rect 39163 24837 39172 24871
rect 39120 24828 39172 24837
rect 39580 24828 39632 24880
rect 41696 24828 41748 24880
rect 41788 24828 41840 24880
rect 38752 24760 38804 24812
rect 40868 24803 40920 24812
rect 40868 24769 40877 24803
rect 40877 24769 40911 24803
rect 40911 24769 40920 24803
rect 40868 24760 40920 24769
rect 40960 24803 41012 24812
rect 40960 24769 40969 24803
rect 40969 24769 41003 24803
rect 41003 24769 41012 24803
rect 40960 24760 41012 24769
rect 41328 24803 41380 24812
rect 41328 24769 41337 24803
rect 41337 24769 41371 24803
rect 41371 24769 41380 24803
rect 41328 24760 41380 24769
rect 39580 24692 39632 24744
rect 38752 24624 38804 24676
rect 40592 24735 40644 24744
rect 40592 24701 40601 24735
rect 40601 24701 40635 24735
rect 40635 24701 40644 24735
rect 40592 24692 40644 24701
rect 41788 24667 41840 24676
rect 41788 24633 41797 24667
rect 41797 24633 41831 24667
rect 41831 24633 41840 24667
rect 41788 24624 41840 24633
rect 33508 24599 33560 24608
rect 33508 24565 33517 24599
rect 33517 24565 33551 24599
rect 33551 24565 33560 24599
rect 33508 24556 33560 24565
rect 35624 24556 35676 24608
rect 37280 24556 37332 24608
rect 38660 24556 38712 24608
rect 39672 24556 39724 24608
rect 41420 24556 41472 24608
rect 41512 24599 41564 24608
rect 41512 24565 41521 24599
rect 41521 24565 41555 24599
rect 41555 24565 41564 24599
rect 41512 24556 41564 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3516 24216 3568 24268
rect 2964 24148 3016 24200
rect 3792 24148 3844 24200
rect 6552 24352 6604 24404
rect 7288 24352 7340 24404
rect 8024 24395 8076 24404
rect 8024 24361 8033 24395
rect 8033 24361 8067 24395
rect 8067 24361 8076 24395
rect 8024 24352 8076 24361
rect 8392 24352 8444 24404
rect 9312 24352 9364 24404
rect 11336 24395 11388 24404
rect 11336 24361 11345 24395
rect 11345 24361 11379 24395
rect 11379 24361 11388 24395
rect 11336 24352 11388 24361
rect 12992 24352 13044 24404
rect 2136 24080 2188 24132
rect 4252 24080 4304 24132
rect 4804 24148 4856 24200
rect 5172 24191 5224 24200
rect 5172 24157 5181 24191
rect 5181 24157 5215 24191
rect 5215 24157 5224 24191
rect 5172 24148 5224 24157
rect 7380 24284 7432 24336
rect 8208 24284 8260 24336
rect 6184 24216 6236 24268
rect 6092 24191 6144 24200
rect 6092 24157 6101 24191
rect 6101 24157 6135 24191
rect 6135 24157 6144 24191
rect 6092 24148 6144 24157
rect 6460 24148 6512 24200
rect 7564 24259 7616 24268
rect 7564 24225 7573 24259
rect 7573 24225 7607 24259
rect 7607 24225 7616 24259
rect 7564 24216 7616 24225
rect 7656 24216 7708 24268
rect 14740 24352 14792 24404
rect 14004 24284 14056 24336
rect 14096 24216 14148 24268
rect 6828 24191 6880 24200
rect 6828 24157 6837 24191
rect 6837 24157 6871 24191
rect 6871 24157 6880 24191
rect 6828 24148 6880 24157
rect 4620 24080 4672 24132
rect 5632 24080 5684 24132
rect 7104 24191 7156 24200
rect 7104 24157 7113 24191
rect 7113 24157 7147 24191
rect 7147 24157 7156 24191
rect 7104 24148 7156 24157
rect 7472 24148 7524 24200
rect 8208 24148 8260 24200
rect 7748 24080 7800 24132
rect 7840 24123 7892 24132
rect 7840 24089 7865 24123
rect 7865 24089 7892 24123
rect 7840 24080 7892 24089
rect 8024 24080 8076 24132
rect 8944 24148 8996 24200
rect 9220 24191 9272 24200
rect 9220 24157 9229 24191
rect 9229 24157 9263 24191
rect 9263 24157 9272 24191
rect 9220 24148 9272 24157
rect 9312 24191 9364 24200
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 9496 24191 9548 24200
rect 9496 24157 9505 24191
rect 9505 24157 9539 24191
rect 9539 24157 9548 24191
rect 9496 24148 9548 24157
rect 9588 24191 9640 24200
rect 9588 24157 9597 24191
rect 9597 24157 9631 24191
rect 9631 24157 9640 24191
rect 9588 24148 9640 24157
rect 9128 24080 9180 24132
rect 9956 24191 10008 24200
rect 9956 24157 9965 24191
rect 9965 24157 9999 24191
rect 9999 24157 10008 24191
rect 9956 24148 10008 24157
rect 11796 24191 11848 24200
rect 11796 24157 11805 24191
rect 11805 24157 11839 24191
rect 11839 24157 11848 24191
rect 11796 24148 11848 24157
rect 12532 24148 12584 24200
rect 2780 24012 2832 24064
rect 4160 24012 4212 24064
rect 4712 24012 4764 24064
rect 5080 24012 5132 24064
rect 5448 24012 5500 24064
rect 6920 24012 6972 24064
rect 7104 24012 7156 24064
rect 7564 24012 7616 24064
rect 9404 24012 9456 24064
rect 14832 24148 14884 24200
rect 17960 24352 18012 24404
rect 19156 24352 19208 24404
rect 19892 24352 19944 24404
rect 20720 24352 20772 24404
rect 22192 24352 22244 24404
rect 26976 24352 27028 24404
rect 27896 24352 27948 24404
rect 28356 24352 28408 24404
rect 28816 24352 28868 24404
rect 18328 24284 18380 24336
rect 17040 24216 17092 24268
rect 18144 24216 18196 24268
rect 18604 24216 18656 24268
rect 16948 24148 17000 24200
rect 17224 24191 17276 24200
rect 17224 24157 17233 24191
rect 17233 24157 17267 24191
rect 17267 24157 17276 24191
rect 17224 24148 17276 24157
rect 18512 24148 18564 24200
rect 19524 24216 19576 24268
rect 18788 24148 18840 24200
rect 16672 24080 16724 24132
rect 18236 24123 18288 24132
rect 18236 24089 18245 24123
rect 18245 24089 18279 24123
rect 18279 24089 18288 24123
rect 19064 24148 19116 24200
rect 19432 24191 19484 24200
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 19708 24191 19760 24200
rect 19708 24157 19717 24191
rect 19717 24157 19751 24191
rect 19751 24157 19760 24191
rect 19708 24148 19760 24157
rect 24216 24284 24268 24336
rect 25136 24284 25188 24336
rect 28632 24284 28684 24336
rect 29644 24284 29696 24336
rect 30380 24352 30432 24404
rect 30564 24352 30616 24404
rect 30840 24352 30892 24404
rect 31668 24352 31720 24404
rect 32956 24395 33008 24404
rect 32956 24361 32965 24395
rect 32965 24361 32999 24395
rect 32999 24361 33008 24395
rect 32956 24352 33008 24361
rect 33140 24352 33192 24404
rect 33600 24352 33652 24404
rect 34612 24352 34664 24404
rect 38660 24352 38712 24404
rect 41328 24352 41380 24404
rect 19984 24216 20036 24268
rect 21824 24259 21876 24268
rect 21824 24225 21833 24259
rect 21833 24225 21867 24259
rect 21867 24225 21876 24259
rect 21824 24216 21876 24225
rect 23480 24216 23532 24268
rect 24676 24216 24728 24268
rect 25780 24259 25832 24268
rect 25780 24225 25789 24259
rect 25789 24225 25823 24259
rect 25823 24225 25832 24259
rect 25780 24216 25832 24225
rect 18236 24080 18288 24089
rect 16396 24012 16448 24064
rect 16764 24012 16816 24064
rect 18420 24055 18472 24064
rect 18420 24021 18429 24055
rect 18429 24021 18463 24055
rect 18463 24021 18472 24055
rect 18420 24012 18472 24021
rect 18788 24012 18840 24064
rect 19156 24012 19208 24064
rect 19340 24055 19392 24064
rect 19340 24021 19349 24055
rect 19349 24021 19383 24055
rect 19383 24021 19392 24055
rect 19340 24012 19392 24021
rect 19524 24055 19576 24064
rect 19524 24021 19533 24055
rect 19533 24021 19567 24055
rect 19567 24021 19576 24055
rect 19524 24012 19576 24021
rect 19892 24123 19944 24132
rect 19892 24089 19901 24123
rect 19901 24089 19935 24123
rect 19935 24089 19944 24123
rect 19892 24080 19944 24089
rect 24584 24191 24636 24200
rect 24584 24157 24593 24191
rect 24593 24157 24627 24191
rect 24627 24157 24636 24191
rect 24584 24148 24636 24157
rect 24860 24191 24912 24200
rect 24860 24157 24869 24191
rect 24869 24157 24903 24191
rect 24903 24157 24912 24191
rect 24860 24148 24912 24157
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 25136 24191 25188 24200
rect 25136 24157 25145 24191
rect 25145 24157 25179 24191
rect 25179 24157 25188 24191
rect 25136 24148 25188 24157
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 25688 24148 25740 24200
rect 26056 24148 26108 24200
rect 26240 24191 26292 24200
rect 26240 24157 26249 24191
rect 26249 24157 26283 24191
rect 26283 24157 26292 24191
rect 26240 24148 26292 24157
rect 20444 24080 20496 24132
rect 21916 24080 21968 24132
rect 22468 24123 22520 24132
rect 22468 24089 22477 24123
rect 22477 24089 22511 24123
rect 22511 24089 22520 24123
rect 22468 24080 22520 24089
rect 25596 24080 25648 24132
rect 26148 24123 26200 24132
rect 26148 24089 26157 24123
rect 26157 24089 26191 24123
rect 26191 24089 26200 24123
rect 26148 24080 26200 24089
rect 20260 24012 20312 24064
rect 24584 24012 24636 24064
rect 26516 24191 26568 24200
rect 26516 24157 26525 24191
rect 26525 24157 26559 24191
rect 26559 24157 26568 24191
rect 26516 24148 26568 24157
rect 27620 24216 27672 24268
rect 28172 24216 28224 24268
rect 33508 24284 33560 24336
rect 26792 24191 26844 24200
rect 26792 24157 26801 24191
rect 26801 24157 26835 24191
rect 26835 24157 26844 24191
rect 26792 24148 26844 24157
rect 28448 24148 28500 24200
rect 27160 24123 27212 24132
rect 27160 24089 27169 24123
rect 27169 24089 27203 24123
rect 27203 24089 27212 24123
rect 27160 24080 27212 24089
rect 28816 24012 28868 24064
rect 29828 24080 29880 24132
rect 30472 24191 30524 24200
rect 30472 24157 30481 24191
rect 30481 24157 30515 24191
rect 30515 24157 30524 24191
rect 30472 24148 30524 24157
rect 30656 24148 30708 24200
rect 30840 24191 30892 24200
rect 30840 24157 30849 24191
rect 30849 24157 30883 24191
rect 30883 24157 30892 24191
rect 30840 24148 30892 24157
rect 31208 24148 31260 24200
rect 31392 24148 31444 24200
rect 31852 24148 31904 24200
rect 30932 24080 30984 24132
rect 31024 24080 31076 24132
rect 30840 24012 30892 24064
rect 31668 24080 31720 24132
rect 32956 24216 33008 24268
rect 33048 24216 33100 24268
rect 35900 24259 35952 24268
rect 35900 24225 35909 24259
rect 35909 24225 35943 24259
rect 35943 24225 35952 24259
rect 35900 24216 35952 24225
rect 35992 24216 36044 24268
rect 36452 24284 36504 24336
rect 37004 24259 37056 24268
rect 37004 24225 37013 24259
rect 37013 24225 37047 24259
rect 37047 24225 37056 24259
rect 37004 24216 37056 24225
rect 37280 24259 37332 24268
rect 37280 24225 37289 24259
rect 37289 24225 37323 24259
rect 37323 24225 37332 24259
rect 37280 24216 37332 24225
rect 38752 24216 38804 24268
rect 39764 24216 39816 24268
rect 40776 24216 40828 24268
rect 32680 24148 32732 24200
rect 34612 24148 34664 24200
rect 34980 24148 35032 24200
rect 35624 24191 35676 24200
rect 35624 24157 35633 24191
rect 35633 24157 35667 24191
rect 35667 24157 35676 24191
rect 35624 24148 35676 24157
rect 34796 24080 34848 24132
rect 35164 24080 35216 24132
rect 36084 24080 36136 24132
rect 39580 24148 39632 24200
rect 40040 24191 40092 24200
rect 40040 24157 40049 24191
rect 40049 24157 40083 24191
rect 40083 24157 40092 24191
rect 40040 24148 40092 24157
rect 40408 24191 40460 24200
rect 40408 24157 40417 24191
rect 40417 24157 40451 24191
rect 40451 24157 40460 24191
rect 40408 24148 40460 24157
rect 41788 24148 41840 24200
rect 31484 24012 31536 24064
rect 32496 24012 32548 24064
rect 32956 24012 33008 24064
rect 34520 24012 34572 24064
rect 36728 24012 36780 24064
rect 37556 24012 37608 24064
rect 39304 24123 39356 24132
rect 39304 24089 39313 24123
rect 39313 24089 39347 24123
rect 39347 24089 39356 24123
rect 39304 24080 39356 24089
rect 39488 24123 39540 24132
rect 39488 24089 39497 24123
rect 39497 24089 39531 24123
rect 39531 24089 39540 24123
rect 39488 24080 39540 24089
rect 39028 24012 39080 24064
rect 40684 24080 40736 24132
rect 39764 24012 39816 24064
rect 40224 24055 40276 24064
rect 40224 24021 40233 24055
rect 40233 24021 40267 24055
rect 40267 24021 40276 24055
rect 40224 24012 40276 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 3976 23851 4028 23860
rect 3976 23817 3985 23851
rect 3985 23817 4019 23851
rect 4019 23817 4028 23851
rect 3976 23808 4028 23817
rect 2504 23740 2556 23792
rect 2688 23740 2740 23792
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 2780 23672 2832 23724
rect 3792 23715 3844 23724
rect 3792 23681 3801 23715
rect 3801 23681 3835 23715
rect 3835 23681 3844 23715
rect 3792 23672 3844 23681
rect 4620 23783 4672 23792
rect 4620 23749 4629 23783
rect 4629 23749 4663 23783
rect 4663 23749 4672 23783
rect 4620 23740 4672 23749
rect 7748 23808 7800 23860
rect 8944 23851 8996 23860
rect 8944 23817 8953 23851
rect 8953 23817 8987 23851
rect 8987 23817 8996 23851
rect 8944 23808 8996 23817
rect 7288 23740 7340 23792
rect 5724 23672 5776 23724
rect 6552 23672 6604 23724
rect 7196 23715 7248 23724
rect 7196 23681 7205 23715
rect 7205 23681 7239 23715
rect 7239 23681 7248 23715
rect 7196 23672 7248 23681
rect 7380 23715 7432 23724
rect 7380 23681 7389 23715
rect 7389 23681 7423 23715
rect 7423 23681 7432 23715
rect 7380 23672 7432 23681
rect 2136 23579 2188 23588
rect 2136 23545 2145 23579
rect 2145 23545 2179 23579
rect 2179 23545 2188 23579
rect 2136 23536 2188 23545
rect 4252 23604 4304 23656
rect 6000 23604 6052 23656
rect 7656 23672 7708 23724
rect 4160 23536 4212 23588
rect 6828 23536 6880 23588
rect 9036 23672 9088 23724
rect 9404 23672 9456 23724
rect 12992 23808 13044 23860
rect 13084 23808 13136 23860
rect 10232 23783 10284 23792
rect 10232 23749 10266 23783
rect 10266 23749 10284 23783
rect 10232 23740 10284 23749
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 11796 23672 11848 23724
rect 14280 23740 14332 23792
rect 9864 23604 9916 23656
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 5816 23468 5868 23520
rect 7196 23468 7248 23520
rect 7288 23468 7340 23520
rect 10232 23468 10284 23520
rect 10324 23468 10376 23520
rect 13268 23536 13320 23588
rect 18052 23808 18104 23860
rect 18420 23808 18472 23860
rect 19708 23808 19760 23860
rect 20260 23808 20312 23860
rect 20444 23808 20496 23860
rect 21916 23851 21968 23860
rect 21916 23817 21925 23851
rect 21925 23817 21959 23851
rect 21959 23817 21968 23851
rect 21916 23808 21968 23817
rect 22468 23808 22520 23860
rect 23020 23808 23072 23860
rect 19432 23740 19484 23792
rect 19800 23740 19852 23792
rect 20168 23740 20220 23792
rect 13912 23647 13964 23656
rect 13912 23613 13921 23647
rect 13921 23613 13955 23647
rect 13955 23613 13964 23647
rect 13912 23604 13964 23613
rect 14004 23647 14056 23656
rect 14004 23613 14013 23647
rect 14013 23613 14047 23647
rect 14047 23613 14056 23647
rect 14004 23604 14056 23613
rect 16396 23715 16448 23724
rect 16396 23681 16405 23715
rect 16405 23681 16439 23715
rect 16439 23681 16448 23715
rect 16396 23672 16448 23681
rect 16580 23672 16632 23724
rect 17040 23715 17092 23724
rect 17040 23681 17049 23715
rect 17049 23681 17083 23715
rect 17083 23681 17092 23715
rect 17040 23672 17092 23681
rect 17592 23672 17644 23724
rect 17132 23647 17184 23656
rect 17132 23613 17141 23647
rect 17141 23613 17175 23647
rect 17175 23613 17184 23647
rect 17132 23604 17184 23613
rect 17960 23715 18012 23724
rect 17960 23681 18005 23715
rect 18005 23681 18012 23715
rect 17960 23672 18012 23681
rect 18328 23672 18380 23724
rect 18604 23604 18656 23656
rect 18788 23715 18840 23724
rect 18788 23681 18797 23715
rect 18797 23681 18831 23715
rect 18831 23681 18840 23715
rect 18788 23672 18840 23681
rect 20076 23672 20128 23724
rect 22560 23740 22612 23792
rect 24952 23808 25004 23860
rect 27160 23808 27212 23860
rect 22744 23672 22796 23724
rect 26148 23740 26200 23792
rect 26240 23740 26292 23792
rect 27344 23740 27396 23792
rect 27436 23740 27488 23792
rect 30748 23808 30800 23860
rect 27988 23740 28040 23792
rect 24216 23672 24268 23724
rect 24308 23715 24360 23724
rect 24308 23681 24317 23715
rect 24317 23681 24351 23715
rect 24351 23681 24360 23715
rect 24308 23672 24360 23681
rect 26056 23672 26108 23724
rect 27804 23672 27856 23724
rect 19248 23604 19300 23656
rect 19340 23604 19392 23656
rect 18052 23536 18104 23588
rect 19892 23536 19944 23588
rect 25044 23604 25096 23656
rect 26792 23604 26844 23656
rect 27896 23604 27948 23656
rect 28724 23672 28776 23724
rect 30656 23672 30708 23724
rect 28080 23647 28132 23656
rect 28080 23613 28089 23647
rect 28089 23613 28123 23647
rect 28123 23613 28132 23647
rect 28080 23604 28132 23613
rect 28356 23604 28408 23656
rect 31024 23672 31076 23724
rect 31668 23808 31720 23860
rect 34980 23851 35032 23860
rect 34980 23817 35005 23851
rect 35005 23817 35032 23851
rect 34980 23808 35032 23817
rect 31300 23783 31352 23792
rect 31300 23749 31309 23783
rect 31309 23749 31343 23783
rect 31343 23749 31352 23783
rect 31300 23740 31352 23749
rect 34704 23740 34756 23792
rect 25688 23536 25740 23588
rect 25872 23536 25924 23588
rect 27252 23536 27304 23588
rect 12992 23468 13044 23520
rect 13820 23468 13872 23520
rect 15660 23468 15712 23520
rect 15936 23468 15988 23520
rect 17960 23468 18012 23520
rect 18604 23468 18656 23520
rect 20168 23511 20220 23520
rect 20168 23477 20177 23511
rect 20177 23477 20211 23511
rect 20211 23477 20220 23511
rect 20168 23468 20220 23477
rect 24308 23468 24360 23520
rect 25136 23468 25188 23520
rect 25780 23468 25832 23520
rect 31760 23672 31812 23724
rect 32312 23672 32364 23724
rect 34612 23672 34664 23724
rect 35164 23740 35216 23792
rect 34980 23672 35032 23724
rect 35440 23715 35492 23724
rect 35440 23681 35449 23715
rect 35449 23681 35483 23715
rect 35483 23681 35492 23715
rect 35440 23672 35492 23681
rect 37004 23672 37056 23724
rect 37556 23783 37608 23792
rect 37556 23749 37565 23783
rect 37565 23749 37599 23783
rect 37599 23749 37608 23783
rect 37556 23740 37608 23749
rect 40408 23808 40460 23860
rect 39764 23783 39816 23792
rect 39764 23749 39773 23783
rect 39773 23749 39807 23783
rect 39807 23749 39816 23783
rect 39764 23740 39816 23749
rect 41052 23740 41104 23792
rect 41696 23783 41748 23792
rect 41696 23749 41705 23783
rect 41705 23749 41739 23783
rect 41739 23749 41748 23783
rect 41696 23740 41748 23749
rect 41144 23672 41196 23724
rect 29736 23536 29788 23588
rect 32772 23604 32824 23656
rect 34520 23604 34572 23656
rect 36176 23604 36228 23656
rect 38752 23604 38804 23656
rect 39028 23647 39080 23656
rect 39028 23613 39037 23647
rect 39037 23613 39071 23647
rect 39071 23613 39080 23647
rect 39028 23604 39080 23613
rect 41420 23672 41472 23724
rect 41604 23715 41656 23724
rect 41604 23681 41613 23715
rect 41613 23681 41647 23715
rect 41647 23681 41656 23715
rect 41604 23672 41656 23681
rect 42064 23672 42116 23724
rect 31668 23536 31720 23588
rect 35716 23536 35768 23588
rect 31484 23511 31536 23520
rect 31484 23477 31493 23511
rect 31493 23477 31527 23511
rect 31527 23477 31536 23511
rect 31484 23468 31536 23477
rect 34796 23468 34848 23520
rect 34980 23511 35032 23520
rect 34980 23477 34989 23511
rect 34989 23477 35023 23511
rect 35023 23477 35032 23511
rect 34980 23468 35032 23477
rect 36544 23468 36596 23520
rect 41328 23511 41380 23520
rect 41328 23477 41337 23511
rect 41337 23477 41371 23511
rect 41371 23477 41380 23511
rect 41328 23468 41380 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1400 23307 1452 23316
rect 1400 23273 1409 23307
rect 1409 23273 1443 23307
rect 1443 23273 1452 23307
rect 1400 23264 1452 23273
rect 5448 23307 5500 23316
rect 5448 23273 5457 23307
rect 5457 23273 5491 23307
rect 5491 23273 5500 23307
rect 5448 23264 5500 23273
rect 5632 23307 5684 23316
rect 5632 23273 5641 23307
rect 5641 23273 5675 23307
rect 5675 23273 5684 23307
rect 5632 23264 5684 23273
rect 112 23128 164 23180
rect 7380 23239 7432 23248
rect 7380 23205 7389 23239
rect 7389 23205 7423 23239
rect 7423 23205 7432 23239
rect 7380 23196 7432 23205
rect 12440 23196 12492 23248
rect 12164 23128 12216 23180
rect 15476 23196 15528 23248
rect 17040 23196 17092 23248
rect 13912 23128 13964 23180
rect 14188 23171 14240 23180
rect 14188 23137 14197 23171
rect 14197 23137 14231 23171
rect 14231 23137 14240 23171
rect 14188 23128 14240 23137
rect 14556 23128 14608 23180
rect 3240 23060 3292 23112
rect 7104 23103 7156 23112
rect 7104 23069 7113 23103
rect 7113 23069 7147 23103
rect 7147 23069 7156 23103
rect 7104 23060 7156 23069
rect 7196 23060 7248 23112
rect 7380 23060 7432 23112
rect 7472 23103 7524 23112
rect 7472 23069 7481 23103
rect 7481 23069 7515 23103
rect 7515 23069 7524 23103
rect 7472 23060 7524 23069
rect 7656 23060 7708 23112
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 10232 23060 10284 23112
rect 12992 23060 13044 23112
rect 13176 23060 13228 23112
rect 13636 23103 13688 23112
rect 13636 23069 13645 23103
rect 13645 23069 13679 23103
rect 13679 23069 13688 23103
rect 13636 23060 13688 23069
rect 2412 22992 2464 23044
rect 2872 23035 2924 23044
rect 2872 23001 2881 23035
rect 2881 23001 2915 23035
rect 2915 23001 2924 23035
rect 2872 22992 2924 23001
rect 5356 22992 5408 23044
rect 13728 22992 13780 23044
rect 14464 23103 14516 23112
rect 14464 23069 14473 23103
rect 14473 23069 14507 23103
rect 14507 23069 14516 23103
rect 14464 23060 14516 23069
rect 16672 23128 16724 23180
rect 14832 23103 14884 23112
rect 14832 23069 14841 23103
rect 14841 23069 14875 23103
rect 14875 23069 14884 23103
rect 14832 23060 14884 23069
rect 15108 23103 15160 23112
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 15292 23103 15344 23112
rect 15292 23069 15301 23103
rect 15301 23069 15335 23103
rect 15335 23069 15344 23103
rect 15292 23060 15344 23069
rect 6000 22924 6052 22976
rect 7748 22967 7800 22976
rect 7748 22933 7757 22967
rect 7757 22933 7791 22967
rect 7791 22933 7800 22967
rect 7748 22924 7800 22933
rect 12624 22924 12676 22976
rect 14188 22967 14240 22976
rect 14188 22933 14197 22967
rect 14197 22933 14231 22967
rect 14231 22933 14240 22967
rect 14188 22924 14240 22933
rect 15568 23060 15620 23112
rect 19524 23128 19576 23180
rect 19892 23171 19944 23180
rect 19892 23137 19901 23171
rect 19901 23137 19935 23171
rect 19935 23137 19944 23171
rect 19892 23128 19944 23137
rect 18144 23060 18196 23112
rect 21732 23264 21784 23316
rect 21916 23307 21968 23316
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 28724 23264 28776 23316
rect 29000 23196 29052 23248
rect 30564 23128 30616 23180
rect 31300 23128 31352 23180
rect 32036 23128 32088 23180
rect 32220 23128 32272 23180
rect 34704 23196 34756 23248
rect 22836 23060 22888 23112
rect 24676 23060 24728 23112
rect 25504 23060 25556 23112
rect 25596 23103 25648 23112
rect 25596 23069 25605 23103
rect 25605 23069 25639 23103
rect 25639 23069 25648 23103
rect 25596 23060 25648 23069
rect 25872 23103 25924 23112
rect 25872 23069 25881 23103
rect 25881 23069 25915 23103
rect 25915 23069 25924 23103
rect 25872 23060 25924 23069
rect 25964 23103 26016 23112
rect 25964 23069 25973 23103
rect 25973 23069 26007 23103
rect 26007 23069 26016 23103
rect 25964 23060 26016 23069
rect 27712 23060 27764 23112
rect 28908 23060 28960 23112
rect 31484 23103 31536 23112
rect 31484 23069 31493 23103
rect 31493 23069 31527 23103
rect 31527 23069 31536 23103
rect 31484 23060 31536 23069
rect 33416 23060 33468 23112
rect 33508 23103 33560 23112
rect 33508 23069 33517 23103
rect 33517 23069 33551 23103
rect 33551 23069 33560 23103
rect 33508 23060 33560 23069
rect 34520 23171 34572 23180
rect 34520 23137 34529 23171
rect 34529 23137 34563 23171
rect 34563 23137 34572 23171
rect 34520 23128 34572 23137
rect 35532 23128 35584 23180
rect 35716 23171 35768 23180
rect 35716 23137 35725 23171
rect 35725 23137 35759 23171
rect 35759 23137 35768 23171
rect 35716 23128 35768 23137
rect 35256 23060 35308 23112
rect 35992 23128 36044 23180
rect 15936 23035 15988 23044
rect 15936 23001 15945 23035
rect 15945 23001 15979 23035
rect 15979 23001 15988 23035
rect 15936 22992 15988 23001
rect 18052 22992 18104 23044
rect 19616 23035 19668 23044
rect 19616 23001 19625 23035
rect 19625 23001 19659 23035
rect 19659 23001 19668 23035
rect 19616 22992 19668 23001
rect 25228 22992 25280 23044
rect 29092 22992 29144 23044
rect 31760 22992 31812 23044
rect 16580 22924 16632 22976
rect 18788 22924 18840 22976
rect 22468 22924 22520 22976
rect 23388 22924 23440 22976
rect 26424 22924 26476 22976
rect 27160 22924 27212 22976
rect 30288 22924 30340 22976
rect 32128 22967 32180 22976
rect 32128 22933 32137 22967
rect 32137 22933 32171 22967
rect 32171 22933 32180 22967
rect 32128 22924 32180 22933
rect 36544 23103 36596 23111
rect 36544 23069 36553 23103
rect 36553 23069 36587 23103
rect 36587 23069 36596 23103
rect 36544 23059 36596 23069
rect 38660 23103 38712 23112
rect 38660 23069 38669 23103
rect 38669 23069 38703 23103
rect 38703 23069 38712 23103
rect 38660 23060 38712 23069
rect 39304 23264 39356 23316
rect 39396 23103 39448 23112
rect 39396 23069 39405 23103
rect 39405 23069 39439 23103
rect 39439 23069 39448 23103
rect 39396 23060 39448 23069
rect 41696 23264 41748 23316
rect 40040 23060 40092 23112
rect 40408 23103 40460 23112
rect 40408 23069 40417 23103
rect 40417 23069 40451 23103
rect 40451 23069 40460 23103
rect 40408 23060 40460 23069
rect 34612 22924 34664 22976
rect 34888 22924 34940 22976
rect 34980 22924 35032 22976
rect 36268 22967 36320 22976
rect 36268 22933 36277 22967
rect 36277 22933 36311 22967
rect 36311 22933 36320 22967
rect 36268 22924 36320 22933
rect 37004 22992 37056 23044
rect 37096 22992 37148 23044
rect 36820 22924 36872 22976
rect 37740 22924 37792 22976
rect 41144 22992 41196 23044
rect 41328 22924 41380 22976
rect 42064 22924 42116 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 2412 22652 2464 22704
rect 5724 22720 5776 22772
rect 7104 22720 7156 22772
rect 7932 22763 7984 22772
rect 7932 22729 7941 22763
rect 7941 22729 7975 22763
rect 7975 22729 7984 22763
rect 7932 22720 7984 22729
rect 9864 22720 9916 22772
rect 12624 22763 12676 22772
rect 12624 22729 12633 22763
rect 12633 22729 12667 22763
rect 12667 22729 12676 22763
rect 12624 22720 12676 22729
rect 14464 22720 14516 22772
rect 15292 22720 15344 22772
rect 5540 22652 5592 22704
rect 5632 22652 5684 22704
rect 8024 22695 8076 22704
rect 8024 22661 8033 22695
rect 8033 22661 8067 22695
rect 8067 22661 8076 22695
rect 8024 22652 8076 22661
rect 7748 22627 7800 22636
rect 7748 22593 7757 22627
rect 7757 22593 7791 22627
rect 7791 22593 7800 22627
rect 7748 22584 7800 22593
rect 10140 22652 10192 22704
rect 11152 22652 11204 22704
rect 12072 22652 12124 22704
rect 13728 22652 13780 22704
rect 14188 22652 14240 22704
rect 16488 22720 16540 22772
rect 18052 22720 18104 22772
rect 17592 22695 17644 22704
rect 17592 22661 17601 22695
rect 17601 22661 17635 22695
rect 17635 22661 17644 22695
rect 17592 22652 17644 22661
rect 18788 22695 18840 22704
rect 18788 22661 18797 22695
rect 18797 22661 18831 22695
rect 18831 22661 18840 22695
rect 18788 22652 18840 22661
rect 19616 22720 19668 22772
rect 19800 22720 19852 22772
rect 20720 22695 20772 22704
rect 20720 22661 20729 22695
rect 20729 22661 20763 22695
rect 20763 22661 20772 22695
rect 20720 22652 20772 22661
rect 2780 22516 2832 22568
rect 3240 22516 3292 22568
rect 4712 22516 4764 22568
rect 7656 22559 7708 22568
rect 7656 22525 7665 22559
rect 7665 22525 7699 22559
rect 7699 22525 7708 22559
rect 7656 22516 7708 22525
rect 1400 22423 1452 22432
rect 1400 22389 1409 22423
rect 1409 22389 1443 22423
rect 1443 22389 1452 22423
rect 1400 22380 1452 22389
rect 4804 22380 4856 22432
rect 6828 22380 6880 22432
rect 7748 22380 7800 22432
rect 11428 22584 11480 22636
rect 14280 22627 14332 22636
rect 14280 22593 14289 22627
rect 14289 22593 14323 22627
rect 14323 22593 14332 22627
rect 14280 22584 14332 22593
rect 16212 22627 16264 22636
rect 16212 22593 16221 22627
rect 16221 22593 16255 22627
rect 16255 22593 16264 22627
rect 16212 22584 16264 22593
rect 17960 22627 18012 22636
rect 17960 22593 17969 22627
rect 17969 22593 18003 22627
rect 18003 22593 18012 22627
rect 17960 22584 18012 22593
rect 18144 22627 18196 22636
rect 18144 22593 18153 22627
rect 18153 22593 18187 22627
rect 18187 22593 18196 22627
rect 18144 22584 18196 22593
rect 18236 22627 18288 22636
rect 18236 22593 18245 22627
rect 18245 22593 18279 22627
rect 18279 22593 18288 22627
rect 18236 22584 18288 22593
rect 20628 22627 20680 22636
rect 20628 22593 20637 22627
rect 20637 22593 20671 22627
rect 20671 22593 20680 22627
rect 20628 22584 20680 22593
rect 22560 22720 22612 22772
rect 24216 22763 24268 22772
rect 24216 22729 24225 22763
rect 24225 22729 24259 22763
rect 24259 22729 24268 22763
rect 24216 22720 24268 22729
rect 22468 22652 22520 22704
rect 14004 22559 14056 22568
rect 14004 22525 14013 22559
rect 14013 22525 14047 22559
rect 14047 22525 14056 22559
rect 14004 22516 14056 22525
rect 15568 22516 15620 22568
rect 16672 22516 16724 22568
rect 12440 22448 12492 22500
rect 21456 22627 21508 22636
rect 21456 22593 21465 22627
rect 21465 22593 21499 22627
rect 21499 22593 21508 22627
rect 24676 22695 24728 22704
rect 24676 22661 24685 22695
rect 24685 22661 24719 22695
rect 24719 22661 24728 22695
rect 24676 22652 24728 22661
rect 24768 22652 24820 22704
rect 24860 22652 24912 22704
rect 25596 22720 25648 22772
rect 26148 22763 26200 22772
rect 26148 22729 26157 22763
rect 26157 22729 26191 22763
rect 26191 22729 26200 22763
rect 26148 22720 26200 22729
rect 26240 22720 26292 22772
rect 21456 22584 21508 22593
rect 23112 22584 23164 22636
rect 27896 22652 27948 22704
rect 30288 22695 30340 22704
rect 30288 22661 30297 22695
rect 30297 22661 30331 22695
rect 30331 22661 30340 22695
rect 30288 22652 30340 22661
rect 31760 22763 31812 22772
rect 31760 22729 31769 22763
rect 31769 22729 31803 22763
rect 31803 22729 31812 22763
rect 31760 22720 31812 22729
rect 32496 22720 32548 22772
rect 33416 22763 33468 22772
rect 33416 22729 33425 22763
rect 33425 22729 33459 22763
rect 33459 22729 33468 22763
rect 33416 22720 33468 22729
rect 33508 22720 33560 22772
rect 33232 22652 33284 22704
rect 34888 22695 34940 22704
rect 34888 22661 34897 22695
rect 34897 22661 34931 22695
rect 34931 22661 34940 22695
rect 34888 22652 34940 22661
rect 35256 22763 35308 22772
rect 35256 22729 35265 22763
rect 35265 22729 35299 22763
rect 35299 22729 35308 22763
rect 35256 22720 35308 22729
rect 36176 22720 36228 22772
rect 25504 22584 25556 22636
rect 21088 22448 21140 22500
rect 21824 22559 21876 22568
rect 21824 22525 21833 22559
rect 21833 22525 21867 22559
rect 21867 22525 21876 22559
rect 21824 22516 21876 22525
rect 22376 22516 22428 22568
rect 23756 22516 23808 22568
rect 24124 22448 24176 22500
rect 24860 22516 24912 22568
rect 25780 22627 25832 22636
rect 25780 22593 25789 22627
rect 25789 22593 25823 22627
rect 25823 22593 25832 22627
rect 25780 22584 25832 22593
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 27712 22584 27764 22636
rect 28172 22584 28224 22636
rect 32128 22584 32180 22636
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 36268 22652 36320 22704
rect 35440 22627 35492 22636
rect 35440 22593 35449 22627
rect 35449 22593 35483 22627
rect 35483 22593 35492 22627
rect 35440 22584 35492 22593
rect 37188 22720 37240 22772
rect 38016 22720 38068 22772
rect 38200 22720 38252 22772
rect 40316 22763 40368 22772
rect 40316 22729 40325 22763
rect 40325 22729 40359 22763
rect 40359 22729 40368 22763
rect 40316 22720 40368 22729
rect 41236 22720 41288 22772
rect 26240 22516 26292 22568
rect 26976 22516 27028 22568
rect 34796 22516 34848 22568
rect 35348 22516 35400 22568
rect 37740 22584 37792 22636
rect 42064 22652 42116 22704
rect 40960 22584 41012 22636
rect 41972 22584 42024 22636
rect 36452 22516 36504 22568
rect 26516 22448 26568 22500
rect 28080 22448 28132 22500
rect 31852 22448 31904 22500
rect 41328 22516 41380 22568
rect 12256 22423 12308 22432
rect 12256 22389 12265 22423
rect 12265 22389 12299 22423
rect 12299 22389 12308 22423
rect 12256 22380 12308 22389
rect 12808 22380 12860 22432
rect 16396 22423 16448 22432
rect 16396 22389 16405 22423
rect 16405 22389 16439 22423
rect 16439 22389 16448 22423
rect 16396 22380 16448 22389
rect 17500 22380 17552 22432
rect 20444 22423 20496 22432
rect 20444 22389 20453 22423
rect 20453 22389 20487 22423
rect 20487 22389 20496 22423
rect 20444 22380 20496 22389
rect 20536 22380 20588 22432
rect 21732 22380 21784 22432
rect 22560 22380 22612 22432
rect 25964 22423 26016 22432
rect 25964 22389 25973 22423
rect 25973 22389 26007 22423
rect 26007 22389 26016 22423
rect 25964 22380 26016 22389
rect 28540 22380 28592 22432
rect 39396 22448 39448 22500
rect 42156 22448 42208 22500
rect 36912 22423 36964 22432
rect 36912 22389 36921 22423
rect 36921 22389 36955 22423
rect 36955 22389 36964 22423
rect 36912 22380 36964 22389
rect 37556 22380 37608 22432
rect 40132 22380 40184 22432
rect 40684 22423 40736 22432
rect 40684 22389 40693 22423
rect 40693 22389 40727 22423
rect 40727 22389 40736 22423
rect 40684 22380 40736 22389
rect 40960 22380 41012 22432
rect 41144 22380 41196 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 5540 22176 5592 22228
rect 7656 22176 7708 22228
rect 14464 22176 14516 22228
rect 15108 22176 15160 22228
rect 3240 22040 3292 22092
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 4252 22015 4304 22024
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 7104 22108 7156 22160
rect 6368 21972 6420 22024
rect 6828 22015 6880 22024
rect 6828 21981 6837 22015
rect 6837 21981 6871 22015
rect 6871 21981 6880 22015
rect 6828 21972 6880 21981
rect 10140 22040 10192 22092
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 7472 22015 7524 22024
rect 7472 21981 7481 22015
rect 7481 21981 7515 22015
rect 7515 21981 7524 22015
rect 7472 21972 7524 21981
rect 7748 22015 7800 22024
rect 7748 21981 7757 22015
rect 7757 21981 7791 22015
rect 7791 21981 7800 22015
rect 7748 21972 7800 21981
rect 8852 21972 8904 22024
rect 11612 21972 11664 22024
rect 12808 22015 12860 22024
rect 12808 21981 12842 22015
rect 12842 21981 12860 22015
rect 12808 21972 12860 21981
rect 16396 22176 16448 22228
rect 17500 22219 17552 22228
rect 17500 22185 17530 22219
rect 17530 22185 17552 22219
rect 17500 22176 17552 22185
rect 18236 22176 18288 22228
rect 20628 22176 20680 22228
rect 16948 22108 17000 22160
rect 23112 22219 23164 22228
rect 23112 22185 23121 22219
rect 23121 22185 23155 22219
rect 23155 22185 23164 22219
rect 23112 22176 23164 22185
rect 25780 22176 25832 22228
rect 34060 22176 34112 22228
rect 34612 22176 34664 22228
rect 36912 22176 36964 22228
rect 41328 22176 41380 22228
rect 15476 22040 15528 22092
rect 5908 21904 5960 21956
rect 6460 21904 6512 21956
rect 9036 21904 9088 21956
rect 9404 21947 9456 21956
rect 9404 21913 9413 21947
rect 9413 21913 9447 21947
rect 9447 21913 9456 21947
rect 9404 21904 9456 21913
rect 1308 21836 1360 21888
rect 5724 21836 5776 21888
rect 6184 21836 6236 21888
rect 6920 21879 6972 21888
rect 6920 21845 6929 21879
rect 6929 21845 6963 21879
rect 6963 21845 6972 21879
rect 6920 21836 6972 21845
rect 7012 21836 7064 21888
rect 7932 21836 7984 21888
rect 11152 21947 11204 21956
rect 11152 21913 11161 21947
rect 11161 21913 11195 21947
rect 11195 21913 11204 21947
rect 11152 21904 11204 21913
rect 15384 21947 15436 21956
rect 15384 21913 15393 21947
rect 15393 21913 15427 21947
rect 15427 21913 15436 21947
rect 15384 21904 15436 21913
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 15660 22015 15712 22024
rect 15660 21981 15669 22015
rect 15669 21981 15703 22015
rect 15703 21981 15712 22015
rect 15660 21972 15712 21981
rect 16304 22040 16356 22092
rect 16672 22040 16724 22092
rect 24032 22108 24084 22160
rect 27896 22108 27948 22160
rect 23756 22083 23808 22092
rect 23756 22049 23765 22083
rect 23765 22049 23799 22083
rect 23799 22049 23808 22083
rect 23756 22040 23808 22049
rect 24124 22040 24176 22092
rect 31760 22108 31812 22160
rect 31208 22040 31260 22092
rect 16396 21972 16448 22024
rect 16856 21904 16908 21956
rect 15016 21879 15068 21888
rect 15016 21845 15025 21879
rect 15025 21845 15059 21879
rect 15059 21845 15068 21879
rect 15016 21836 15068 21845
rect 16304 21879 16356 21888
rect 16304 21845 16313 21879
rect 16313 21845 16347 21879
rect 16347 21845 16356 21879
rect 16304 21836 16356 21845
rect 18880 21972 18932 22024
rect 21456 22015 21508 22024
rect 21456 21981 21465 22015
rect 21465 21981 21499 22015
rect 21499 21981 21508 22015
rect 21456 21972 21508 21981
rect 21732 22015 21784 22024
rect 21732 21981 21766 22015
rect 21766 21981 21784 22015
rect 21732 21972 21784 21981
rect 23204 21972 23256 22024
rect 18512 21904 18564 21956
rect 20444 21904 20496 21956
rect 18144 21836 18196 21888
rect 20628 21836 20680 21888
rect 20996 21836 21048 21888
rect 21824 21836 21876 21888
rect 22836 21879 22888 21888
rect 22836 21845 22845 21879
rect 22845 21845 22879 21879
rect 22879 21845 22888 21879
rect 22836 21836 22888 21845
rect 23296 21836 23348 21888
rect 24952 21836 25004 21888
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 28816 21972 28868 22024
rect 25596 21904 25648 21956
rect 26424 21904 26476 21956
rect 26976 21904 27028 21956
rect 28172 21904 28224 21956
rect 28448 21904 28500 21956
rect 29000 21947 29052 21956
rect 29000 21913 29009 21947
rect 29009 21913 29043 21947
rect 29043 21913 29052 21947
rect 29000 21904 29052 21913
rect 30104 21904 30156 21956
rect 30932 22015 30984 22024
rect 30932 21981 30941 22015
rect 30941 21981 30975 22015
rect 30975 21981 30984 22015
rect 30932 21972 30984 21981
rect 31392 22015 31444 22024
rect 31392 21981 31401 22015
rect 31401 21981 31435 22015
rect 31435 21981 31444 22015
rect 31392 21972 31444 21981
rect 34796 22040 34848 22092
rect 32128 22015 32180 22024
rect 32128 21981 32137 22015
rect 32137 21981 32171 22015
rect 32171 21981 32180 22015
rect 32128 21972 32180 21981
rect 25688 21836 25740 21888
rect 26608 21836 26660 21888
rect 27068 21836 27120 21888
rect 29552 21879 29604 21888
rect 29552 21845 29561 21879
rect 29561 21845 29595 21879
rect 29595 21845 29604 21879
rect 29552 21836 29604 21845
rect 29828 21836 29880 21888
rect 31116 21879 31168 21888
rect 31116 21845 31125 21879
rect 31125 21845 31159 21879
rect 31159 21845 31168 21879
rect 31116 21836 31168 21845
rect 31484 21947 31536 21956
rect 31484 21913 31493 21947
rect 31493 21913 31527 21947
rect 31527 21913 31536 21947
rect 31484 21904 31536 21913
rect 33140 21972 33192 22024
rect 32404 21947 32456 21956
rect 32404 21913 32438 21947
rect 32438 21913 32456 21947
rect 32404 21904 32456 21913
rect 33416 21904 33468 21956
rect 32496 21836 32548 21888
rect 33048 21836 33100 21888
rect 33508 21879 33560 21888
rect 33508 21845 33517 21879
rect 33517 21845 33551 21879
rect 33551 21845 33560 21879
rect 34428 21972 34480 22024
rect 36268 22083 36320 22092
rect 36268 22049 36277 22083
rect 36277 22049 36311 22083
rect 36311 22049 36320 22083
rect 36268 22040 36320 22049
rect 36544 22040 36596 22092
rect 38016 22083 38068 22092
rect 38016 22049 38025 22083
rect 38025 22049 38059 22083
rect 38059 22049 38068 22083
rect 38016 22040 38068 22049
rect 41972 22083 42024 22092
rect 41972 22049 41981 22083
rect 41981 22049 42015 22083
rect 42015 22049 42024 22083
rect 41972 22040 42024 22049
rect 38752 21972 38804 22024
rect 40408 21972 40460 22024
rect 41328 22015 41380 22024
rect 41328 21981 41337 22015
rect 41337 21981 41371 22015
rect 41371 21981 41380 22015
rect 41328 21972 41380 21981
rect 34704 21904 34756 21956
rect 35072 21947 35124 21956
rect 35072 21913 35081 21947
rect 35081 21913 35115 21947
rect 35115 21913 35124 21947
rect 35072 21904 35124 21913
rect 38200 21947 38252 21956
rect 38200 21913 38209 21947
rect 38209 21913 38243 21947
rect 38243 21913 38252 21947
rect 38200 21904 38252 21913
rect 40132 21947 40184 21956
rect 40132 21913 40166 21947
rect 40166 21913 40184 21947
rect 40132 21904 40184 21913
rect 33508 21836 33560 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 4712 21632 4764 21684
rect 4252 21564 4304 21616
rect 3148 21471 3200 21480
rect 3148 21437 3157 21471
rect 3157 21437 3191 21471
rect 3191 21437 3200 21471
rect 3148 21428 3200 21437
rect 4804 21496 4856 21548
rect 5816 21632 5868 21684
rect 6828 21632 6880 21684
rect 9404 21632 9456 21684
rect 12992 21675 13044 21684
rect 12992 21641 13001 21675
rect 13001 21641 13035 21675
rect 13035 21641 13044 21675
rect 12992 21632 13044 21641
rect 15568 21675 15620 21684
rect 15568 21641 15577 21675
rect 15577 21641 15611 21675
rect 15611 21641 15620 21675
rect 15568 21632 15620 21641
rect 17224 21632 17276 21684
rect 21364 21632 21416 21684
rect 22652 21632 22704 21684
rect 24860 21675 24912 21684
rect 24860 21641 24869 21675
rect 24869 21641 24903 21675
rect 24903 21641 24912 21675
rect 24860 21632 24912 21641
rect 25596 21675 25648 21684
rect 25596 21641 25605 21675
rect 25605 21641 25639 21675
rect 25639 21641 25648 21675
rect 25596 21632 25648 21641
rect 25688 21632 25740 21684
rect 5264 21539 5316 21548
rect 5264 21505 5273 21539
rect 5273 21505 5307 21539
rect 5307 21505 5316 21539
rect 5264 21496 5316 21505
rect 5724 21564 5776 21616
rect 7104 21564 7156 21616
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 5264 21360 5316 21412
rect 6276 21428 6328 21480
rect 6644 21428 6696 21480
rect 6736 21471 6788 21480
rect 6736 21437 6745 21471
rect 6745 21437 6779 21471
rect 6779 21437 6788 21471
rect 6736 21428 6788 21437
rect 7288 21428 7340 21480
rect 11152 21564 11204 21616
rect 12256 21564 12308 21616
rect 16580 21564 16632 21616
rect 16948 21564 17000 21616
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 8852 21471 8904 21480
rect 8852 21437 8861 21471
rect 8861 21437 8895 21471
rect 8895 21437 8904 21471
rect 8852 21428 8904 21437
rect 8944 21428 8996 21480
rect 11612 21539 11664 21548
rect 11612 21505 11621 21539
rect 11621 21505 11655 21539
rect 11655 21505 11664 21539
rect 11612 21496 11664 21505
rect 15016 21496 15068 21548
rect 15384 21496 15436 21548
rect 16120 21471 16172 21480
rect 16120 21437 16129 21471
rect 16129 21437 16163 21471
rect 16163 21437 16172 21471
rect 16120 21428 16172 21437
rect 16304 21496 16356 21548
rect 20536 21564 20588 21616
rect 23204 21564 23256 21616
rect 24216 21564 24268 21616
rect 25320 21607 25372 21616
rect 25320 21573 25329 21607
rect 25329 21573 25363 21607
rect 25363 21573 25372 21607
rect 25320 21564 25372 21573
rect 18052 21496 18104 21548
rect 18512 21496 18564 21548
rect 18880 21539 18932 21548
rect 18880 21505 18889 21539
rect 18889 21505 18923 21539
rect 18923 21505 18932 21539
rect 18880 21496 18932 21505
rect 19156 21539 19208 21548
rect 19156 21505 19190 21539
rect 19190 21505 19208 21539
rect 19156 21496 19208 21505
rect 17960 21428 18012 21480
rect 2596 21335 2648 21344
rect 2596 21301 2605 21335
rect 2605 21301 2639 21335
rect 2639 21301 2648 21335
rect 2596 21292 2648 21301
rect 6000 21335 6052 21344
rect 6000 21301 6009 21335
rect 6009 21301 6043 21335
rect 6043 21301 6052 21335
rect 6000 21292 6052 21301
rect 6184 21292 6236 21344
rect 7564 21292 7616 21344
rect 14372 21292 14424 21344
rect 17960 21292 18012 21344
rect 21088 21496 21140 21548
rect 22284 21496 22336 21548
rect 21180 21428 21232 21480
rect 25136 21496 25188 21548
rect 25228 21539 25280 21548
rect 25228 21505 25237 21539
rect 25237 21505 25271 21539
rect 25271 21505 25280 21539
rect 25228 21496 25280 21505
rect 25964 21496 26016 21548
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 27528 21496 27580 21548
rect 28356 21675 28408 21684
rect 28356 21641 28365 21675
rect 28365 21641 28399 21675
rect 28399 21641 28408 21675
rect 28356 21632 28408 21641
rect 30932 21632 30984 21684
rect 32404 21675 32456 21684
rect 32404 21641 32413 21675
rect 32413 21641 32447 21675
rect 32447 21641 32456 21675
rect 32404 21632 32456 21641
rect 29552 21564 29604 21616
rect 31484 21564 31536 21616
rect 33048 21564 33100 21616
rect 35072 21632 35124 21684
rect 36452 21632 36504 21684
rect 41328 21675 41380 21684
rect 41328 21641 41337 21675
rect 41337 21641 41371 21675
rect 41371 21641 41380 21675
rect 41328 21632 41380 21641
rect 35348 21564 35400 21616
rect 32496 21496 32548 21548
rect 20628 21360 20680 21412
rect 23204 21471 23256 21480
rect 23204 21437 23213 21471
rect 23213 21437 23247 21471
rect 23247 21437 23256 21471
rect 23204 21428 23256 21437
rect 20444 21292 20496 21344
rect 21824 21335 21876 21344
rect 21824 21301 21833 21335
rect 21833 21301 21867 21335
rect 21867 21301 21876 21335
rect 21824 21292 21876 21301
rect 22468 21360 22520 21412
rect 26608 21428 26660 21480
rect 28448 21471 28500 21480
rect 28448 21437 28457 21471
rect 28457 21437 28491 21471
rect 28491 21437 28500 21471
rect 28448 21428 28500 21437
rect 30104 21428 30156 21480
rect 31852 21471 31904 21480
rect 31852 21437 31861 21471
rect 31861 21437 31895 21471
rect 31895 21437 31904 21471
rect 31852 21428 31904 21437
rect 23756 21292 23808 21344
rect 25964 21292 26016 21344
rect 28816 21292 28868 21344
rect 29920 21292 29972 21344
rect 31208 21335 31260 21344
rect 31208 21301 31217 21335
rect 31217 21301 31251 21335
rect 31251 21301 31260 21335
rect 31208 21292 31260 21301
rect 32588 21360 32640 21412
rect 33416 21496 33468 21548
rect 34060 21539 34112 21548
rect 34060 21505 34069 21539
rect 34069 21505 34103 21539
rect 34103 21505 34112 21539
rect 34060 21496 34112 21505
rect 33692 21428 33744 21480
rect 34612 21496 34664 21548
rect 40408 21564 40460 21616
rect 40684 21496 40736 21548
rect 35624 21471 35676 21480
rect 35624 21437 35633 21471
rect 35633 21437 35667 21471
rect 35667 21437 35676 21471
rect 35624 21428 35676 21437
rect 33140 21292 33192 21344
rect 33784 21335 33836 21344
rect 33784 21301 33793 21335
rect 33793 21301 33827 21335
rect 33827 21301 33836 21335
rect 33784 21292 33836 21301
rect 33876 21335 33928 21344
rect 33876 21301 33885 21335
rect 33885 21301 33919 21335
rect 33919 21301 33928 21335
rect 33876 21292 33928 21301
rect 35992 21292 36044 21344
rect 36728 21292 36780 21344
rect 40224 21292 40276 21344
rect 40960 21292 41012 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 5632 21088 5684 21140
rect 6736 21088 6788 21140
rect 8852 21088 8904 21140
rect 16120 21088 16172 21140
rect 4620 21020 4672 21072
rect 1676 20884 1728 20936
rect 2596 20884 2648 20936
rect 3056 20884 3108 20936
rect 3976 20884 4028 20936
rect 4804 20927 4856 20936
rect 4804 20893 4813 20927
rect 4813 20893 4847 20927
rect 4847 20893 4856 20927
rect 4804 20884 4856 20893
rect 5264 20952 5316 21004
rect 6644 20952 6696 21004
rect 10784 20952 10836 21004
rect 11796 20995 11848 21004
rect 11796 20961 11805 20995
rect 11805 20961 11839 20995
rect 11839 20961 11848 20995
rect 11796 20952 11848 20961
rect 16028 20995 16080 21004
rect 16028 20961 16037 20995
rect 16037 20961 16071 20995
rect 16071 20961 16080 20995
rect 16028 20952 16080 20961
rect 17408 20952 17460 21004
rect 19156 21088 19208 21140
rect 23204 21088 23256 21140
rect 29092 21088 29144 21140
rect 38660 21131 38712 21140
rect 38660 21097 38669 21131
rect 38669 21097 38703 21131
rect 38703 21097 38712 21131
rect 38660 21088 38712 21097
rect 20628 21020 20680 21072
rect 27896 21020 27948 21072
rect 24768 20952 24820 21004
rect 24952 20995 25004 21004
rect 24952 20961 24961 20995
rect 24961 20961 24995 20995
rect 24995 20961 25004 20995
rect 24952 20952 25004 20961
rect 28448 21020 28500 21072
rect 29828 20952 29880 21004
rect 5356 20884 5408 20936
rect 4160 20816 4212 20868
rect 4528 20859 4580 20868
rect 4528 20825 4537 20859
rect 4537 20825 4571 20859
rect 4571 20825 4580 20859
rect 4528 20816 4580 20825
rect 6184 20927 6236 20936
rect 6184 20893 6193 20927
rect 6193 20893 6227 20927
rect 6227 20893 6236 20927
rect 6184 20884 6236 20893
rect 8392 20884 8444 20936
rect 10140 20884 10192 20936
rect 13176 20927 13228 20936
rect 13176 20893 13185 20927
rect 13185 20893 13219 20927
rect 13219 20893 13228 20927
rect 13176 20884 13228 20893
rect 16580 20884 16632 20936
rect 17224 20927 17276 20936
rect 17224 20893 17233 20927
rect 17233 20893 17267 20927
rect 17267 20893 17276 20927
rect 17224 20884 17276 20893
rect 6368 20816 6420 20868
rect 6920 20816 6972 20868
rect 9772 20859 9824 20868
rect 9772 20825 9806 20859
rect 9806 20825 9824 20859
rect 9772 20816 9824 20825
rect 14372 20859 14424 20868
rect 14372 20825 14406 20859
rect 14406 20825 14424 20859
rect 14372 20816 14424 20825
rect 14464 20816 14516 20868
rect 3332 20791 3384 20800
rect 3332 20757 3341 20791
rect 3341 20757 3375 20791
rect 3375 20757 3384 20791
rect 3332 20748 3384 20757
rect 3424 20748 3476 20800
rect 4712 20791 4764 20800
rect 4712 20757 4721 20791
rect 4721 20757 4755 20791
rect 4755 20757 4764 20791
rect 4712 20748 4764 20757
rect 7012 20748 7064 20800
rect 10968 20791 11020 20800
rect 10968 20757 10977 20791
rect 10977 20757 11011 20791
rect 11011 20757 11020 20791
rect 10968 20748 11020 20757
rect 12256 20791 12308 20800
rect 12256 20757 12265 20791
rect 12265 20757 12299 20791
rect 12299 20757 12308 20791
rect 12256 20748 12308 20757
rect 15568 20791 15620 20800
rect 15568 20757 15577 20791
rect 15577 20757 15611 20791
rect 15611 20757 15620 20791
rect 15568 20748 15620 20757
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 18144 20927 18196 20936
rect 18144 20893 18153 20927
rect 18153 20893 18187 20927
rect 18187 20893 18196 20927
rect 18144 20884 18196 20893
rect 19340 20884 19392 20936
rect 20076 20884 20128 20936
rect 21456 20884 21508 20936
rect 22468 20884 22520 20936
rect 25780 20927 25832 20936
rect 25780 20893 25789 20927
rect 25789 20893 25823 20927
rect 25823 20893 25832 20927
rect 25780 20884 25832 20893
rect 26976 20884 27028 20936
rect 28540 20884 28592 20936
rect 28724 20927 28776 20936
rect 28724 20893 28733 20927
rect 28733 20893 28767 20927
rect 28767 20893 28776 20927
rect 28724 20884 28776 20893
rect 28816 20927 28868 20936
rect 28816 20893 28825 20927
rect 28825 20893 28859 20927
rect 28859 20893 28868 20927
rect 28816 20884 28868 20893
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 18236 20816 18288 20868
rect 21824 20816 21876 20868
rect 26332 20816 26384 20868
rect 19064 20791 19116 20800
rect 19064 20757 19073 20791
rect 19073 20757 19107 20791
rect 19107 20757 19116 20791
rect 19064 20748 19116 20757
rect 23480 20748 23532 20800
rect 25320 20748 25372 20800
rect 25872 20748 25924 20800
rect 39212 20995 39264 21004
rect 39212 20961 39221 20995
rect 39221 20961 39255 20995
rect 39255 20961 39264 20995
rect 39212 20952 39264 20961
rect 39396 20995 39448 21004
rect 39396 20961 39405 20995
rect 39405 20961 39439 20995
rect 39439 20961 39448 20995
rect 39396 20952 39448 20961
rect 40040 20952 40092 21004
rect 40408 20995 40460 21004
rect 40408 20961 40417 20995
rect 40417 20961 40451 20995
rect 40451 20961 40460 20995
rect 40408 20952 40460 20961
rect 31116 20884 31168 20936
rect 31760 20884 31812 20936
rect 32128 20884 32180 20936
rect 33876 20884 33928 20936
rect 35992 20884 36044 20936
rect 36544 20927 36596 20936
rect 36544 20893 36553 20927
rect 36553 20893 36587 20927
rect 36587 20893 36596 20927
rect 36544 20884 36596 20893
rect 37188 20884 37240 20936
rect 37556 20927 37608 20936
rect 37556 20893 37590 20927
rect 37590 20893 37608 20927
rect 37556 20884 37608 20893
rect 27620 20748 27672 20800
rect 29092 20748 29144 20800
rect 34336 20816 34388 20868
rect 40408 20816 40460 20868
rect 40684 20859 40736 20868
rect 40684 20825 40693 20859
rect 40693 20825 40727 20859
rect 40727 20825 40736 20859
rect 40684 20816 40736 20825
rect 41236 20816 41288 20868
rect 31484 20748 31536 20800
rect 31852 20791 31904 20800
rect 31852 20757 31861 20791
rect 31861 20757 31895 20791
rect 31895 20757 31904 20791
rect 31852 20748 31904 20757
rect 32312 20748 32364 20800
rect 32496 20748 32548 20800
rect 32772 20748 32824 20800
rect 33692 20748 33744 20800
rect 34612 20748 34664 20800
rect 35624 20748 35676 20800
rect 38752 20791 38804 20800
rect 38752 20757 38761 20791
rect 38761 20757 38795 20791
rect 38795 20757 38804 20791
rect 38752 20748 38804 20757
rect 39580 20748 39632 20800
rect 42156 20791 42208 20800
rect 42156 20757 42165 20791
rect 42165 20757 42199 20791
rect 42199 20757 42208 20791
rect 42156 20748 42208 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 3148 20544 3200 20596
rect 4528 20587 4580 20596
rect 4528 20553 4537 20587
rect 4537 20553 4571 20587
rect 4571 20553 4580 20587
rect 4528 20544 4580 20553
rect 6276 20544 6328 20596
rect 9772 20587 9824 20596
rect 9772 20553 9781 20587
rect 9781 20553 9815 20587
rect 9815 20553 9824 20587
rect 9772 20544 9824 20553
rect 13176 20544 13228 20596
rect 18604 20544 18656 20596
rect 22284 20587 22336 20596
rect 22284 20553 22293 20587
rect 22293 20553 22327 20587
rect 22327 20553 22336 20587
rect 22284 20544 22336 20553
rect 25780 20544 25832 20596
rect 26332 20544 26384 20596
rect 27712 20544 27764 20596
rect 29000 20544 29052 20596
rect 32404 20544 32456 20596
rect 8392 20519 8444 20528
rect 8392 20485 8401 20519
rect 8401 20485 8435 20519
rect 8435 20485 8444 20519
rect 8392 20476 8444 20485
rect 12256 20476 12308 20528
rect 15568 20476 15620 20528
rect 19064 20476 19116 20528
rect 23480 20476 23532 20528
rect 25504 20476 25556 20528
rect 26056 20476 26108 20528
rect 29184 20476 29236 20528
rect 1676 20408 1728 20460
rect 1860 20451 1912 20460
rect 1860 20417 1894 20451
rect 1894 20417 1912 20451
rect 1860 20408 1912 20417
rect 3424 20451 3476 20460
rect 3424 20417 3433 20451
rect 3433 20417 3467 20451
rect 3467 20417 3476 20451
rect 3424 20408 3476 20417
rect 4620 20451 4672 20460
rect 4620 20417 4629 20451
rect 4629 20417 4663 20451
rect 4663 20417 4672 20451
rect 4620 20408 4672 20417
rect 5264 20408 5316 20460
rect 6552 20408 6604 20460
rect 8944 20408 8996 20460
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 9128 20408 9180 20417
rect 10968 20408 11020 20460
rect 11612 20408 11664 20460
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 20720 20408 20772 20460
rect 3332 20383 3384 20392
rect 3332 20349 3341 20383
rect 3341 20349 3375 20383
rect 3375 20349 3384 20383
rect 3332 20340 3384 20349
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 6276 20340 6328 20392
rect 8484 20340 8536 20392
rect 14464 20383 14516 20392
rect 14464 20349 14473 20383
rect 14473 20349 14507 20383
rect 14507 20349 14516 20383
rect 14464 20340 14516 20349
rect 16580 20340 16632 20392
rect 17316 20340 17368 20392
rect 17960 20340 18012 20392
rect 21088 20383 21140 20392
rect 21088 20349 21097 20383
rect 21097 20349 21131 20383
rect 21131 20349 21140 20383
rect 21088 20340 21140 20349
rect 22376 20383 22428 20392
rect 22376 20349 22385 20383
rect 22385 20349 22419 20383
rect 22419 20349 22428 20383
rect 22376 20340 22428 20349
rect 22468 20340 22520 20392
rect 25964 20451 26016 20460
rect 25964 20417 25973 20451
rect 25973 20417 26007 20451
rect 26007 20417 26016 20451
rect 25964 20408 26016 20417
rect 28356 20451 28408 20460
rect 28356 20417 28365 20451
rect 28365 20417 28399 20451
rect 28399 20417 28408 20451
rect 28356 20408 28408 20417
rect 40224 20587 40276 20596
rect 40224 20553 40233 20587
rect 40233 20553 40267 20587
rect 40267 20553 40276 20587
rect 40224 20544 40276 20553
rect 40684 20544 40736 20596
rect 41972 20544 42024 20596
rect 32772 20476 32824 20528
rect 33324 20476 33376 20528
rect 34796 20476 34848 20528
rect 37188 20476 37240 20528
rect 33140 20408 33192 20460
rect 34428 20408 34480 20460
rect 35348 20408 35400 20460
rect 39948 20476 40000 20528
rect 40500 20476 40552 20528
rect 38752 20408 38804 20460
rect 38844 20451 38896 20460
rect 38844 20417 38853 20451
rect 38853 20417 38887 20451
rect 38887 20417 38896 20451
rect 38844 20408 38896 20417
rect 25872 20340 25924 20392
rect 26976 20272 27028 20324
rect 27620 20272 27672 20324
rect 3056 20204 3108 20256
rect 3700 20204 3752 20256
rect 5264 20247 5316 20256
rect 5264 20213 5273 20247
rect 5273 20213 5307 20247
rect 5307 20213 5316 20247
rect 5264 20204 5316 20213
rect 6828 20204 6880 20256
rect 17132 20204 17184 20256
rect 20076 20247 20128 20256
rect 20076 20213 20085 20247
rect 20085 20213 20119 20247
rect 20119 20213 20128 20247
rect 20076 20204 20128 20213
rect 22008 20204 22060 20256
rect 26884 20204 26936 20256
rect 28080 20383 28132 20392
rect 28080 20349 28089 20383
rect 28089 20349 28123 20383
rect 28123 20349 28132 20383
rect 28080 20340 28132 20349
rect 29092 20340 29144 20392
rect 30104 20383 30156 20392
rect 30104 20349 30113 20383
rect 30113 20349 30147 20383
rect 30147 20349 30156 20383
rect 30104 20340 30156 20349
rect 32128 20340 32180 20392
rect 33508 20340 33560 20392
rect 29276 20204 29328 20256
rect 33876 20204 33928 20256
rect 33968 20247 34020 20256
rect 33968 20213 33977 20247
rect 33977 20213 34011 20247
rect 34011 20213 34020 20247
rect 33968 20204 34020 20213
rect 34152 20204 34204 20256
rect 36912 20383 36964 20392
rect 36912 20349 36921 20383
rect 36921 20349 36955 20383
rect 36955 20349 36964 20383
rect 36912 20340 36964 20349
rect 40960 20408 41012 20460
rect 41512 20451 41564 20460
rect 41512 20417 41521 20451
rect 41521 20417 41555 20451
rect 41555 20417 41564 20451
rect 41512 20408 41564 20417
rect 40408 20340 40460 20392
rect 41696 20383 41748 20392
rect 41696 20349 41705 20383
rect 41705 20349 41739 20383
rect 41739 20349 41748 20383
rect 41696 20340 41748 20349
rect 36176 20247 36228 20256
rect 36176 20213 36185 20247
rect 36185 20213 36219 20247
rect 36219 20213 36228 20247
rect 36176 20204 36228 20213
rect 39028 20204 39080 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3884 20000 3936 20052
rect 4712 20000 4764 20052
rect 6460 20000 6512 20052
rect 10048 20000 10100 20052
rect 11796 20000 11848 20052
rect 17316 20043 17368 20052
rect 17316 20009 17325 20043
rect 17325 20009 17359 20043
rect 17359 20009 17368 20043
rect 17316 20000 17368 20009
rect 19340 20000 19392 20052
rect 20536 20000 20588 20052
rect 6644 19932 6696 19984
rect 8392 19932 8444 19984
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 3240 19796 3292 19848
rect 3700 19796 3752 19848
rect 4160 19839 4212 19848
rect 4160 19805 4169 19839
rect 4169 19805 4203 19839
rect 4203 19805 4212 19839
rect 4160 19796 4212 19805
rect 6092 19864 6144 19916
rect 6828 19864 6880 19916
rect 10508 19975 10560 19984
rect 10508 19941 10517 19975
rect 10517 19941 10551 19975
rect 10551 19941 10560 19975
rect 10508 19932 10560 19941
rect 11612 19932 11664 19984
rect 3056 19728 3108 19780
rect 4344 19728 4396 19780
rect 8116 19839 8168 19848
rect 6368 19771 6420 19780
rect 6368 19737 6377 19771
rect 6377 19737 6411 19771
rect 6411 19737 6420 19771
rect 6368 19728 6420 19737
rect 6828 19728 6880 19780
rect 8116 19805 8125 19839
rect 8125 19805 8159 19839
rect 8159 19805 8168 19839
rect 8116 19796 8168 19805
rect 7104 19771 7156 19780
rect 7104 19737 7113 19771
rect 7113 19737 7147 19771
rect 7147 19737 7156 19771
rect 7104 19728 7156 19737
rect 4620 19660 4672 19712
rect 5908 19660 5960 19712
rect 6460 19660 6512 19712
rect 7012 19660 7064 19712
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 8484 19839 8536 19848
rect 8484 19805 8493 19839
rect 8493 19805 8527 19839
rect 8527 19805 8536 19839
rect 8484 19796 8536 19805
rect 8668 19796 8720 19848
rect 9772 19796 9824 19848
rect 10140 19796 10192 19848
rect 10968 19796 11020 19848
rect 11520 19839 11572 19848
rect 11520 19805 11529 19839
rect 11529 19805 11563 19839
rect 11563 19805 11572 19839
rect 11520 19796 11572 19805
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 18052 19864 18104 19916
rect 18604 19864 18656 19916
rect 13820 19796 13872 19848
rect 14464 19796 14516 19848
rect 9312 19728 9364 19780
rect 8852 19660 8904 19712
rect 9680 19660 9732 19712
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 10416 19660 10468 19669
rect 12072 19660 12124 19712
rect 12256 19771 12308 19780
rect 12256 19737 12290 19771
rect 12290 19737 12308 19771
rect 12256 19728 12308 19737
rect 15752 19771 15804 19780
rect 15752 19737 15761 19771
rect 15761 19737 15795 19771
rect 15795 19737 15804 19771
rect 15752 19728 15804 19737
rect 13176 19660 13228 19712
rect 16212 19728 16264 19780
rect 18420 19796 18472 19848
rect 20628 19864 20680 19916
rect 22008 19907 22060 19916
rect 22008 19873 22017 19907
rect 22017 19873 22051 19907
rect 22051 19873 22060 19907
rect 22008 19864 22060 19873
rect 18604 19728 18656 19780
rect 19800 19839 19852 19848
rect 19800 19805 19809 19839
rect 19809 19805 19843 19839
rect 19843 19805 19852 19839
rect 19800 19796 19852 19805
rect 29000 20000 29052 20052
rect 31944 20000 31996 20052
rect 33048 20000 33100 20052
rect 35348 20000 35400 20052
rect 37924 20000 37976 20052
rect 41696 20000 41748 20052
rect 28356 19864 28408 19916
rect 32864 19864 32916 19916
rect 33048 19907 33100 19916
rect 33048 19873 33057 19907
rect 33057 19873 33091 19907
rect 33091 19873 33100 19907
rect 33048 19864 33100 19873
rect 33876 19864 33928 19916
rect 20444 19728 20496 19780
rect 20720 19728 20772 19780
rect 23756 19796 23808 19848
rect 22468 19771 22520 19780
rect 22468 19737 22477 19771
rect 22477 19737 22511 19771
rect 22511 19737 22520 19771
rect 22468 19728 22520 19737
rect 26884 19771 26936 19780
rect 26884 19737 26893 19771
rect 26893 19737 26927 19771
rect 26927 19737 26936 19771
rect 26884 19728 26936 19737
rect 29000 19728 29052 19780
rect 29184 19728 29236 19780
rect 17224 19703 17276 19712
rect 17224 19669 17233 19703
rect 17233 19669 17267 19703
rect 17267 19669 17276 19703
rect 17224 19660 17276 19669
rect 17776 19703 17828 19712
rect 17776 19669 17785 19703
rect 17785 19669 17819 19703
rect 17819 19669 17828 19703
rect 17776 19660 17828 19669
rect 21088 19660 21140 19712
rect 21824 19660 21876 19712
rect 23480 19703 23532 19712
rect 23480 19669 23489 19703
rect 23489 19669 23523 19703
rect 23523 19669 23532 19703
rect 23480 19660 23532 19669
rect 23572 19660 23624 19712
rect 25044 19660 25096 19712
rect 25504 19660 25556 19712
rect 27712 19660 27764 19712
rect 29828 19660 29880 19712
rect 34428 19796 34480 19848
rect 34704 19839 34756 19848
rect 34704 19805 34713 19839
rect 34713 19805 34747 19839
rect 34747 19805 34756 19839
rect 34704 19796 34756 19805
rect 36176 19864 36228 19916
rect 36636 19796 36688 19848
rect 38844 19907 38896 19916
rect 38844 19873 38853 19907
rect 38853 19873 38887 19907
rect 38887 19873 38896 19907
rect 38844 19864 38896 19873
rect 39028 19839 39080 19848
rect 39028 19805 39037 19839
rect 39037 19805 39071 19839
rect 39071 19805 39080 19839
rect 39028 19796 39080 19805
rect 31760 19660 31812 19712
rect 36544 19771 36596 19780
rect 36544 19737 36553 19771
rect 36553 19737 36587 19771
rect 36587 19737 36596 19771
rect 36544 19728 36596 19737
rect 34428 19660 34480 19712
rect 36912 19660 36964 19712
rect 37188 19660 37240 19712
rect 38476 19728 38528 19780
rect 40224 19771 40276 19780
rect 40224 19737 40233 19771
rect 40233 19737 40267 19771
rect 40267 19737 40276 19771
rect 40224 19728 40276 19737
rect 41236 19728 41288 19780
rect 38660 19660 38712 19712
rect 39580 19703 39632 19712
rect 39580 19669 39589 19703
rect 39589 19669 39623 19703
rect 39623 19669 39632 19703
rect 39580 19660 39632 19669
rect 40868 19660 40920 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 1860 19456 1912 19508
rect 3056 19456 3108 19508
rect 8300 19456 8352 19508
rect 9128 19456 9180 19508
rect 10508 19456 10560 19508
rect 10876 19456 10928 19508
rect 12256 19456 12308 19508
rect 15752 19456 15804 19508
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 3240 19431 3292 19440
rect 3240 19397 3249 19431
rect 3249 19397 3283 19431
rect 3283 19397 3292 19431
rect 3240 19388 3292 19397
rect 4160 19388 4212 19440
rect 4896 19388 4948 19440
rect 4712 19320 4764 19372
rect 5908 19388 5960 19440
rect 5264 19320 5316 19372
rect 6644 19363 6696 19372
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 3332 19252 3384 19304
rect 4344 19252 4396 19304
rect 4620 19252 4672 19304
rect 5724 19295 5776 19304
rect 5724 19261 5733 19295
rect 5733 19261 5767 19295
rect 5767 19261 5776 19295
rect 5724 19252 5776 19261
rect 4804 19184 4856 19236
rect 6092 19252 6144 19304
rect 7196 19388 7248 19440
rect 8668 19431 8720 19440
rect 8668 19397 8677 19431
rect 8677 19397 8711 19431
rect 8711 19397 8720 19431
rect 8668 19388 8720 19397
rect 8852 19431 8904 19440
rect 8852 19397 8861 19431
rect 8861 19397 8895 19431
rect 8895 19397 8904 19431
rect 8852 19388 8904 19397
rect 6920 19363 6972 19372
rect 6920 19329 6954 19363
rect 6954 19329 6972 19363
rect 6920 19320 6972 19329
rect 8116 19320 8168 19372
rect 10416 19388 10468 19440
rect 10968 19388 11020 19440
rect 6828 19116 6880 19168
rect 8116 19116 8168 19168
rect 9680 19320 9732 19372
rect 9772 19363 9824 19372
rect 9772 19329 9781 19363
rect 9781 19329 9815 19363
rect 9815 19329 9824 19363
rect 9772 19320 9824 19329
rect 11796 19320 11848 19372
rect 17776 19456 17828 19508
rect 9220 19295 9272 19304
rect 9220 19261 9229 19295
rect 9229 19261 9263 19295
rect 9263 19261 9272 19295
rect 9220 19252 9272 19261
rect 9404 19295 9456 19304
rect 9404 19261 9413 19295
rect 9413 19261 9447 19295
rect 9447 19261 9456 19295
rect 9404 19252 9456 19261
rect 11336 19252 11388 19304
rect 11520 19252 11572 19304
rect 12072 19295 12124 19304
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 12072 19252 12124 19261
rect 12256 19363 12308 19372
rect 12256 19329 12265 19363
rect 12265 19329 12299 19363
rect 12299 19329 12308 19363
rect 12256 19320 12308 19329
rect 12532 19252 12584 19304
rect 13820 19320 13872 19372
rect 14372 19320 14424 19372
rect 17960 19388 18012 19440
rect 18420 19388 18472 19440
rect 20720 19388 20772 19440
rect 22468 19456 22520 19508
rect 25412 19456 25464 19508
rect 26792 19456 26844 19508
rect 23572 19388 23624 19440
rect 25504 19388 25556 19440
rect 13452 19252 13504 19304
rect 13176 19184 13228 19236
rect 9956 19116 10008 19168
rect 17684 19116 17736 19168
rect 18328 19252 18380 19304
rect 19248 19252 19300 19304
rect 20720 19252 20772 19304
rect 20904 19252 20956 19304
rect 22744 19252 22796 19304
rect 26332 19363 26384 19372
rect 26332 19329 26341 19363
rect 26341 19329 26375 19363
rect 26375 19329 26384 19363
rect 28632 19456 28684 19508
rect 29828 19456 29880 19508
rect 31576 19499 31628 19508
rect 31576 19465 31585 19499
rect 31585 19465 31619 19499
rect 31619 19465 31628 19499
rect 31576 19456 31628 19465
rect 32128 19499 32180 19508
rect 32128 19465 32137 19499
rect 32137 19465 32171 19499
rect 32171 19465 32180 19499
rect 32128 19456 32180 19465
rect 32588 19456 32640 19508
rect 29000 19388 29052 19440
rect 26332 19320 26384 19329
rect 23756 19227 23808 19236
rect 23756 19193 23765 19227
rect 23765 19193 23799 19227
rect 23799 19193 23808 19227
rect 23756 19184 23808 19193
rect 22376 19116 22428 19168
rect 24124 19295 24176 19304
rect 24124 19261 24133 19295
rect 24133 19261 24167 19295
rect 24167 19261 24176 19295
rect 24124 19252 24176 19261
rect 26516 19295 26568 19304
rect 26516 19261 26525 19295
rect 26525 19261 26559 19295
rect 26559 19261 26568 19295
rect 26516 19252 26568 19261
rect 26700 19252 26752 19304
rect 28264 19295 28316 19304
rect 28264 19261 28273 19295
rect 28273 19261 28307 19295
rect 28307 19261 28316 19295
rect 28264 19252 28316 19261
rect 29000 19252 29052 19304
rect 33140 19388 33192 19440
rect 29828 19363 29880 19372
rect 29828 19329 29837 19363
rect 29837 19329 29871 19363
rect 29871 19329 29880 19363
rect 29828 19320 29880 19329
rect 34704 19456 34756 19508
rect 36360 19456 36412 19508
rect 38476 19499 38528 19508
rect 38476 19465 38485 19499
rect 38485 19465 38519 19499
rect 38519 19465 38528 19499
rect 38476 19456 38528 19465
rect 40224 19499 40276 19508
rect 40224 19465 40233 19499
rect 40233 19465 40267 19499
rect 40267 19465 40276 19499
rect 40224 19456 40276 19465
rect 40960 19456 41012 19508
rect 41512 19499 41564 19508
rect 41512 19465 41521 19499
rect 41521 19465 41555 19499
rect 41555 19465 41564 19499
rect 41512 19456 41564 19465
rect 33968 19388 34020 19440
rect 34428 19431 34480 19440
rect 34428 19397 34437 19431
rect 34437 19397 34471 19431
rect 34471 19397 34480 19431
rect 34428 19388 34480 19397
rect 39580 19388 39632 19440
rect 29644 19252 29696 19304
rect 30472 19252 30524 19304
rect 34336 19252 34388 19304
rect 25228 19116 25280 19168
rect 25964 19159 26016 19168
rect 25964 19125 25973 19159
rect 25973 19125 26007 19159
rect 26007 19125 26016 19159
rect 25964 19116 26016 19125
rect 33232 19116 33284 19168
rect 34704 19252 34756 19304
rect 35348 19295 35400 19304
rect 35348 19261 35357 19295
rect 35357 19261 35391 19295
rect 35391 19261 35400 19295
rect 35348 19252 35400 19261
rect 38108 19363 38160 19372
rect 38108 19329 38117 19363
rect 38117 19329 38151 19363
rect 38151 19329 38160 19363
rect 38108 19320 38160 19329
rect 40592 19363 40644 19372
rect 40592 19329 40601 19363
rect 40601 19329 40635 19363
rect 40635 19329 40644 19363
rect 40592 19320 40644 19329
rect 40868 19320 40920 19372
rect 36544 19252 36596 19304
rect 37924 19295 37976 19304
rect 37924 19261 37933 19295
rect 37933 19261 37967 19295
rect 37967 19261 37976 19295
rect 37924 19252 37976 19261
rect 41052 19184 41104 19236
rect 42156 19295 42208 19304
rect 42156 19261 42165 19295
rect 42165 19261 42199 19295
rect 42199 19261 42208 19295
rect 42156 19252 42208 19261
rect 41328 19116 41380 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4712 18912 4764 18964
rect 5724 18912 5776 18964
rect 6368 18912 6420 18964
rect 6828 18955 6880 18964
rect 6828 18921 6837 18955
rect 6837 18921 6871 18955
rect 6871 18921 6880 18955
rect 6828 18912 6880 18921
rect 3976 18844 4028 18896
rect 6920 18844 6972 18896
rect 7012 18844 7064 18896
rect 3700 18708 3752 18760
rect 3976 18708 4028 18760
rect 4804 18708 4856 18760
rect 7748 18683 7800 18692
rect 7748 18649 7757 18683
rect 7757 18649 7791 18683
rect 7791 18649 7800 18683
rect 7748 18640 7800 18649
rect 8484 18776 8536 18828
rect 9680 18844 9732 18896
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 10784 18912 10836 18964
rect 12256 18912 12308 18964
rect 17776 18912 17828 18964
rect 18328 18955 18380 18964
rect 18328 18921 18337 18955
rect 18337 18921 18371 18955
rect 18371 18921 18380 18955
rect 18328 18912 18380 18921
rect 18420 18912 18472 18964
rect 20720 18955 20772 18964
rect 20720 18921 20729 18955
rect 20729 18921 20763 18955
rect 20763 18921 20772 18955
rect 20720 18912 20772 18921
rect 22744 18955 22796 18964
rect 22744 18921 22753 18955
rect 22753 18921 22787 18955
rect 22787 18921 22796 18955
rect 22744 18912 22796 18921
rect 24124 18912 24176 18964
rect 24952 18912 25004 18964
rect 26700 18955 26752 18964
rect 26700 18921 26709 18955
rect 26709 18921 26743 18955
rect 26743 18921 26752 18955
rect 26700 18912 26752 18921
rect 28264 18912 28316 18964
rect 30472 18955 30524 18964
rect 30472 18921 30481 18955
rect 30481 18921 30515 18955
rect 30515 18921 30524 18955
rect 30472 18912 30524 18921
rect 33600 18912 33652 18964
rect 10508 18776 10560 18828
rect 8392 18751 8444 18760
rect 8392 18717 8401 18751
rect 8401 18717 8435 18751
rect 8435 18717 8444 18751
rect 8392 18708 8444 18717
rect 9220 18708 9272 18760
rect 10048 18708 10100 18760
rect 10876 18751 10928 18760
rect 10876 18717 10885 18751
rect 10885 18717 10919 18751
rect 10919 18717 10928 18751
rect 10876 18708 10928 18717
rect 4896 18572 4948 18624
rect 8668 18640 8720 18692
rect 9956 18683 10008 18692
rect 9956 18649 9965 18683
rect 9965 18649 9999 18683
rect 9999 18649 10008 18683
rect 9956 18640 10008 18649
rect 7932 18572 7984 18624
rect 9404 18572 9456 18624
rect 9864 18615 9916 18624
rect 9864 18581 9873 18615
rect 9873 18581 9907 18615
rect 9907 18581 9916 18615
rect 10784 18640 10836 18692
rect 11336 18683 11388 18692
rect 11336 18649 11345 18683
rect 11345 18649 11379 18683
rect 11379 18649 11388 18683
rect 11336 18640 11388 18649
rect 12072 18751 12124 18760
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 12532 18819 12584 18828
rect 12532 18785 12541 18819
rect 12541 18785 12575 18819
rect 12575 18785 12584 18819
rect 12532 18776 12584 18785
rect 12532 18640 12584 18692
rect 9864 18572 9916 18581
rect 10232 18572 10284 18624
rect 12716 18751 12768 18760
rect 12716 18717 12726 18751
rect 12726 18717 12760 18751
rect 12760 18717 12768 18751
rect 12716 18708 12768 18717
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13636 18751 13688 18760
rect 13636 18717 13645 18751
rect 13645 18717 13679 18751
rect 13679 18717 13688 18751
rect 13636 18708 13688 18717
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 18052 18776 18104 18828
rect 19248 18708 19300 18760
rect 20904 18708 20956 18760
rect 13084 18640 13136 18692
rect 13176 18683 13228 18692
rect 13176 18649 13185 18683
rect 13185 18649 13219 18683
rect 13219 18649 13228 18683
rect 13176 18640 13228 18649
rect 19708 18683 19760 18692
rect 19708 18649 19717 18683
rect 19717 18649 19751 18683
rect 19751 18649 19760 18683
rect 19708 18640 19760 18649
rect 19800 18640 19852 18692
rect 23204 18819 23256 18828
rect 23204 18785 23213 18819
rect 23213 18785 23247 18819
rect 23247 18785 23256 18819
rect 23204 18776 23256 18785
rect 23388 18708 23440 18760
rect 28080 18776 28132 18828
rect 31024 18819 31076 18828
rect 31024 18785 31033 18819
rect 31033 18785 31067 18819
rect 31067 18785 31076 18819
rect 31024 18776 31076 18785
rect 33324 18776 33376 18828
rect 25228 18708 25280 18760
rect 25964 18708 26016 18760
rect 29644 18708 29696 18760
rect 31576 18708 31628 18760
rect 31760 18708 31812 18760
rect 32588 18751 32640 18760
rect 32588 18717 32597 18751
rect 32597 18717 32631 18751
rect 32631 18717 32640 18751
rect 32588 18708 32640 18717
rect 36544 18912 36596 18964
rect 38108 18912 38160 18964
rect 40592 18912 40644 18964
rect 42064 18844 42116 18896
rect 34704 18776 34756 18828
rect 37188 18776 37240 18828
rect 39304 18751 39356 18760
rect 39304 18717 39313 18751
rect 39313 18717 39347 18751
rect 39347 18717 39356 18751
rect 39304 18708 39356 18717
rect 24400 18640 24452 18692
rect 33140 18640 33192 18692
rect 14188 18572 14240 18624
rect 19340 18572 19392 18624
rect 21456 18572 21508 18624
rect 25412 18572 25464 18624
rect 28908 18615 28960 18624
rect 28908 18581 28917 18615
rect 28917 18581 28951 18615
rect 28951 18581 28960 18615
rect 28908 18572 28960 18581
rect 30932 18615 30984 18624
rect 30932 18581 30941 18615
rect 30941 18581 30975 18615
rect 30975 18581 30984 18615
rect 30932 18572 30984 18581
rect 36544 18640 36596 18692
rect 40868 18708 40920 18760
rect 41604 18708 41656 18760
rect 41052 18640 41104 18692
rect 35440 18572 35492 18624
rect 36084 18572 36136 18624
rect 37924 18572 37976 18624
rect 40224 18572 40276 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 8392 18368 8444 18420
rect 10140 18368 10192 18420
rect 11612 18368 11664 18420
rect 9864 18343 9916 18352
rect 9864 18309 9873 18343
rect 9873 18309 9907 18343
rect 9907 18309 9916 18343
rect 9864 18300 9916 18309
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 8484 18232 8536 18284
rect 9220 18275 9272 18284
rect 9220 18241 9229 18275
rect 9229 18241 9263 18275
rect 9263 18241 9272 18275
rect 9220 18232 9272 18241
rect 9680 18232 9732 18284
rect 10048 18275 10100 18284
rect 10048 18241 10057 18275
rect 10057 18241 10091 18275
rect 10091 18241 10100 18275
rect 10048 18232 10100 18241
rect 8852 18207 8904 18216
rect 8852 18173 8861 18207
rect 8861 18173 8895 18207
rect 8895 18173 8904 18207
rect 8852 18164 8904 18173
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 12532 18300 12584 18352
rect 14188 18343 14240 18352
rect 14188 18309 14206 18343
rect 14206 18309 14240 18343
rect 14188 18300 14240 18309
rect 18420 18300 18472 18352
rect 19984 18368 20036 18420
rect 20812 18368 20864 18420
rect 26332 18411 26384 18420
rect 26332 18377 26341 18411
rect 26341 18377 26375 18411
rect 26375 18377 26384 18411
rect 26332 18368 26384 18377
rect 20352 18300 20404 18352
rect 25044 18300 25096 18352
rect 31944 18368 31996 18420
rect 33140 18368 33192 18420
rect 33600 18368 33652 18420
rect 35348 18368 35400 18420
rect 36360 18368 36412 18420
rect 38660 18368 38712 18420
rect 29092 18300 29144 18352
rect 32588 18300 32640 18352
rect 37924 18300 37976 18352
rect 13176 18232 13228 18284
rect 14372 18232 14424 18284
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 17960 18232 18012 18284
rect 19708 18232 19760 18284
rect 28632 18232 28684 18284
rect 31576 18232 31628 18284
rect 32404 18232 32456 18284
rect 34520 18232 34572 18284
rect 40224 18300 40276 18352
rect 41052 18368 41104 18420
rect 42064 18300 42116 18352
rect 42248 18300 42300 18352
rect 6368 18096 6420 18148
rect 8116 18096 8168 18148
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 4804 18028 4856 18080
rect 7380 18028 7432 18080
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 12532 18207 12584 18216
rect 12532 18173 12541 18207
rect 12541 18173 12575 18207
rect 12575 18173 12584 18207
rect 12532 18164 12584 18173
rect 12808 18164 12860 18216
rect 17408 18164 17460 18216
rect 18420 18207 18472 18216
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 22192 18164 22244 18216
rect 24308 18164 24360 18216
rect 24952 18164 25004 18216
rect 27528 18207 27580 18216
rect 27528 18173 27537 18207
rect 27537 18173 27571 18207
rect 27571 18173 27580 18207
rect 27528 18164 27580 18173
rect 29000 18207 29052 18216
rect 29000 18173 29009 18207
rect 29009 18173 29043 18207
rect 29043 18173 29052 18207
rect 29000 18164 29052 18173
rect 31024 18164 31076 18216
rect 36452 18207 36504 18216
rect 36452 18173 36461 18207
rect 36461 18173 36495 18207
rect 36495 18173 36504 18207
rect 36452 18164 36504 18173
rect 37464 18164 37516 18216
rect 20904 18096 20956 18148
rect 34796 18096 34848 18148
rect 35992 18096 36044 18148
rect 12808 18028 12860 18080
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 25504 18028 25556 18080
rect 30472 18071 30524 18080
rect 30472 18037 30481 18071
rect 30481 18037 30515 18071
rect 30515 18037 30524 18071
rect 30472 18028 30524 18037
rect 30748 18028 30800 18080
rect 35532 18028 35584 18080
rect 36360 18028 36412 18080
rect 37188 18028 37240 18080
rect 37832 18207 37884 18216
rect 37832 18173 37841 18207
rect 37841 18173 37875 18207
rect 37875 18173 37884 18207
rect 37832 18164 37884 18173
rect 41328 18164 41380 18216
rect 39304 18071 39356 18080
rect 39304 18037 39313 18071
rect 39313 18037 39347 18071
rect 39347 18037 39356 18071
rect 39304 18028 39356 18037
rect 41420 18028 41472 18080
rect 41696 18071 41748 18080
rect 41696 18037 41705 18071
rect 41705 18037 41739 18071
rect 41739 18037 41748 18071
rect 41696 18028 41748 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 5816 17824 5868 17876
rect 10876 17867 10928 17876
rect 10876 17833 10885 17867
rect 10885 17833 10919 17867
rect 10919 17833 10928 17867
rect 10876 17824 10928 17833
rect 18420 17824 18472 17876
rect 23756 17824 23808 17876
rect 24400 17867 24452 17876
rect 24400 17833 24409 17867
rect 24409 17833 24443 17867
rect 24443 17833 24452 17867
rect 24400 17824 24452 17833
rect 26516 17824 26568 17876
rect 27528 17824 27580 17876
rect 35440 17824 35492 17876
rect 41604 17867 41656 17876
rect 41604 17833 41613 17867
rect 41613 17833 41647 17867
rect 41647 17833 41656 17867
rect 41604 17824 41656 17833
rect 4620 17756 4672 17808
rect 5172 17756 5224 17808
rect 5908 17756 5960 17808
rect 6000 17756 6052 17808
rect 1584 17688 1636 17740
rect 5448 17688 5500 17740
rect 5540 17688 5592 17740
rect 1676 17620 1728 17672
rect 4712 17620 4764 17672
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 2780 17552 2832 17604
rect 4804 17552 4856 17604
rect 6000 17663 6052 17672
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 10232 17731 10284 17740
rect 10232 17697 10241 17731
rect 10241 17697 10275 17731
rect 10275 17697 10284 17731
rect 10232 17688 10284 17697
rect 12532 17731 12584 17740
rect 12532 17697 12541 17731
rect 12541 17697 12575 17731
rect 12575 17697 12584 17731
rect 12532 17688 12584 17697
rect 12808 17731 12860 17740
rect 12808 17697 12817 17731
rect 12817 17697 12851 17731
rect 12851 17697 12860 17731
rect 12808 17688 12860 17697
rect 17040 17688 17092 17740
rect 7656 17620 7708 17672
rect 10140 17620 10192 17672
rect 10508 17620 10560 17672
rect 3056 17484 3108 17536
rect 6552 17552 6604 17604
rect 7472 17552 7524 17604
rect 9772 17552 9824 17604
rect 6092 17484 6144 17536
rect 8852 17484 8904 17536
rect 9404 17484 9456 17536
rect 9864 17527 9916 17536
rect 9864 17493 9873 17527
rect 9873 17493 9907 17527
rect 9907 17493 9916 17527
rect 9864 17484 9916 17493
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 16672 17620 16724 17672
rect 17684 17731 17736 17740
rect 17684 17697 17693 17731
rect 17693 17697 17727 17731
rect 17727 17697 17736 17731
rect 17684 17688 17736 17697
rect 18328 17688 18380 17740
rect 22008 17756 22060 17808
rect 19708 17688 19760 17740
rect 19892 17688 19944 17740
rect 24952 17731 25004 17740
rect 24952 17697 24961 17731
rect 24961 17697 24995 17731
rect 24995 17697 25004 17731
rect 24952 17688 25004 17697
rect 25228 17731 25280 17740
rect 25228 17697 25237 17731
rect 25237 17697 25271 17731
rect 25271 17697 25280 17731
rect 25228 17688 25280 17697
rect 25504 17731 25556 17740
rect 25504 17697 25513 17731
rect 25513 17697 25547 17731
rect 25547 17697 25556 17731
rect 25504 17688 25556 17697
rect 19984 17620 20036 17672
rect 22468 17663 22520 17672
rect 22468 17629 22477 17663
rect 22477 17629 22511 17663
rect 22511 17629 22520 17663
rect 22468 17620 22520 17629
rect 30196 17688 30248 17740
rect 12348 17595 12400 17604
rect 12348 17561 12366 17595
rect 12366 17561 12400 17595
rect 12348 17552 12400 17561
rect 13912 17552 13964 17604
rect 20904 17595 20956 17604
rect 20904 17561 20913 17595
rect 20913 17561 20947 17595
rect 20947 17561 20956 17595
rect 20904 17552 20956 17561
rect 12716 17484 12768 17536
rect 13544 17484 13596 17536
rect 17040 17527 17092 17536
rect 17040 17493 17049 17527
rect 17049 17493 17083 17527
rect 17083 17493 17092 17527
rect 17040 17484 17092 17493
rect 17408 17527 17460 17536
rect 17408 17493 17417 17527
rect 17417 17493 17451 17527
rect 17451 17493 17460 17527
rect 17408 17484 17460 17493
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 22744 17595 22796 17604
rect 22744 17561 22753 17595
rect 22753 17561 22787 17595
rect 22787 17561 22796 17595
rect 22744 17552 22796 17561
rect 25044 17552 25096 17604
rect 27344 17595 27396 17604
rect 27344 17561 27353 17595
rect 27353 17561 27387 17595
rect 27387 17561 27396 17595
rect 27344 17552 27396 17561
rect 29092 17552 29144 17604
rect 30472 17620 30524 17672
rect 31760 17688 31812 17740
rect 33324 17756 33376 17808
rect 35072 17756 35124 17808
rect 36452 17688 36504 17740
rect 39580 17756 39632 17808
rect 31116 17595 31168 17604
rect 31116 17561 31125 17595
rect 31125 17561 31159 17595
rect 31159 17561 31168 17595
rect 31116 17552 31168 17561
rect 27620 17484 27672 17536
rect 28724 17484 28776 17536
rect 29460 17484 29512 17536
rect 29736 17484 29788 17536
rect 30196 17484 30248 17536
rect 30656 17484 30708 17536
rect 33508 17620 33560 17672
rect 34520 17620 34572 17672
rect 34796 17620 34848 17672
rect 34980 17620 35032 17672
rect 37004 17620 37056 17672
rect 37464 17620 37516 17672
rect 39948 17688 40000 17740
rect 41052 17688 41104 17740
rect 39856 17620 39908 17672
rect 41420 17620 41472 17672
rect 33784 17552 33836 17604
rect 34704 17552 34756 17604
rect 35532 17595 35584 17604
rect 35532 17561 35541 17595
rect 35541 17561 35575 17595
rect 35575 17561 35584 17595
rect 35532 17552 35584 17561
rect 36084 17595 36136 17604
rect 36084 17561 36093 17595
rect 36093 17561 36127 17595
rect 36127 17561 36136 17595
rect 36084 17552 36136 17561
rect 38016 17552 38068 17604
rect 38660 17552 38712 17604
rect 33508 17527 33560 17536
rect 33508 17493 33517 17527
rect 33517 17493 33551 17527
rect 33551 17493 33560 17527
rect 33508 17484 33560 17493
rect 34520 17484 34572 17536
rect 35440 17484 35492 17536
rect 38844 17484 38896 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 4804 17280 4856 17332
rect 5264 17280 5316 17332
rect 848 17144 900 17196
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 3976 17144 4028 17196
rect 4988 17212 5040 17264
rect 6000 17280 6052 17332
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 10600 17280 10652 17332
rect 12440 17280 12492 17332
rect 12808 17280 12860 17332
rect 4896 17187 4948 17196
rect 4896 17153 4905 17187
rect 4905 17153 4939 17187
rect 4939 17153 4948 17187
rect 4896 17144 4948 17153
rect 5264 17144 5316 17196
rect 12348 17212 12400 17264
rect 17408 17280 17460 17332
rect 22468 17280 22520 17332
rect 1768 17076 1820 17128
rect 5172 17076 5224 17128
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6092 17144 6144 17196
rect 6552 17144 6604 17196
rect 5632 17119 5684 17128
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 6368 17119 6420 17128
rect 6368 17085 6377 17119
rect 6377 17085 6411 17119
rect 6411 17085 6420 17119
rect 6368 17076 6420 17085
rect 6736 17144 6788 17196
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 7932 17144 7984 17196
rect 8116 17187 8168 17196
rect 8116 17153 8150 17187
rect 8150 17153 8168 17187
rect 8116 17144 8168 17153
rect 9404 17187 9456 17196
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 7656 17076 7708 17128
rect 9956 17144 10008 17196
rect 11428 17144 11480 17196
rect 11060 17076 11112 17128
rect 12624 17144 12676 17196
rect 20812 17212 20864 17264
rect 23756 17255 23808 17264
rect 23756 17221 23765 17255
rect 23765 17221 23799 17255
rect 23799 17221 23808 17255
rect 23756 17212 23808 17221
rect 13268 17144 13320 17196
rect 19892 17187 19944 17196
rect 19892 17153 19901 17187
rect 19901 17153 19935 17187
rect 19935 17153 19944 17187
rect 19892 17144 19944 17153
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 12532 17076 12584 17128
rect 12808 17076 12860 17128
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 18144 17119 18196 17128
rect 18144 17085 18153 17119
rect 18153 17085 18187 17119
rect 18187 17085 18196 17119
rect 18144 17076 18196 17085
rect 20812 17076 20864 17128
rect 12992 17008 13044 17060
rect 22100 17008 22152 17060
rect 22744 17008 22796 17060
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 4620 16983 4672 16992
rect 4620 16949 4629 16983
rect 4629 16949 4663 16983
rect 4663 16949 4672 16983
rect 4620 16940 4672 16949
rect 5448 16940 5500 16992
rect 5908 16940 5960 16992
rect 6552 16940 6604 16992
rect 9220 16983 9272 16992
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 9404 16940 9456 16992
rect 10324 16940 10376 16992
rect 10508 16940 10560 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 21364 16940 21416 16992
rect 22560 16940 22612 16992
rect 23848 17187 23900 17196
rect 23848 17153 23857 17187
rect 23857 17153 23891 17187
rect 23891 17153 23900 17187
rect 23848 17144 23900 17153
rect 25228 17280 25280 17332
rect 27344 17280 27396 17332
rect 29000 17280 29052 17332
rect 24400 17255 24452 17264
rect 24400 17221 24409 17255
rect 24409 17221 24443 17255
rect 24443 17221 24452 17255
rect 24400 17212 24452 17221
rect 25044 17212 25096 17264
rect 24492 17076 24544 17128
rect 28908 17212 28960 17264
rect 27436 17187 27488 17196
rect 27436 17153 27445 17187
rect 27445 17153 27479 17187
rect 27479 17153 27488 17187
rect 27436 17144 27488 17153
rect 27712 17144 27764 17196
rect 28080 17187 28132 17196
rect 28080 17153 28089 17187
rect 28089 17153 28123 17187
rect 28123 17153 28132 17187
rect 28080 17144 28132 17153
rect 28172 17187 28224 17196
rect 28172 17153 28181 17187
rect 28181 17153 28215 17187
rect 28215 17153 28224 17187
rect 28172 17144 28224 17153
rect 28724 17187 28776 17196
rect 28724 17153 28733 17187
rect 28733 17153 28767 17187
rect 28767 17153 28776 17187
rect 28724 17144 28776 17153
rect 29736 17255 29788 17264
rect 29736 17221 29745 17255
rect 29745 17221 29779 17255
rect 29779 17221 29788 17255
rect 29736 17212 29788 17221
rect 30656 17255 30708 17264
rect 30656 17221 30665 17255
rect 30665 17221 30699 17255
rect 30699 17221 30708 17255
rect 30656 17212 30708 17221
rect 31116 17323 31168 17332
rect 31116 17289 31125 17323
rect 31125 17289 31159 17323
rect 31159 17289 31168 17323
rect 31116 17280 31168 17289
rect 32036 17212 32088 17264
rect 29644 17187 29696 17196
rect 29644 17153 29653 17187
rect 29653 17153 29687 17187
rect 29687 17153 29696 17187
rect 29644 17144 29696 17153
rect 26056 17076 26108 17128
rect 25504 17008 25556 17060
rect 29000 17076 29052 17128
rect 30196 17187 30248 17196
rect 30196 17153 30205 17187
rect 30205 17153 30239 17187
rect 30239 17153 30248 17187
rect 30196 17144 30248 17153
rect 30564 17144 30616 17196
rect 30748 17187 30800 17196
rect 30748 17153 30757 17187
rect 30757 17153 30791 17187
rect 30791 17153 30800 17187
rect 30748 17144 30800 17153
rect 30380 17076 30432 17128
rect 31944 17144 31996 17196
rect 34428 17255 34480 17264
rect 34428 17221 34437 17255
rect 34437 17221 34471 17255
rect 34471 17221 34480 17255
rect 34428 17212 34480 17221
rect 37832 17280 37884 17332
rect 38016 17280 38068 17332
rect 36544 17212 36596 17264
rect 33232 17187 33284 17196
rect 33232 17153 33241 17187
rect 33241 17153 33275 17187
rect 33275 17153 33284 17187
rect 33232 17144 33284 17153
rect 33600 17187 33652 17196
rect 33600 17153 33609 17187
rect 33609 17153 33643 17187
rect 33643 17153 33652 17187
rect 33600 17144 33652 17153
rect 33784 17187 33836 17196
rect 33784 17153 33793 17187
rect 33793 17153 33827 17187
rect 33827 17153 33836 17187
rect 33784 17144 33836 17153
rect 33508 17119 33560 17128
rect 25412 16940 25464 16992
rect 33508 17085 33517 17119
rect 33517 17085 33551 17119
rect 33551 17085 33560 17119
rect 33508 17076 33560 17085
rect 34520 17187 34572 17196
rect 34520 17153 34529 17187
rect 34529 17153 34563 17187
rect 34563 17153 34572 17187
rect 34520 17144 34572 17153
rect 34796 17187 34848 17196
rect 34796 17153 34805 17187
rect 34805 17153 34839 17187
rect 34839 17153 34848 17187
rect 34796 17144 34848 17153
rect 34980 17187 35032 17196
rect 34980 17153 34989 17187
rect 34989 17153 35023 17187
rect 35023 17153 35032 17187
rect 34980 17144 35032 17153
rect 31852 17008 31904 17060
rect 27804 16983 27856 16992
rect 27804 16949 27813 16983
rect 27813 16949 27847 16983
rect 27847 16949 27856 16983
rect 27804 16940 27856 16949
rect 30288 16940 30340 16992
rect 32496 16983 32548 16992
rect 32496 16949 32505 16983
rect 32505 16949 32539 16983
rect 32539 16949 32548 16983
rect 32496 16940 32548 16949
rect 33324 16983 33376 16992
rect 33324 16949 33333 16983
rect 33333 16949 33367 16983
rect 33367 16949 33376 16983
rect 33324 16940 33376 16949
rect 34060 16940 34112 16992
rect 34520 17008 34572 17060
rect 35072 17076 35124 17128
rect 38016 17144 38068 17196
rect 35256 17119 35308 17128
rect 35256 17085 35265 17119
rect 35265 17085 35299 17119
rect 35299 17085 35308 17119
rect 35256 17076 35308 17085
rect 35716 16940 35768 16992
rect 37004 16983 37056 16992
rect 37004 16949 37013 16983
rect 37013 16949 37047 16983
rect 37047 16949 37056 16983
rect 37004 16940 37056 16949
rect 37556 17119 37608 17128
rect 37556 17085 37565 17119
rect 37565 17085 37599 17119
rect 37599 17085 37608 17119
rect 37556 17076 37608 17085
rect 37924 17076 37976 17128
rect 38844 17255 38896 17264
rect 38844 17221 38853 17255
rect 38853 17221 38887 17255
rect 38887 17221 38896 17255
rect 38844 17212 38896 17221
rect 40040 17280 40092 17332
rect 40132 17280 40184 17332
rect 38476 17187 38528 17196
rect 38476 17153 38485 17187
rect 38485 17153 38519 17187
rect 38519 17153 38528 17187
rect 38476 17144 38528 17153
rect 38568 17144 38620 17196
rect 38476 17008 38528 17060
rect 39580 17187 39632 17196
rect 39580 17153 39589 17187
rect 39589 17153 39623 17187
rect 39623 17153 39632 17187
rect 39580 17144 39632 17153
rect 39856 17187 39908 17196
rect 39856 17153 39865 17187
rect 39865 17153 39899 17187
rect 39899 17153 39908 17187
rect 39856 17144 39908 17153
rect 39948 17187 40000 17196
rect 39948 17153 39957 17187
rect 39957 17153 39991 17187
rect 39991 17153 40000 17187
rect 39948 17144 40000 17153
rect 41972 17144 42024 17196
rect 42156 17144 42208 17196
rect 41696 17008 41748 17060
rect 39580 16940 39632 16992
rect 40408 16940 40460 16992
rect 40500 16940 40552 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 5632 16736 5684 16788
rect 6000 16736 6052 16788
rect 6552 16736 6604 16788
rect 8116 16736 8168 16788
rect 4896 16668 4948 16720
rect 1584 16600 1636 16652
rect 5264 16643 5316 16652
rect 5264 16609 5273 16643
rect 5273 16609 5307 16643
rect 5307 16609 5316 16643
rect 5264 16600 5316 16609
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 5908 16668 5960 16720
rect 10876 16736 10928 16788
rect 11428 16779 11480 16788
rect 11428 16745 11437 16779
rect 11437 16745 11471 16779
rect 11471 16745 11480 16779
rect 11428 16736 11480 16745
rect 6184 16600 6236 16652
rect 1676 16532 1728 16584
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 11060 16668 11112 16720
rect 9956 16600 10008 16652
rect 4804 16532 4856 16541
rect 2780 16464 2832 16516
rect 3976 16464 4028 16516
rect 4896 16507 4948 16516
rect 4896 16473 4905 16507
rect 4905 16473 4939 16507
rect 4939 16473 4948 16507
rect 4896 16464 4948 16473
rect 5172 16464 5224 16516
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 8668 16464 8720 16516
rect 8852 16464 8904 16516
rect 9404 16575 9456 16584
rect 9404 16541 9413 16575
rect 9413 16541 9447 16575
rect 9447 16541 9456 16575
rect 9404 16532 9456 16541
rect 12348 16736 12400 16788
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 12900 16736 12952 16788
rect 13268 16779 13320 16788
rect 13268 16745 13277 16779
rect 13277 16745 13311 16779
rect 13311 16745 13320 16779
rect 13268 16736 13320 16745
rect 13912 16779 13964 16788
rect 13912 16745 13921 16779
rect 13921 16745 13955 16779
rect 13955 16745 13964 16779
rect 13912 16736 13964 16745
rect 20812 16779 20864 16788
rect 20812 16745 20821 16779
rect 20821 16745 20855 16779
rect 20855 16745 20864 16779
rect 20812 16736 20864 16745
rect 23848 16736 23900 16788
rect 24400 16779 24452 16788
rect 24400 16745 24409 16779
rect 24409 16745 24443 16779
rect 24443 16745 24452 16779
rect 24400 16736 24452 16745
rect 24768 16736 24820 16788
rect 28080 16736 28132 16788
rect 29092 16736 29144 16788
rect 30288 16736 30340 16788
rect 32496 16736 32548 16788
rect 17040 16668 17092 16720
rect 13636 16643 13688 16652
rect 9680 16464 9732 16516
rect 10324 16464 10376 16516
rect 11980 16464 12032 16516
rect 2964 16396 3016 16448
rect 5632 16396 5684 16448
rect 11888 16396 11940 16448
rect 12440 16507 12492 16516
rect 12440 16473 12449 16507
rect 12449 16473 12483 16507
rect 12483 16473 12492 16507
rect 12440 16464 12492 16473
rect 12624 16507 12676 16516
rect 12624 16473 12665 16507
rect 12665 16473 12676 16507
rect 13636 16609 13645 16643
rect 13645 16609 13679 16643
rect 13679 16609 13688 16643
rect 13636 16600 13688 16609
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 15200 16532 15252 16584
rect 15476 16532 15528 16584
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 18144 16532 18196 16584
rect 18696 16575 18748 16584
rect 12624 16464 12676 16473
rect 12900 16507 12952 16516
rect 12900 16473 12909 16507
rect 12909 16473 12943 16507
rect 12943 16473 12952 16507
rect 12900 16464 12952 16473
rect 12992 16464 13044 16516
rect 15384 16464 15436 16516
rect 16212 16464 16264 16516
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 18972 16532 19024 16584
rect 19708 16532 19760 16584
rect 19800 16575 19852 16584
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 12808 16396 12860 16448
rect 19524 16507 19576 16516
rect 19524 16473 19533 16507
rect 19533 16473 19567 16507
rect 19567 16473 19576 16507
rect 19524 16464 19576 16473
rect 19892 16464 19944 16516
rect 20260 16532 20312 16584
rect 20720 16532 20772 16584
rect 18144 16439 18196 16448
rect 18144 16405 18153 16439
rect 18153 16405 18187 16439
rect 18187 16405 18196 16439
rect 18144 16396 18196 16405
rect 18420 16439 18472 16448
rect 18420 16405 18429 16439
rect 18429 16405 18463 16439
rect 18463 16405 18472 16439
rect 18420 16396 18472 16405
rect 18788 16396 18840 16448
rect 19156 16396 19208 16448
rect 20628 16396 20680 16448
rect 21180 16507 21232 16516
rect 21180 16473 21189 16507
rect 21189 16473 21223 16507
rect 21223 16473 21232 16507
rect 21180 16464 21232 16473
rect 21456 16575 21508 16584
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 22100 16643 22152 16652
rect 22100 16609 22109 16643
rect 22109 16609 22143 16643
rect 22143 16609 22152 16643
rect 22100 16600 22152 16609
rect 21732 16532 21784 16584
rect 24124 16643 24176 16652
rect 24124 16609 24133 16643
rect 24133 16609 24167 16643
rect 24167 16609 24176 16643
rect 24124 16600 24176 16609
rect 25872 16668 25924 16720
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 22928 16532 22980 16584
rect 24216 16532 24268 16584
rect 24952 16532 25004 16584
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 25504 16532 25556 16541
rect 25596 16532 25648 16584
rect 26056 16575 26108 16584
rect 26056 16541 26065 16575
rect 26065 16541 26099 16575
rect 26099 16541 26108 16575
rect 26056 16532 26108 16541
rect 26884 16600 26936 16652
rect 27988 16668 28040 16720
rect 28172 16668 28224 16720
rect 28540 16532 28592 16584
rect 22836 16464 22888 16516
rect 26148 16464 26200 16516
rect 29460 16532 29512 16584
rect 30196 16600 30248 16652
rect 33508 16668 33560 16720
rect 34796 16779 34848 16788
rect 34796 16745 34805 16779
rect 34805 16745 34839 16779
rect 34839 16745 34848 16779
rect 34796 16736 34848 16745
rect 34888 16736 34940 16788
rect 38016 16736 38068 16788
rect 38568 16736 38620 16788
rect 31760 16600 31812 16652
rect 31944 16600 31996 16652
rect 33324 16600 33376 16652
rect 34888 16600 34940 16652
rect 37464 16600 37516 16652
rect 31392 16507 31444 16516
rect 31392 16473 31401 16507
rect 31401 16473 31435 16507
rect 31435 16473 31444 16507
rect 31392 16464 31444 16473
rect 31760 16507 31812 16516
rect 31760 16473 31769 16507
rect 31769 16473 31803 16507
rect 31803 16473 31812 16507
rect 31760 16464 31812 16473
rect 32036 16464 32088 16516
rect 22100 16396 22152 16448
rect 22192 16439 22244 16448
rect 22192 16405 22201 16439
rect 22201 16405 22235 16439
rect 22235 16405 22244 16439
rect 22192 16396 22244 16405
rect 25044 16396 25096 16448
rect 27252 16396 27304 16448
rect 29368 16396 29420 16448
rect 30380 16396 30432 16448
rect 32220 16439 32272 16448
rect 32220 16405 32229 16439
rect 32229 16405 32263 16439
rect 32263 16405 32272 16439
rect 32220 16396 32272 16405
rect 34060 16575 34112 16584
rect 34060 16541 34069 16575
rect 34069 16541 34103 16575
rect 34103 16541 34112 16575
rect 34060 16532 34112 16541
rect 34980 16532 35032 16584
rect 35256 16532 35308 16584
rect 33232 16464 33284 16516
rect 33784 16439 33836 16448
rect 33784 16405 33793 16439
rect 33793 16405 33827 16439
rect 33827 16405 33836 16439
rect 33784 16396 33836 16405
rect 34060 16396 34112 16448
rect 34796 16464 34848 16516
rect 35164 16464 35216 16516
rect 35716 16532 35768 16584
rect 36360 16575 36412 16584
rect 36360 16541 36369 16575
rect 36369 16541 36403 16575
rect 36403 16541 36412 16575
rect 36360 16532 36412 16541
rect 35440 16464 35492 16516
rect 37004 16532 37056 16584
rect 37372 16532 37424 16584
rect 38200 16532 38252 16584
rect 34704 16396 34756 16448
rect 37556 16396 37608 16448
rect 39120 16396 39172 16448
rect 40500 16643 40552 16652
rect 40500 16609 40509 16643
rect 40509 16609 40543 16643
rect 40543 16609 40552 16643
rect 40500 16600 40552 16609
rect 40132 16575 40184 16584
rect 40132 16541 40141 16575
rect 40141 16541 40175 16575
rect 40175 16541 40184 16575
rect 40132 16532 40184 16541
rect 41604 16532 41656 16584
rect 40500 16464 40552 16516
rect 40040 16396 40092 16448
rect 41972 16439 42024 16448
rect 41972 16405 41981 16439
rect 41981 16405 42015 16439
rect 42015 16405 42024 16439
rect 41972 16396 42024 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 6368 16192 6420 16244
rect 8484 16192 8536 16244
rect 8852 16192 8904 16244
rect 12072 16192 12124 16244
rect 12900 16192 12952 16244
rect 13636 16192 13688 16244
rect 15660 16235 15712 16244
rect 15660 16201 15669 16235
rect 15669 16201 15703 16235
rect 15703 16201 15712 16235
rect 15660 16192 15712 16201
rect 18236 16192 18288 16244
rect 3976 16124 4028 16176
rect 5540 16124 5592 16176
rect 8208 16124 8260 16176
rect 9956 16124 10008 16176
rect 11980 16124 12032 16176
rect 12624 16124 12676 16176
rect 848 16056 900 16108
rect 2964 16099 3016 16108
rect 2964 16065 2973 16099
rect 2973 16065 3007 16099
rect 3007 16065 3016 16099
rect 2964 16056 3016 16065
rect 5356 16099 5408 16108
rect 5356 16065 5365 16099
rect 5365 16065 5399 16099
rect 5399 16065 5408 16099
rect 5356 16056 5408 16065
rect 6000 16056 6052 16108
rect 6092 16099 6144 16108
rect 6092 16065 6101 16099
rect 6101 16065 6135 16099
rect 6135 16065 6144 16099
rect 6092 16056 6144 16065
rect 1768 15988 1820 16040
rect 11060 15988 11112 16040
rect 5356 15920 5408 15972
rect 7748 15920 7800 15972
rect 11704 15920 11756 15972
rect 11888 16031 11940 16040
rect 11888 15997 11897 16031
rect 11897 15997 11931 16031
rect 11931 15997 11940 16031
rect 11888 15988 11940 15997
rect 11980 16031 12032 16040
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 1676 15852 1728 15904
rect 9404 15852 9456 15904
rect 10692 15852 10744 15904
rect 11612 15852 11664 15904
rect 12440 15920 12492 15972
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 20904 16192 20956 16244
rect 21180 16192 21232 16244
rect 24124 16235 24176 16244
rect 24124 16201 24133 16235
rect 24133 16201 24167 16235
rect 24167 16201 24176 16235
rect 24124 16192 24176 16201
rect 24216 16235 24268 16244
rect 24216 16201 24225 16235
rect 24225 16201 24259 16235
rect 24259 16201 24268 16235
rect 24216 16192 24268 16201
rect 24860 16192 24912 16244
rect 25596 16192 25648 16244
rect 29000 16192 29052 16244
rect 29368 16235 29420 16244
rect 29368 16201 29377 16235
rect 29377 16201 29411 16235
rect 29411 16201 29420 16235
rect 29368 16192 29420 16201
rect 30932 16192 30984 16244
rect 12716 16056 12768 16065
rect 13268 16056 13320 16108
rect 13820 16056 13872 16108
rect 15384 16056 15436 16108
rect 13360 15920 13412 15972
rect 15200 15920 15252 15972
rect 15844 16056 15896 16108
rect 16488 16031 16540 16040
rect 16488 15997 16497 16031
rect 16497 15997 16531 16031
rect 16531 15997 16540 16031
rect 16488 15988 16540 15997
rect 17132 16099 17184 16108
rect 17132 16065 17141 16099
rect 17141 16065 17175 16099
rect 17175 16065 17184 16099
rect 17132 16056 17184 16065
rect 19708 16124 19760 16176
rect 20812 16124 20864 16176
rect 23756 16167 23808 16176
rect 23756 16133 23765 16167
rect 23765 16133 23799 16167
rect 23799 16133 23808 16167
rect 23756 16124 23808 16133
rect 19432 16056 19484 16108
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 17316 16031 17368 16040
rect 17316 15997 17325 16031
rect 17325 15997 17359 16031
rect 17359 15997 17368 16031
rect 17316 15988 17368 15997
rect 17408 15988 17460 16040
rect 20168 15988 20220 16040
rect 21824 16099 21876 16108
rect 21824 16065 21833 16099
rect 21833 16065 21867 16099
rect 21867 16065 21876 16099
rect 21824 16056 21876 16065
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 23940 16099 23992 16108
rect 23940 16065 23949 16099
rect 23949 16065 23983 16099
rect 23983 16065 23992 16099
rect 23940 16056 23992 16065
rect 27252 16167 27304 16176
rect 27252 16133 27261 16167
rect 27261 16133 27295 16167
rect 27295 16133 27304 16167
rect 27252 16124 27304 16133
rect 29092 16124 29144 16176
rect 31392 16192 31444 16244
rect 34704 16192 34756 16244
rect 32220 16124 32272 16176
rect 33784 16167 33836 16176
rect 33784 16133 33793 16167
rect 33793 16133 33827 16167
rect 33827 16133 33836 16167
rect 33784 16124 33836 16133
rect 35256 16235 35308 16244
rect 35256 16201 35265 16235
rect 35265 16201 35299 16235
rect 35299 16201 35308 16235
rect 35256 16192 35308 16201
rect 37740 16235 37792 16244
rect 37740 16201 37749 16235
rect 37749 16201 37783 16235
rect 37783 16201 37792 16235
rect 37740 16192 37792 16201
rect 25044 16099 25096 16108
rect 25044 16065 25053 16099
rect 25053 16065 25087 16099
rect 25087 16065 25096 16099
rect 25044 16056 25096 16065
rect 30380 16056 30432 16108
rect 12808 15852 12860 15904
rect 12992 15852 13044 15904
rect 15384 15852 15436 15904
rect 15844 15895 15896 15904
rect 15844 15861 15853 15895
rect 15853 15861 15887 15895
rect 15887 15861 15896 15895
rect 15844 15852 15896 15861
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 17316 15852 17368 15904
rect 18144 15852 18196 15904
rect 20260 15852 20312 15904
rect 22192 15988 22244 16040
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 20904 15920 20956 15972
rect 21364 15963 21416 15972
rect 21364 15929 21373 15963
rect 21373 15929 21407 15963
rect 21407 15929 21416 15963
rect 21364 15920 21416 15929
rect 25044 15920 25096 15972
rect 20720 15852 20772 15904
rect 22100 15852 22152 15904
rect 22928 15852 22980 15904
rect 26792 15920 26844 15972
rect 26424 15852 26476 15904
rect 27804 15988 27856 16040
rect 28724 15988 28776 16040
rect 28632 15920 28684 15972
rect 29276 16031 29328 16040
rect 29276 15997 29285 16031
rect 29285 15997 29319 16031
rect 29319 15997 29328 16031
rect 29276 15988 29328 15997
rect 27620 15852 27672 15904
rect 28540 15852 28592 15904
rect 28816 15895 28868 15904
rect 28816 15861 28825 15895
rect 28825 15861 28859 15895
rect 28859 15861 28868 15895
rect 28816 15852 28868 15861
rect 31668 16056 31720 16108
rect 31944 16056 31996 16108
rect 35256 16056 35308 16108
rect 37464 16124 37516 16176
rect 36360 16056 36412 16108
rect 33876 15988 33928 16040
rect 34428 15988 34480 16040
rect 35164 15988 35216 16040
rect 40040 16099 40092 16108
rect 40040 16065 40048 16099
rect 40048 16065 40082 16099
rect 40082 16065 40092 16099
rect 40040 16056 40092 16065
rect 40132 16099 40184 16108
rect 40132 16065 40141 16099
rect 40141 16065 40175 16099
rect 40175 16065 40184 16099
rect 40132 16056 40184 16065
rect 41328 16056 41380 16108
rect 41972 16124 42024 16176
rect 42064 16056 42116 16108
rect 34980 15920 35032 15972
rect 37004 15920 37056 15972
rect 39488 16031 39540 16040
rect 39488 15997 39497 16031
rect 39497 15997 39531 16031
rect 39531 15997 39540 16031
rect 39488 15988 39540 15997
rect 38108 15920 38160 15972
rect 40224 16031 40276 16040
rect 40224 15997 40233 16031
rect 40233 15997 40267 16031
rect 40267 15997 40276 16031
rect 40224 15988 40276 15997
rect 40500 16031 40552 16040
rect 40500 15997 40509 16031
rect 40509 15997 40543 16031
rect 40543 15997 40552 16031
rect 40500 15988 40552 15997
rect 42248 15988 42300 16040
rect 35256 15852 35308 15904
rect 36544 15852 36596 15904
rect 37280 15895 37332 15904
rect 37280 15861 37289 15895
rect 37289 15861 37323 15895
rect 37323 15861 37332 15895
rect 37280 15852 37332 15861
rect 37556 15852 37608 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4804 15648 4856 15700
rect 5724 15691 5776 15700
rect 5724 15657 5733 15691
rect 5733 15657 5767 15691
rect 5767 15657 5776 15691
rect 5724 15648 5776 15657
rect 6460 15648 6512 15700
rect 8208 15648 8260 15700
rect 1768 15555 1820 15564
rect 1768 15521 1777 15555
rect 1777 15521 1811 15555
rect 1811 15521 1820 15555
rect 1768 15512 1820 15521
rect 5356 15555 5408 15564
rect 5356 15521 5365 15555
rect 5365 15521 5399 15555
rect 5399 15521 5408 15555
rect 5356 15512 5408 15521
rect 9036 15580 9088 15632
rect 9128 15580 9180 15632
rect 11612 15648 11664 15700
rect 11796 15648 11848 15700
rect 11980 15648 12032 15700
rect 13820 15691 13872 15700
rect 13820 15657 13829 15691
rect 13829 15657 13863 15691
rect 13863 15657 13872 15691
rect 13820 15648 13872 15657
rect 17500 15648 17552 15700
rect 18420 15648 18472 15700
rect 18880 15691 18932 15700
rect 18880 15657 18889 15691
rect 18889 15657 18923 15691
rect 18923 15657 18932 15691
rect 18880 15648 18932 15657
rect 19432 15648 19484 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 20352 15648 20404 15700
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2228 15444 2280 15496
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 7564 15444 7616 15496
rect 8208 15444 8260 15496
rect 3976 15376 4028 15428
rect 6644 15376 6696 15428
rect 7932 15419 7984 15428
rect 7932 15385 7941 15419
rect 7941 15385 7975 15419
rect 7975 15385 7984 15419
rect 7932 15376 7984 15385
rect 9588 15444 9640 15496
rect 9956 15512 10008 15564
rect 10692 15623 10744 15632
rect 10692 15589 10701 15623
rect 10701 15589 10735 15623
rect 10735 15589 10744 15623
rect 10692 15580 10744 15589
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 8484 15308 8536 15360
rect 12808 15444 12860 15496
rect 12992 15444 13044 15496
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 19156 15580 19208 15632
rect 19248 15580 19300 15632
rect 18696 15512 18748 15564
rect 13636 15487 13688 15496
rect 13636 15453 13645 15487
rect 13645 15453 13679 15487
rect 13679 15453 13688 15487
rect 13636 15444 13688 15453
rect 15200 15444 15252 15496
rect 12624 15308 12676 15360
rect 13544 15376 13596 15428
rect 16672 15376 16724 15428
rect 18236 15444 18288 15496
rect 18788 15487 18840 15496
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 19064 15555 19116 15564
rect 19064 15521 19073 15555
rect 19073 15521 19107 15555
rect 19107 15521 19116 15555
rect 19064 15512 19116 15521
rect 20812 15691 20864 15700
rect 20812 15657 20821 15691
rect 20821 15657 20855 15691
rect 20855 15657 20864 15691
rect 20812 15648 20864 15657
rect 20904 15648 20956 15700
rect 22192 15580 22244 15632
rect 21364 15512 21416 15564
rect 17040 15376 17092 15428
rect 17408 15376 17460 15428
rect 18972 15376 19024 15428
rect 20536 15376 20588 15428
rect 14372 15308 14424 15360
rect 18880 15308 18932 15360
rect 19892 15308 19944 15360
rect 20444 15308 20496 15360
rect 21824 15487 21876 15496
rect 21824 15453 21863 15487
rect 21863 15453 21876 15487
rect 21824 15444 21876 15453
rect 22284 15444 22336 15496
rect 22468 15580 22520 15632
rect 24768 15580 24820 15632
rect 22468 15444 22520 15496
rect 23756 15512 23808 15564
rect 26332 15580 26384 15632
rect 28540 15648 28592 15700
rect 27436 15580 27488 15632
rect 29276 15580 29328 15632
rect 23664 15444 23716 15496
rect 23940 15444 23992 15496
rect 25044 15487 25096 15496
rect 25044 15453 25053 15487
rect 25053 15453 25087 15487
rect 25087 15453 25096 15487
rect 25044 15444 25096 15453
rect 26056 15512 26108 15564
rect 26516 15512 26568 15564
rect 20996 15308 21048 15360
rect 22192 15308 22244 15360
rect 22284 15308 22336 15360
rect 23940 15308 23992 15360
rect 25596 15351 25648 15360
rect 25596 15317 25605 15351
rect 25605 15317 25639 15351
rect 25639 15317 25648 15351
rect 25596 15308 25648 15317
rect 26056 15376 26108 15428
rect 26332 15419 26384 15428
rect 26332 15385 26341 15419
rect 26341 15385 26375 15419
rect 26375 15385 26384 15419
rect 26332 15376 26384 15385
rect 26516 15419 26568 15428
rect 26516 15385 26525 15419
rect 26525 15385 26559 15419
rect 26559 15385 26568 15419
rect 26516 15376 26568 15385
rect 27252 15419 27304 15428
rect 27252 15385 27261 15419
rect 27261 15385 27295 15419
rect 27295 15385 27304 15419
rect 27252 15376 27304 15385
rect 27620 15487 27672 15496
rect 27620 15453 27629 15487
rect 27629 15453 27663 15487
rect 27663 15453 27672 15487
rect 27620 15444 27672 15453
rect 28632 15487 28684 15496
rect 28632 15453 28641 15487
rect 28641 15453 28675 15487
rect 28675 15453 28684 15487
rect 28632 15444 28684 15453
rect 29460 15512 29512 15564
rect 37096 15648 37148 15700
rect 37280 15648 37332 15700
rect 38660 15648 38712 15700
rect 41604 15691 41656 15700
rect 41604 15657 41613 15691
rect 41613 15657 41647 15691
rect 41647 15657 41656 15691
rect 41604 15648 41656 15657
rect 31300 15512 31352 15564
rect 33048 15512 33100 15564
rect 35256 15555 35308 15564
rect 35256 15521 35265 15555
rect 35265 15521 35299 15555
rect 35299 15521 35308 15555
rect 35256 15512 35308 15521
rect 37464 15512 37516 15564
rect 38660 15512 38712 15564
rect 27712 15376 27764 15428
rect 29736 15487 29788 15496
rect 29736 15453 29745 15487
rect 29745 15453 29779 15487
rect 29779 15453 29788 15487
rect 29736 15444 29788 15453
rect 31760 15444 31812 15496
rect 31852 15487 31904 15496
rect 31852 15453 31861 15487
rect 31861 15453 31895 15487
rect 31895 15453 31904 15487
rect 31852 15444 31904 15453
rect 32772 15376 32824 15428
rect 35440 15376 35492 15428
rect 26700 15308 26752 15360
rect 26792 15308 26844 15360
rect 27528 15308 27580 15360
rect 28356 15308 28408 15360
rect 29736 15308 29788 15360
rect 31024 15351 31076 15360
rect 31024 15317 31033 15351
rect 31033 15317 31067 15351
rect 31067 15317 31076 15351
rect 31024 15308 31076 15317
rect 36544 15308 36596 15360
rect 39488 15512 39540 15564
rect 39856 15512 39908 15564
rect 39120 15487 39172 15496
rect 39120 15453 39129 15487
rect 39129 15453 39163 15487
rect 39163 15453 39172 15487
rect 39120 15444 39172 15453
rect 39580 15487 39632 15496
rect 39580 15453 39589 15487
rect 39589 15453 39623 15487
rect 39623 15453 39632 15487
rect 39580 15444 39632 15453
rect 39028 15376 39080 15428
rect 40040 15487 40092 15496
rect 40040 15453 40049 15487
rect 40049 15453 40083 15487
rect 40083 15453 40092 15487
rect 40040 15444 40092 15453
rect 40408 15487 40460 15496
rect 40408 15453 40417 15487
rect 40417 15453 40451 15487
rect 40451 15453 40460 15487
rect 40408 15444 40460 15453
rect 39212 15351 39264 15360
rect 39212 15317 39221 15351
rect 39221 15317 39255 15351
rect 39255 15317 39264 15351
rect 39212 15308 39264 15317
rect 39304 15351 39356 15360
rect 39304 15317 39313 15351
rect 39313 15317 39347 15351
rect 39347 15317 39356 15351
rect 39304 15308 39356 15317
rect 40040 15308 40092 15360
rect 41420 15487 41472 15496
rect 41420 15453 41429 15487
rect 41429 15453 41463 15487
rect 41463 15453 41472 15487
rect 41420 15444 41472 15453
rect 41788 15376 41840 15428
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 4620 15104 4672 15156
rect 5172 15104 5224 15156
rect 5540 15104 5592 15156
rect 7104 15104 7156 15156
rect 7932 15104 7984 15156
rect 10048 15104 10100 15156
rect 3976 15036 4028 15088
rect 5264 15036 5316 15088
rect 5724 15036 5776 15088
rect 8300 15036 8352 15088
rect 13544 15147 13596 15156
rect 13544 15113 13553 15147
rect 13553 15113 13587 15147
rect 13587 15113 13596 15147
rect 13544 15104 13596 15113
rect 16488 15147 16540 15156
rect 16488 15113 16497 15147
rect 16497 15113 16531 15147
rect 16531 15113 16540 15147
rect 16488 15104 16540 15113
rect 18144 15147 18196 15156
rect 18144 15113 18153 15147
rect 18153 15113 18187 15147
rect 18187 15113 18196 15147
rect 18144 15104 18196 15113
rect 19064 15147 19116 15156
rect 19064 15113 19073 15147
rect 19073 15113 19107 15147
rect 19107 15113 19116 15147
rect 19064 15104 19116 15113
rect 19340 15104 19392 15156
rect 19708 15104 19760 15156
rect 19984 15104 20036 15156
rect 20904 15104 20956 15156
rect 2688 14943 2740 14952
rect 2688 14909 2697 14943
rect 2697 14909 2731 14943
rect 2731 14909 2740 14943
rect 2688 14900 2740 14909
rect 3792 14900 3844 14952
rect 5908 14968 5960 15020
rect 5816 14900 5868 14952
rect 5724 14832 5776 14884
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 8484 14968 8536 15020
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 15200 14968 15252 15020
rect 15384 15011 15436 15020
rect 15384 14977 15418 15011
rect 15418 14977 15436 15011
rect 15384 14968 15436 14977
rect 16580 14968 16632 15020
rect 17960 14968 18012 15020
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 10324 14900 10376 14952
rect 12992 14900 13044 14952
rect 17040 14900 17092 14952
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 18420 14900 18472 14952
rect 19892 15011 19944 15020
rect 19892 14977 19901 15011
rect 19901 14977 19935 15011
rect 19935 14977 19944 15011
rect 19892 14968 19944 14977
rect 20352 15079 20404 15088
rect 20352 15045 20361 15079
rect 20361 15045 20395 15079
rect 20395 15045 20404 15079
rect 20352 15036 20404 15045
rect 20444 15036 20496 15088
rect 20628 15036 20680 15088
rect 22836 15036 22888 15088
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 22284 15011 22336 15020
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 29092 15104 29144 15156
rect 29460 15104 29512 15156
rect 31668 15104 31720 15156
rect 31852 15147 31904 15156
rect 31852 15113 31861 15147
rect 31861 15113 31895 15147
rect 31895 15113 31904 15147
rect 31852 15104 31904 15113
rect 32772 15147 32824 15156
rect 32772 15113 32781 15147
rect 32781 15113 32815 15147
rect 32815 15113 32824 15147
rect 32772 15104 32824 15113
rect 26240 15079 26292 15088
rect 26240 15045 26249 15079
rect 26249 15045 26283 15079
rect 26283 15045 26292 15079
rect 26240 15036 26292 15045
rect 20444 14900 20496 14952
rect 22192 14900 22244 14952
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 5448 14807 5500 14816
rect 5448 14773 5457 14807
rect 5457 14773 5491 14807
rect 5491 14773 5500 14807
rect 5448 14764 5500 14773
rect 6276 14764 6328 14816
rect 12348 14832 12400 14884
rect 18788 14832 18840 14884
rect 10048 14807 10100 14816
rect 10048 14773 10057 14807
rect 10057 14773 10091 14807
rect 10091 14773 10100 14807
rect 10048 14764 10100 14773
rect 16212 14764 16264 14816
rect 18880 14764 18932 14816
rect 19248 14764 19300 14816
rect 21640 14832 21692 14884
rect 24492 14900 24544 14952
rect 25872 14968 25924 15020
rect 26424 15011 26476 15020
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 26424 14968 26476 14977
rect 27620 15036 27672 15088
rect 25320 14900 25372 14952
rect 25596 14900 25648 14952
rect 27436 15011 27488 15020
rect 27436 14977 27445 15011
rect 27445 14977 27479 15011
rect 27479 14977 27488 15011
rect 27436 14968 27488 14977
rect 28816 14968 28868 15020
rect 29092 15011 29144 15020
rect 29092 14977 29101 15011
rect 29101 14977 29135 15011
rect 29135 14977 29144 15011
rect 29092 14968 29144 14977
rect 28172 14900 28224 14952
rect 28724 14943 28776 14952
rect 28724 14909 28733 14943
rect 28733 14909 28767 14943
rect 28767 14909 28776 14943
rect 28724 14900 28776 14909
rect 21456 14764 21508 14816
rect 21732 14764 21784 14816
rect 26424 14832 26476 14884
rect 26792 14832 26844 14884
rect 28540 14832 28592 14884
rect 29368 15011 29420 15020
rect 29368 14977 29377 15011
rect 29377 14977 29411 15011
rect 29411 14977 29420 15011
rect 29368 14968 29420 14977
rect 31024 15036 31076 15088
rect 34428 15036 34480 15088
rect 29828 14832 29880 14884
rect 33140 14900 33192 14952
rect 33876 14943 33928 14952
rect 33876 14909 33885 14943
rect 33885 14909 33919 14943
rect 33919 14909 33928 14943
rect 33876 14900 33928 14909
rect 30472 14832 30524 14884
rect 31576 14832 31628 14884
rect 34520 14968 34572 15020
rect 35440 15104 35492 15156
rect 37096 15104 37148 15156
rect 37464 15104 37516 15156
rect 38016 15036 38068 15088
rect 38752 15036 38804 15088
rect 39212 15036 39264 15088
rect 39856 15036 39908 15088
rect 37280 14968 37332 15020
rect 37464 15011 37516 15020
rect 37464 14977 37473 15011
rect 37473 14977 37507 15011
rect 37507 14977 37516 15011
rect 37464 14968 37516 14977
rect 41420 15104 41472 15156
rect 35440 14900 35492 14952
rect 23112 14764 23164 14816
rect 24124 14764 24176 14816
rect 25872 14764 25924 14816
rect 26240 14764 26292 14816
rect 27252 14764 27304 14816
rect 32220 14764 32272 14816
rect 34060 14764 34112 14816
rect 35348 14832 35400 14884
rect 36544 14943 36596 14952
rect 36544 14909 36553 14943
rect 36553 14909 36587 14943
rect 36587 14909 36596 14943
rect 36544 14900 36596 14909
rect 37740 14943 37792 14952
rect 37740 14909 37749 14943
rect 37749 14909 37783 14943
rect 37783 14909 37792 14943
rect 37740 14900 37792 14909
rect 40868 14900 40920 14952
rect 41604 14900 41656 14952
rect 36452 14764 36504 14816
rect 40132 14832 40184 14884
rect 38476 14764 38528 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3792 14603 3844 14612
rect 3792 14569 3801 14603
rect 3801 14569 3835 14603
rect 3835 14569 3844 14603
rect 3792 14560 3844 14569
rect 4896 14560 4948 14612
rect 10324 14603 10376 14612
rect 10324 14569 10333 14603
rect 10333 14569 10367 14603
rect 10367 14569 10376 14603
rect 10324 14560 10376 14569
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 22376 14560 22428 14612
rect 28632 14560 28684 14612
rect 37740 14560 37792 14612
rect 39580 14603 39632 14612
rect 39580 14569 39589 14603
rect 39589 14569 39623 14603
rect 39623 14569 39632 14603
rect 39580 14560 39632 14569
rect 40868 14603 40920 14612
rect 40868 14569 40877 14603
rect 40877 14569 40911 14603
rect 40911 14569 40920 14603
rect 40868 14560 40920 14569
rect 41788 14603 41840 14612
rect 41788 14569 41797 14603
rect 41797 14569 41831 14603
rect 41831 14569 41840 14603
rect 41788 14560 41840 14569
rect 18328 14492 18380 14544
rect 19432 14492 19484 14544
rect 20260 14492 20312 14544
rect 2688 14424 2740 14476
rect 1676 14356 1728 14408
rect 7564 14424 7616 14476
rect 8300 14424 8352 14476
rect 12164 14424 12216 14476
rect 16948 14424 17000 14476
rect 20536 14467 20588 14476
rect 9036 14356 9088 14408
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 11980 14356 12032 14408
rect 18788 14356 18840 14408
rect 20536 14433 20545 14467
rect 20545 14433 20579 14467
rect 20579 14433 20588 14467
rect 20536 14424 20588 14433
rect 19708 14399 19760 14408
rect 19708 14365 19743 14399
rect 19743 14365 19760 14399
rect 19708 14356 19760 14365
rect 20720 14356 20772 14408
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 21732 14492 21784 14544
rect 35440 14492 35492 14544
rect 27620 14424 27672 14476
rect 29828 14467 29880 14476
rect 29828 14433 29837 14467
rect 29837 14433 29871 14467
rect 29871 14433 29880 14467
rect 29828 14424 29880 14433
rect 29920 14424 29972 14476
rect 2780 14288 2832 14340
rect 3976 14288 4028 14340
rect 4620 14288 4672 14340
rect 9864 14288 9916 14340
rect 16212 14331 16264 14340
rect 16212 14297 16221 14331
rect 16221 14297 16255 14331
rect 16255 14297 16264 14331
rect 16212 14288 16264 14297
rect 18512 14288 18564 14340
rect 19156 14288 19208 14340
rect 20260 14288 20312 14340
rect 21456 14331 21508 14340
rect 21456 14297 21465 14331
rect 21465 14297 21499 14331
rect 21499 14297 21508 14331
rect 21456 14288 21508 14297
rect 26792 14399 26844 14408
rect 26792 14365 26801 14399
rect 26801 14365 26835 14399
rect 26835 14365 26844 14399
rect 26792 14356 26844 14365
rect 31944 14467 31996 14476
rect 31944 14433 31953 14467
rect 31953 14433 31987 14467
rect 31987 14433 31996 14467
rect 31944 14424 31996 14433
rect 32220 14467 32272 14476
rect 32220 14433 32229 14467
rect 32229 14433 32263 14467
rect 32263 14433 32272 14467
rect 32220 14424 32272 14433
rect 38108 14424 38160 14476
rect 22100 14288 22152 14340
rect 22836 14288 22888 14340
rect 23756 14288 23808 14340
rect 25320 14288 25372 14340
rect 6000 14220 6052 14272
rect 11704 14220 11756 14272
rect 12808 14220 12860 14272
rect 17960 14220 18012 14272
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 21088 14263 21140 14272
rect 21088 14229 21097 14263
rect 21097 14229 21131 14263
rect 21131 14229 21140 14263
rect 21088 14220 21140 14229
rect 24768 14220 24820 14272
rect 26516 14288 26568 14340
rect 26884 14288 26936 14340
rect 26700 14263 26752 14272
rect 26700 14229 26709 14263
rect 26709 14229 26743 14263
rect 26743 14229 26752 14263
rect 26700 14220 26752 14229
rect 34336 14356 34388 14408
rect 35164 14399 35216 14408
rect 35164 14365 35173 14399
rect 35173 14365 35207 14399
rect 35207 14365 35216 14399
rect 35164 14356 35216 14365
rect 38384 14399 38436 14408
rect 38384 14365 38393 14399
rect 38393 14365 38427 14399
rect 38427 14365 38436 14399
rect 38384 14356 38436 14365
rect 38476 14399 38528 14408
rect 38476 14365 38511 14399
rect 38511 14365 38528 14399
rect 38476 14356 38528 14365
rect 38660 14399 38712 14408
rect 38660 14365 38669 14399
rect 38669 14365 38703 14399
rect 38703 14365 38712 14399
rect 38660 14356 38712 14365
rect 28356 14220 28408 14272
rect 29092 14288 29144 14340
rect 30380 14288 30432 14340
rect 31852 14331 31904 14340
rect 31852 14297 31861 14331
rect 31861 14297 31895 14331
rect 31895 14297 31904 14331
rect 31852 14288 31904 14297
rect 32956 14288 33008 14340
rect 34428 14288 34480 14340
rect 39120 14399 39172 14408
rect 39120 14365 39129 14399
rect 39129 14365 39163 14399
rect 39163 14365 39172 14399
rect 39120 14356 39172 14365
rect 39212 14356 39264 14408
rect 39580 14424 39632 14476
rect 39488 14399 39540 14408
rect 39488 14365 39497 14399
rect 39497 14365 39531 14399
rect 39531 14365 39540 14399
rect 39488 14356 39540 14365
rect 39764 14356 39816 14408
rect 39856 14399 39908 14408
rect 39856 14365 39865 14399
rect 39865 14365 39899 14399
rect 39899 14365 39908 14399
rect 39856 14356 39908 14365
rect 40040 14424 40092 14476
rect 41512 14399 41564 14408
rect 41512 14365 41521 14399
rect 41521 14365 41555 14399
rect 41555 14365 41564 14399
rect 41512 14356 41564 14365
rect 28816 14220 28868 14272
rect 29276 14220 29328 14272
rect 30564 14220 30616 14272
rect 33876 14220 33928 14272
rect 34612 14220 34664 14272
rect 35348 14220 35400 14272
rect 37924 14220 37976 14272
rect 38384 14220 38436 14272
rect 39120 14220 39172 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 2228 14016 2280 14068
rect 4804 14016 4856 14068
rect 5632 14016 5684 14068
rect 11704 14059 11756 14068
rect 4620 13948 4672 14000
rect 4712 13948 4764 14000
rect 5356 13948 5408 14000
rect 6000 13991 6052 14000
rect 6000 13957 6009 13991
rect 6009 13957 6043 13991
rect 6043 13957 6052 13991
rect 6000 13948 6052 13957
rect 6092 13948 6144 14000
rect 6552 13948 6604 14000
rect 9864 13991 9916 14000
rect 9864 13957 9873 13991
rect 9873 13957 9907 13991
rect 9907 13957 9916 13991
rect 9864 13948 9916 13957
rect 10324 13948 10376 14000
rect 5632 13880 5684 13932
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 3332 13855 3384 13864
rect 3332 13821 3341 13855
rect 3341 13821 3375 13855
rect 3375 13821 3384 13855
rect 3332 13812 3384 13821
rect 5448 13812 5500 13864
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 5448 13719 5500 13728
rect 5448 13685 5457 13719
rect 5457 13685 5491 13719
rect 5491 13685 5500 13719
rect 5448 13676 5500 13685
rect 8300 13880 8352 13932
rect 9404 13880 9456 13932
rect 11704 14025 11713 14059
rect 11713 14025 11747 14059
rect 11747 14025 11756 14059
rect 11704 14016 11756 14025
rect 11980 14059 12032 14068
rect 11980 14025 11989 14059
rect 11989 14025 12023 14059
rect 12023 14025 12032 14059
rect 11980 14016 12032 14025
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 12348 14016 12400 14068
rect 12256 13948 12308 14000
rect 18420 14059 18472 14068
rect 18420 14025 18429 14059
rect 18429 14025 18463 14059
rect 18463 14025 18472 14059
rect 18420 14016 18472 14025
rect 18512 13948 18564 14000
rect 19800 14016 19852 14068
rect 20536 14016 20588 14068
rect 22284 14016 22336 14068
rect 23756 14059 23808 14068
rect 23756 14025 23765 14059
rect 23765 14025 23799 14059
rect 23799 14025 23808 14059
rect 23756 14016 23808 14025
rect 5908 13812 5960 13864
rect 11796 13880 11848 13932
rect 11980 13880 12032 13932
rect 12808 13880 12860 13932
rect 8760 13744 8812 13796
rect 11980 13744 12032 13796
rect 18052 13880 18104 13932
rect 22100 13880 22152 13932
rect 22928 13880 22980 13932
rect 23112 13923 23164 13932
rect 23112 13889 23121 13923
rect 23121 13889 23155 13923
rect 23155 13889 23164 13923
rect 23112 13880 23164 13889
rect 25136 14016 25188 14068
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 24124 13991 24176 14000
rect 24124 13957 24133 13991
rect 24133 13957 24167 13991
rect 24167 13957 24176 13991
rect 24124 13948 24176 13957
rect 24768 13948 24820 14000
rect 25596 13880 25648 13932
rect 25780 14016 25832 14068
rect 26884 14016 26936 14068
rect 27436 14016 27488 14068
rect 32404 14016 32456 14068
rect 33048 14016 33100 14068
rect 29092 13991 29144 14000
rect 29092 13957 29101 13991
rect 29101 13957 29135 13991
rect 29135 13957 29144 13991
rect 29092 13948 29144 13957
rect 29276 13948 29328 14000
rect 32956 13948 33008 14000
rect 26700 13880 26752 13932
rect 27896 13880 27948 13932
rect 34796 14016 34848 14068
rect 35164 14016 35216 14068
rect 37280 14016 37332 14068
rect 38384 14016 38436 14068
rect 38568 14016 38620 14068
rect 39948 14016 40000 14068
rect 41144 14016 41196 14068
rect 36452 13991 36504 14000
rect 36452 13957 36461 13991
rect 36461 13957 36495 13991
rect 36495 13957 36504 13991
rect 36452 13948 36504 13957
rect 39764 13948 39816 14000
rect 41420 13948 41472 14000
rect 35348 13880 35400 13932
rect 38292 13880 38344 13932
rect 39120 13880 39172 13932
rect 39304 13880 39356 13932
rect 39488 13880 39540 13932
rect 17040 13812 17092 13864
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 18788 13855 18840 13864
rect 18788 13821 18797 13855
rect 18797 13821 18831 13855
rect 18831 13821 18840 13855
rect 18788 13812 18840 13821
rect 21640 13855 21692 13864
rect 21640 13821 21649 13855
rect 21649 13821 21683 13855
rect 21683 13821 21692 13855
rect 21640 13812 21692 13821
rect 22376 13812 22428 13864
rect 22836 13812 22888 13864
rect 25688 13812 25740 13864
rect 16488 13744 16540 13796
rect 25872 13812 25924 13864
rect 26056 13744 26108 13796
rect 28356 13855 28408 13864
rect 28356 13821 28365 13855
rect 28365 13821 28399 13855
rect 28399 13821 28408 13855
rect 28356 13812 28408 13821
rect 28448 13855 28500 13864
rect 28448 13821 28457 13855
rect 28457 13821 28491 13855
rect 28491 13821 28500 13855
rect 28448 13812 28500 13821
rect 30472 13855 30524 13864
rect 30472 13821 30481 13855
rect 30481 13821 30515 13855
rect 30515 13821 30524 13855
rect 30472 13812 30524 13821
rect 32128 13812 32180 13864
rect 33968 13855 34020 13864
rect 33968 13821 33977 13855
rect 33977 13821 34011 13855
rect 34011 13821 34020 13855
rect 33968 13812 34020 13821
rect 5816 13676 5868 13728
rect 11336 13719 11388 13728
rect 11336 13685 11345 13719
rect 11345 13685 11379 13719
rect 11379 13685 11388 13719
rect 11336 13676 11388 13685
rect 12532 13719 12584 13728
rect 12532 13685 12541 13719
rect 12541 13685 12575 13719
rect 12575 13685 12584 13719
rect 12532 13676 12584 13685
rect 15292 13676 15344 13728
rect 16396 13676 16448 13728
rect 17960 13676 18012 13728
rect 23480 13676 23532 13728
rect 28264 13744 28316 13796
rect 32312 13744 32364 13796
rect 32956 13744 33008 13796
rect 34336 13787 34388 13796
rect 34336 13753 34345 13787
rect 34345 13753 34379 13787
rect 34379 13753 34388 13787
rect 34336 13744 34388 13753
rect 34612 13855 34664 13864
rect 34612 13821 34621 13855
rect 34621 13821 34655 13855
rect 34655 13821 34664 13855
rect 34612 13812 34664 13821
rect 35440 13744 35492 13796
rect 39212 13812 39264 13864
rect 39764 13812 39816 13864
rect 37464 13744 37516 13796
rect 37648 13744 37700 13796
rect 38200 13744 38252 13796
rect 40776 13744 40828 13796
rect 42156 13855 42208 13864
rect 42156 13821 42165 13855
rect 42165 13821 42199 13855
rect 42199 13821 42208 13855
rect 42156 13812 42208 13821
rect 26976 13719 27028 13728
rect 26976 13685 26985 13719
rect 26985 13685 27019 13719
rect 27019 13685 27028 13719
rect 26976 13676 27028 13685
rect 27712 13719 27764 13728
rect 27712 13685 27721 13719
rect 27721 13685 27755 13719
rect 27755 13685 27764 13719
rect 27712 13676 27764 13685
rect 39396 13676 39448 13728
rect 40684 13676 40736 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2964 13472 3016 13524
rect 3332 13472 3384 13524
rect 6552 13515 6604 13524
rect 6552 13481 6561 13515
rect 6561 13481 6595 13515
rect 6595 13481 6604 13515
rect 6552 13472 6604 13481
rect 1584 13336 1636 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 5356 13404 5408 13456
rect 10692 13472 10744 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 11612 13404 11664 13456
rect 5540 13336 5592 13388
rect 5724 13336 5776 13388
rect 2780 13200 2832 13252
rect 4712 13132 4764 13184
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 21916 13472 21968 13524
rect 18788 13404 18840 13456
rect 21640 13404 21692 13456
rect 23572 13404 23624 13456
rect 25228 13447 25280 13456
rect 25228 13413 25237 13447
rect 25237 13413 25271 13447
rect 25271 13413 25280 13447
rect 25228 13404 25280 13413
rect 26884 13404 26936 13456
rect 28448 13404 28500 13456
rect 28540 13404 28592 13456
rect 29000 13404 29052 13456
rect 29920 13404 29972 13456
rect 6736 13268 6788 13320
rect 8760 13268 8812 13320
rect 16396 13336 16448 13388
rect 18420 13336 18472 13388
rect 18512 13336 18564 13388
rect 21088 13336 21140 13388
rect 22376 13336 22428 13388
rect 24860 13336 24912 13388
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 11336 13268 11388 13320
rect 11520 13268 11572 13320
rect 14556 13268 14608 13320
rect 5448 13200 5500 13252
rect 5356 13132 5408 13184
rect 6000 13175 6052 13184
rect 6000 13141 6009 13175
rect 6009 13141 6043 13175
rect 6043 13141 6052 13175
rect 6000 13132 6052 13141
rect 6460 13175 6512 13184
rect 6460 13141 6469 13175
rect 6469 13141 6503 13175
rect 6503 13141 6512 13175
rect 6460 13132 6512 13141
rect 8024 13243 8076 13252
rect 8024 13209 8033 13243
rect 8033 13209 8067 13243
rect 8067 13209 8076 13243
rect 8024 13200 8076 13209
rect 10324 13200 10376 13252
rect 12164 13243 12216 13252
rect 12164 13209 12173 13243
rect 12173 13209 12207 13243
rect 12207 13209 12216 13243
rect 12164 13200 12216 13209
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 19708 13268 19760 13320
rect 19892 13268 19944 13320
rect 24216 13268 24268 13320
rect 24676 13311 24728 13320
rect 24676 13277 24685 13311
rect 24685 13277 24719 13311
rect 24719 13277 24728 13311
rect 24676 13268 24728 13277
rect 25596 13379 25648 13388
rect 25596 13345 25605 13379
rect 25605 13345 25639 13379
rect 25639 13345 25648 13379
rect 25596 13336 25648 13345
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 11428 13132 11480 13184
rect 12992 13132 13044 13184
rect 13452 13132 13504 13184
rect 14924 13200 14976 13252
rect 13728 13132 13780 13184
rect 19524 13243 19576 13252
rect 19524 13209 19533 13243
rect 19533 13209 19567 13243
rect 19567 13209 19576 13243
rect 19524 13200 19576 13209
rect 19984 13200 20036 13252
rect 17868 13132 17920 13184
rect 22468 13200 22520 13252
rect 22836 13200 22888 13252
rect 25136 13268 25188 13320
rect 27528 13311 27580 13320
rect 27528 13277 27537 13311
rect 27537 13277 27571 13311
rect 27571 13277 27580 13311
rect 27528 13268 27580 13277
rect 27712 13311 27764 13320
rect 27712 13277 27721 13311
rect 27721 13277 27755 13311
rect 27755 13277 27764 13311
rect 27712 13268 27764 13277
rect 30564 13336 30616 13388
rect 23756 13132 23808 13184
rect 25872 13200 25924 13252
rect 26056 13200 26108 13252
rect 27252 13200 27304 13252
rect 26976 13132 27028 13184
rect 27620 13132 27672 13184
rect 28540 13243 28592 13252
rect 28540 13209 28549 13243
rect 28549 13209 28583 13243
rect 28583 13209 28592 13243
rect 28540 13200 28592 13209
rect 28724 13311 28776 13320
rect 28724 13277 28733 13311
rect 28733 13277 28767 13311
rect 28767 13277 28776 13311
rect 28724 13268 28776 13277
rect 32404 13472 32456 13524
rect 37372 13472 37424 13524
rect 38108 13472 38160 13524
rect 33968 13404 34020 13456
rect 33048 13379 33100 13388
rect 33048 13345 33057 13379
rect 33057 13345 33091 13379
rect 33091 13345 33100 13379
rect 33048 13336 33100 13345
rect 34888 13311 34940 13320
rect 34888 13277 34897 13311
rect 34897 13277 34931 13311
rect 34931 13277 34940 13311
rect 34888 13268 34940 13277
rect 35440 13336 35492 13388
rect 36820 13404 36872 13456
rect 39028 13472 39080 13524
rect 39396 13515 39448 13524
rect 39396 13481 39405 13515
rect 39405 13481 39439 13515
rect 39439 13481 39448 13515
rect 39396 13472 39448 13481
rect 42156 13515 42208 13524
rect 42156 13481 42165 13515
rect 42165 13481 42199 13515
rect 42199 13481 42208 13515
rect 42156 13472 42208 13481
rect 35072 13311 35124 13320
rect 35072 13277 35081 13311
rect 35081 13277 35115 13311
rect 35115 13277 35124 13311
rect 35072 13268 35124 13277
rect 30104 13200 30156 13252
rect 30656 13200 30708 13252
rect 37464 13311 37516 13320
rect 37464 13277 37473 13311
rect 37473 13277 37507 13311
rect 37507 13277 37516 13311
rect 37464 13268 37516 13277
rect 28264 13175 28316 13184
rect 28264 13141 28273 13175
rect 28273 13141 28307 13175
rect 28307 13141 28316 13175
rect 28264 13132 28316 13141
rect 28908 13175 28960 13184
rect 28908 13141 28917 13175
rect 28917 13141 28951 13175
rect 28951 13141 28960 13175
rect 28908 13132 28960 13141
rect 32128 13132 32180 13184
rect 35072 13132 35124 13184
rect 36084 13200 36136 13252
rect 36268 13200 36320 13252
rect 38476 13200 38528 13252
rect 40684 13379 40736 13388
rect 40684 13345 40693 13379
rect 40693 13345 40727 13379
rect 40727 13345 40736 13379
rect 40684 13336 40736 13345
rect 39120 13311 39172 13320
rect 39120 13277 39129 13311
rect 39129 13277 39163 13311
rect 39163 13277 39172 13311
rect 39120 13268 39172 13277
rect 39212 13311 39264 13320
rect 39212 13277 39221 13311
rect 39221 13277 39255 13311
rect 39255 13277 39264 13311
rect 39212 13268 39264 13277
rect 37280 13132 37332 13184
rect 39120 13132 39172 13184
rect 39488 13268 39540 13320
rect 41144 13200 41196 13252
rect 40224 13132 40276 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 6000 12928 6052 12980
rect 8024 12928 8076 12980
rect 9588 12928 9640 12980
rect 10416 12928 10468 12980
rect 16580 12928 16632 12980
rect 18144 12928 18196 12980
rect 18420 12928 18472 12980
rect 3240 12860 3292 12912
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 4620 12792 4672 12844
rect 5448 12792 5500 12844
rect 12532 12860 12584 12912
rect 13360 12860 13412 12912
rect 13452 12903 13504 12912
rect 13452 12869 13461 12903
rect 13461 12869 13495 12903
rect 13495 12869 13504 12903
rect 13452 12860 13504 12869
rect 14556 12860 14608 12912
rect 14924 12860 14976 12912
rect 15108 12860 15160 12912
rect 6828 12792 6880 12844
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 9956 12792 10008 12844
rect 10692 12792 10744 12844
rect 11244 12792 11296 12844
rect 11888 12792 11940 12844
rect 1400 12724 1452 12776
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 3976 12724 4028 12776
rect 5632 12724 5684 12776
rect 6552 12724 6604 12776
rect 12072 12767 12124 12776
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 13728 12792 13780 12844
rect 16488 12792 16540 12844
rect 19892 12928 19944 12980
rect 22468 12971 22520 12980
rect 22468 12937 22477 12971
rect 22477 12937 22511 12971
rect 22511 12937 22520 12971
rect 22468 12928 22520 12937
rect 22928 12971 22980 12980
rect 22928 12937 22937 12971
rect 22937 12937 22971 12971
rect 22971 12937 22980 12971
rect 22928 12928 22980 12937
rect 20168 12860 20220 12912
rect 28724 12928 28776 12980
rect 29092 12928 29144 12980
rect 29460 12971 29512 12980
rect 29460 12937 29469 12971
rect 29469 12937 29503 12971
rect 29503 12937 29512 12971
rect 29460 12928 29512 12937
rect 30472 12928 30524 12980
rect 32220 12928 32272 12980
rect 33416 12971 33468 12980
rect 33416 12937 33425 12971
rect 33425 12937 33459 12971
rect 33459 12937 33468 12971
rect 33416 12928 33468 12937
rect 35348 12928 35400 12980
rect 35532 12928 35584 12980
rect 36084 12928 36136 12980
rect 36820 12928 36872 12980
rect 25136 12860 25188 12912
rect 26148 12860 26200 12912
rect 2872 12656 2924 12708
rect 3424 12656 3476 12708
rect 6828 12656 6880 12708
rect 8576 12656 8628 12708
rect 9864 12656 9916 12708
rect 11428 12656 11480 12708
rect 12164 12656 12216 12708
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 19432 12792 19484 12844
rect 20076 12792 20128 12844
rect 23572 12792 23624 12844
rect 25320 12792 25372 12844
rect 27344 12792 27396 12844
rect 19340 12724 19392 12776
rect 13636 12656 13688 12708
rect 17868 12656 17920 12708
rect 19616 12656 19668 12708
rect 23480 12724 23532 12776
rect 23664 12724 23716 12776
rect 27620 12835 27672 12844
rect 27620 12801 27629 12835
rect 27629 12801 27663 12835
rect 27663 12801 27672 12835
rect 27620 12792 27672 12801
rect 28908 12860 28960 12912
rect 28080 12792 28132 12844
rect 28172 12835 28224 12844
rect 28172 12801 28181 12835
rect 28181 12801 28215 12835
rect 28215 12801 28224 12835
rect 28172 12792 28224 12801
rect 28724 12792 28776 12844
rect 29368 12860 29420 12912
rect 29644 12860 29696 12912
rect 30380 12860 30432 12912
rect 34428 12860 34480 12912
rect 38568 12928 38620 12980
rect 39396 12928 39448 12980
rect 2780 12588 2832 12640
rect 3056 12588 3108 12640
rect 3700 12588 3752 12640
rect 4712 12588 4764 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 6460 12588 6512 12640
rect 9680 12588 9732 12640
rect 11152 12588 11204 12640
rect 11980 12588 12032 12640
rect 13544 12631 13596 12640
rect 13544 12597 13553 12631
rect 13553 12597 13587 12631
rect 13587 12597 13596 12631
rect 13544 12588 13596 12597
rect 19340 12588 19392 12640
rect 24860 12588 24912 12640
rect 25136 12588 25188 12640
rect 27712 12656 27764 12708
rect 27988 12656 28040 12708
rect 28172 12656 28224 12708
rect 29276 12835 29328 12844
rect 29276 12801 29285 12835
rect 29285 12801 29319 12835
rect 29319 12801 29328 12835
rect 29276 12792 29328 12801
rect 40500 12860 40552 12912
rect 35716 12835 35768 12844
rect 35716 12801 35725 12835
rect 35725 12801 35759 12835
rect 35759 12801 35768 12835
rect 35716 12792 35768 12801
rect 37556 12792 37608 12844
rect 31116 12767 31168 12776
rect 31116 12733 31125 12767
rect 31125 12733 31159 12767
rect 31159 12733 31168 12767
rect 31116 12724 31168 12733
rect 31576 12724 31628 12776
rect 31852 12724 31904 12776
rect 33140 12724 33192 12776
rect 33508 12767 33560 12776
rect 33508 12733 33517 12767
rect 33517 12733 33551 12767
rect 33551 12733 33560 12767
rect 33508 12724 33560 12733
rect 33600 12724 33652 12776
rect 34520 12724 34572 12776
rect 36544 12724 36596 12776
rect 38844 12724 38896 12776
rect 27620 12588 27672 12640
rect 28632 12631 28684 12640
rect 28632 12597 28641 12631
rect 28641 12597 28675 12631
rect 28675 12597 28684 12631
rect 28632 12588 28684 12597
rect 28724 12588 28776 12640
rect 31484 12588 31536 12640
rect 32312 12588 32364 12640
rect 34612 12588 34664 12640
rect 35900 12631 35952 12640
rect 35900 12597 35909 12631
rect 35909 12597 35943 12631
rect 35943 12597 35952 12631
rect 37648 12656 37700 12708
rect 35900 12588 35952 12597
rect 37464 12588 37516 12640
rect 38476 12588 38528 12640
rect 39212 12767 39264 12776
rect 39212 12733 39221 12767
rect 39221 12733 39255 12767
rect 39255 12733 39264 12767
rect 39212 12724 39264 12733
rect 40408 12792 40460 12844
rect 41512 12792 41564 12844
rect 42156 12792 42208 12844
rect 40684 12767 40736 12776
rect 40684 12733 40693 12767
rect 40693 12733 40727 12767
rect 40727 12733 40736 12767
rect 40684 12724 40736 12733
rect 39212 12588 39264 12640
rect 39304 12588 39356 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1768 12384 1820 12436
rect 5632 12384 5684 12436
rect 5724 12427 5776 12436
rect 5724 12393 5733 12427
rect 5733 12393 5767 12427
rect 5767 12393 5776 12427
rect 5724 12384 5776 12393
rect 2688 12316 2740 12368
rect 5448 12248 5500 12300
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 5724 12248 5776 12300
rect 6736 12291 6788 12300
rect 6736 12257 6745 12291
rect 6745 12257 6779 12291
rect 6779 12257 6788 12291
rect 6736 12248 6788 12257
rect 2872 12180 2924 12232
rect 3424 12180 3476 12232
rect 2780 12112 2832 12164
rect 3608 12180 3660 12232
rect 4068 12180 4120 12232
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 4620 12180 4672 12232
rect 5172 12180 5224 12232
rect 4528 12112 4580 12164
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 7012 12180 7064 12232
rect 6644 12155 6696 12164
rect 6644 12121 6653 12155
rect 6653 12121 6687 12155
rect 6687 12121 6696 12155
rect 6644 12112 6696 12121
rect 7472 12180 7524 12232
rect 12072 12384 12124 12436
rect 13452 12384 13504 12436
rect 15016 12384 15068 12436
rect 9404 12291 9456 12300
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 9404 12248 9456 12257
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 11336 12248 11388 12300
rect 10784 12180 10836 12232
rect 11152 12180 11204 12232
rect 12164 12316 12216 12368
rect 12440 12316 12492 12368
rect 3332 12087 3384 12096
rect 3332 12053 3341 12087
rect 3341 12053 3375 12087
rect 3375 12053 3384 12087
rect 3332 12044 3384 12053
rect 4804 12044 4856 12096
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 6736 12044 6788 12096
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 8852 12044 8904 12096
rect 8944 12044 8996 12096
rect 12440 12180 12492 12232
rect 13360 12248 13412 12300
rect 13544 12223 13596 12232
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 13636 12180 13688 12232
rect 12808 12155 12860 12164
rect 12808 12121 12817 12155
rect 12817 12121 12851 12155
rect 12851 12121 12860 12155
rect 12808 12112 12860 12121
rect 15844 12180 15896 12232
rect 12900 12044 12952 12096
rect 14556 12044 14608 12096
rect 16580 12112 16632 12164
rect 17592 12223 17644 12232
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 20168 12359 20220 12368
rect 20168 12325 20177 12359
rect 20177 12325 20211 12359
rect 20211 12325 20220 12359
rect 20168 12316 20220 12325
rect 22192 12427 22244 12436
rect 22192 12393 22201 12427
rect 22201 12393 22235 12427
rect 22235 12393 22244 12427
rect 22192 12384 22244 12393
rect 23204 12384 23256 12436
rect 24308 12384 24360 12436
rect 23664 12316 23716 12368
rect 21456 12248 21508 12300
rect 17868 12223 17920 12232
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 19156 12180 19208 12232
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20260 12180 20312 12189
rect 22376 12180 22428 12232
rect 22652 12291 22704 12300
rect 22652 12257 22661 12291
rect 22661 12257 22695 12291
rect 22695 12257 22704 12291
rect 22652 12248 22704 12257
rect 22928 12248 22980 12300
rect 19800 12112 19852 12164
rect 20168 12112 20220 12164
rect 22192 12112 22244 12164
rect 22284 12112 22336 12164
rect 22744 12112 22796 12164
rect 24952 12291 25004 12300
rect 24952 12257 24961 12291
rect 24961 12257 24995 12291
rect 24995 12257 25004 12291
rect 24952 12248 25004 12257
rect 25228 12384 25280 12436
rect 26424 12384 26476 12436
rect 26976 12384 27028 12436
rect 29552 12384 29604 12436
rect 31116 12384 31168 12436
rect 32956 12427 33008 12436
rect 32956 12393 32965 12427
rect 32965 12393 32999 12427
rect 32999 12393 33008 12427
rect 32956 12384 33008 12393
rect 34704 12384 34756 12436
rect 38384 12384 38436 12436
rect 39396 12384 39448 12436
rect 39488 12384 39540 12436
rect 25872 12248 25924 12300
rect 24124 12180 24176 12232
rect 24768 12180 24820 12232
rect 25780 12180 25832 12232
rect 26056 12223 26108 12232
rect 26056 12189 26065 12223
rect 26065 12189 26099 12223
rect 26099 12189 26108 12223
rect 26056 12180 26108 12189
rect 26148 12180 26200 12232
rect 27988 12248 28040 12300
rect 26516 12112 26568 12164
rect 16120 12044 16172 12096
rect 19524 12044 19576 12096
rect 20076 12044 20128 12096
rect 22468 12044 22520 12096
rect 24492 12087 24544 12096
rect 24492 12053 24501 12087
rect 24501 12053 24535 12087
rect 24535 12053 24544 12087
rect 24492 12044 24544 12053
rect 28908 12112 28960 12164
rect 29460 12248 29512 12300
rect 31668 12248 31720 12300
rect 33324 12248 33376 12300
rect 33692 12291 33744 12300
rect 33692 12257 33701 12291
rect 33701 12257 33735 12291
rect 33735 12257 33744 12291
rect 33692 12248 33744 12257
rect 33876 12291 33928 12300
rect 33876 12257 33885 12291
rect 33885 12257 33919 12291
rect 33919 12257 33928 12291
rect 33876 12248 33928 12257
rect 33968 12248 34020 12300
rect 29184 12223 29236 12232
rect 29184 12189 29193 12223
rect 29193 12189 29227 12223
rect 29227 12189 29236 12223
rect 29184 12180 29236 12189
rect 29276 12180 29328 12232
rect 30196 12180 30248 12232
rect 32588 12223 32640 12232
rect 32588 12189 32597 12223
rect 32597 12189 32631 12223
rect 32631 12189 32640 12223
rect 32588 12180 32640 12189
rect 32956 12223 33008 12232
rect 32956 12189 32965 12223
rect 32965 12189 32999 12223
rect 32999 12189 33008 12223
rect 32956 12180 33008 12189
rect 34612 12248 34664 12300
rect 35992 12316 36044 12368
rect 35900 12248 35952 12300
rect 36912 12248 36964 12300
rect 37464 12248 37516 12300
rect 38844 12248 38896 12300
rect 39028 12248 39080 12300
rect 36360 12223 36412 12232
rect 36360 12189 36369 12223
rect 36369 12189 36403 12223
rect 36403 12189 36412 12223
rect 36360 12180 36412 12189
rect 37188 12223 37240 12232
rect 37188 12189 37197 12223
rect 37197 12189 37231 12223
rect 37231 12189 37240 12223
rect 37188 12180 37240 12189
rect 37556 12180 37608 12232
rect 31024 12112 31076 12164
rect 28632 12044 28684 12096
rect 30380 12044 30432 12096
rect 30840 12087 30892 12096
rect 30840 12053 30849 12087
rect 30849 12053 30883 12087
rect 30883 12053 30892 12087
rect 30840 12044 30892 12053
rect 32312 12155 32364 12164
rect 32312 12121 32321 12155
rect 32321 12121 32355 12155
rect 32355 12121 32364 12155
rect 32312 12112 32364 12121
rect 32680 12155 32732 12164
rect 32680 12121 32689 12155
rect 32689 12121 32723 12155
rect 32723 12121 32732 12155
rect 32680 12112 32732 12121
rect 32864 12044 32916 12096
rect 33048 12044 33100 12096
rect 35348 12112 35400 12164
rect 35532 12112 35584 12164
rect 37372 12155 37424 12164
rect 37372 12121 37381 12155
rect 37381 12121 37415 12155
rect 37415 12121 37424 12155
rect 37372 12112 37424 12121
rect 38200 12112 38252 12164
rect 39212 12180 39264 12232
rect 39580 12316 39632 12368
rect 39948 12248 40000 12300
rect 39580 12180 39632 12232
rect 40224 12223 40276 12232
rect 40224 12189 40233 12223
rect 40233 12189 40267 12223
rect 40267 12189 40276 12223
rect 40224 12180 40276 12189
rect 40500 12291 40552 12300
rect 40500 12257 40509 12291
rect 40509 12257 40543 12291
rect 40543 12257 40552 12291
rect 40500 12248 40552 12257
rect 40684 12248 40736 12300
rect 41512 12223 41564 12232
rect 41512 12189 41521 12223
rect 41521 12189 41555 12223
rect 41555 12189 41564 12223
rect 41512 12180 41564 12189
rect 38936 12112 38988 12164
rect 39304 12155 39356 12164
rect 39304 12121 39313 12155
rect 39313 12121 39347 12155
rect 39347 12121 39356 12155
rect 39304 12112 39356 12121
rect 39764 12112 39816 12164
rect 33232 12087 33284 12096
rect 33232 12053 33241 12087
rect 33241 12053 33275 12087
rect 33275 12053 33284 12087
rect 33232 12044 33284 12053
rect 33324 12044 33376 12096
rect 34152 12044 34204 12096
rect 34796 12044 34848 12096
rect 36728 12044 36780 12096
rect 37924 12044 37976 12096
rect 39212 12044 39264 12096
rect 40592 12087 40644 12096
rect 40592 12053 40601 12087
rect 40601 12053 40635 12087
rect 40635 12053 40644 12087
rect 40592 12044 40644 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 3976 11840 4028 11892
rect 4712 11840 4764 11892
rect 5356 11840 5408 11892
rect 5908 11840 5960 11892
rect 6552 11840 6604 11892
rect 7472 11883 7524 11892
rect 7472 11849 7481 11883
rect 7481 11849 7515 11883
rect 7515 11849 7524 11883
rect 7472 11840 7524 11849
rect 4160 11815 4212 11824
rect 4160 11781 4169 11815
rect 4169 11781 4203 11815
rect 4203 11781 4212 11815
rect 4160 11772 4212 11781
rect 5448 11772 5500 11824
rect 5816 11772 5868 11824
rect 6736 11772 6788 11824
rect 7380 11815 7432 11824
rect 7380 11781 7389 11815
rect 7389 11781 7423 11815
rect 7423 11781 7432 11815
rect 7380 11772 7432 11781
rect 3240 11704 3292 11756
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 4804 11704 4856 11756
rect 5264 11704 5316 11756
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 1492 11679 1544 11688
rect 1492 11645 1501 11679
rect 1501 11645 1535 11679
rect 1535 11645 1544 11679
rect 1492 11636 1544 11645
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 4528 11636 4580 11688
rect 6552 11704 6604 11756
rect 6828 11704 6880 11756
rect 8300 11840 8352 11892
rect 8392 11840 8444 11892
rect 8576 11815 8628 11824
rect 8576 11781 8585 11815
rect 8585 11781 8619 11815
rect 8619 11781 8628 11815
rect 8576 11772 8628 11781
rect 9496 11772 9548 11824
rect 10048 11840 10100 11892
rect 12072 11840 12124 11892
rect 12440 11840 12492 11892
rect 12808 11883 12860 11892
rect 12808 11849 12817 11883
rect 12817 11849 12851 11883
rect 12851 11849 12860 11883
rect 12808 11840 12860 11849
rect 7012 11636 7064 11688
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 8852 11704 8904 11756
rect 3424 11568 3476 11620
rect 9496 11636 9548 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 10692 11636 10744 11688
rect 11888 11636 11940 11688
rect 12164 11704 12216 11756
rect 12532 11772 12584 11824
rect 13360 11840 13412 11892
rect 15108 11840 15160 11892
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 13176 11772 13228 11824
rect 14004 11772 14056 11824
rect 19156 11883 19208 11892
rect 19156 11849 19165 11883
rect 19165 11849 19199 11883
rect 19199 11849 19208 11883
rect 19156 11840 19208 11849
rect 19984 11840 20036 11892
rect 22376 11840 22428 11892
rect 20720 11772 20772 11824
rect 13452 11704 13504 11756
rect 4068 11500 4120 11552
rect 5632 11500 5684 11552
rect 7472 11500 7524 11552
rect 8944 11543 8996 11552
rect 8944 11509 8953 11543
rect 8953 11509 8987 11543
rect 8987 11509 8996 11543
rect 8944 11500 8996 11509
rect 9036 11500 9088 11552
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 12256 11568 12308 11620
rect 10140 11500 10192 11509
rect 11888 11500 11940 11552
rect 13176 11636 13228 11688
rect 13360 11636 13412 11688
rect 12808 11568 12860 11620
rect 14556 11747 14608 11756
rect 14556 11713 14565 11747
rect 14565 11713 14599 11747
rect 14599 11713 14608 11747
rect 14556 11704 14608 11713
rect 15844 11704 15896 11756
rect 16580 11704 16632 11756
rect 22928 11772 22980 11824
rect 24124 11772 24176 11824
rect 13912 11636 13964 11688
rect 14464 11679 14516 11688
rect 14464 11645 14473 11679
rect 14473 11645 14507 11679
rect 14507 11645 14516 11679
rect 14464 11636 14516 11645
rect 16488 11636 16540 11688
rect 19432 11636 19484 11688
rect 19616 11636 19668 11688
rect 21364 11747 21416 11756
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 22376 11747 22428 11756
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 26148 11840 26200 11892
rect 27528 11840 27580 11892
rect 27620 11840 27672 11892
rect 24492 11815 24544 11824
rect 24492 11781 24501 11815
rect 24501 11781 24535 11815
rect 24535 11781 24544 11815
rect 24492 11772 24544 11781
rect 25780 11772 25832 11824
rect 26332 11772 26384 11824
rect 26976 11704 27028 11756
rect 27068 11704 27120 11756
rect 27804 11772 27856 11824
rect 29000 11840 29052 11892
rect 30932 11840 30984 11892
rect 32588 11840 32640 11892
rect 28908 11772 28960 11824
rect 30564 11772 30616 11824
rect 31852 11815 31904 11824
rect 31852 11781 31861 11815
rect 31861 11781 31895 11815
rect 31895 11781 31904 11815
rect 31852 11772 31904 11781
rect 20536 11636 20588 11688
rect 22284 11636 22336 11688
rect 22652 11679 22704 11688
rect 22652 11645 22661 11679
rect 22661 11645 22695 11679
rect 22695 11645 22704 11679
rect 22652 11636 22704 11645
rect 20076 11568 20128 11620
rect 13176 11500 13228 11552
rect 13728 11500 13780 11552
rect 15476 11500 15528 11552
rect 19984 11500 20036 11552
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 24860 11500 24912 11552
rect 25228 11500 25280 11552
rect 25504 11500 25556 11552
rect 26056 11500 26108 11552
rect 26608 11636 26660 11688
rect 27252 11679 27304 11688
rect 27252 11645 27261 11679
rect 27261 11645 27295 11679
rect 27295 11645 27304 11679
rect 27252 11636 27304 11645
rect 27896 11747 27948 11756
rect 27896 11713 27905 11747
rect 27905 11713 27939 11747
rect 27939 11713 27948 11747
rect 27896 11704 27948 11713
rect 31024 11704 31076 11756
rect 33232 11772 33284 11824
rect 33416 11772 33468 11824
rect 36176 11840 36228 11892
rect 36360 11840 36412 11892
rect 36728 11883 36780 11892
rect 36728 11849 36737 11883
rect 36737 11849 36771 11883
rect 36771 11849 36780 11883
rect 36728 11840 36780 11849
rect 36820 11883 36872 11892
rect 36820 11849 36829 11883
rect 36829 11849 36863 11883
rect 36863 11849 36872 11883
rect 36820 11840 36872 11849
rect 34796 11815 34848 11824
rect 34796 11781 34805 11815
rect 34805 11781 34839 11815
rect 34839 11781 34848 11815
rect 34796 11772 34848 11781
rect 35348 11772 35400 11824
rect 40592 11840 40644 11892
rect 40684 11883 40736 11892
rect 40684 11849 40693 11883
rect 40693 11849 40727 11883
rect 40727 11849 40736 11883
rect 40684 11840 40736 11849
rect 30564 11636 30616 11688
rect 31392 11636 31444 11688
rect 31576 11679 31628 11688
rect 31576 11645 31585 11679
rect 31585 11645 31619 11679
rect 31619 11645 31628 11679
rect 31576 11636 31628 11645
rect 29184 11568 29236 11620
rect 32036 11568 32088 11620
rect 32496 11568 32548 11620
rect 34520 11568 34572 11620
rect 36084 11568 36136 11620
rect 37648 11636 37700 11688
rect 37924 11636 37976 11688
rect 38476 11636 38528 11688
rect 41144 11704 41196 11756
rect 37556 11568 37608 11620
rect 38384 11568 38436 11620
rect 38568 11568 38620 11620
rect 28724 11500 28776 11552
rect 29828 11500 29880 11552
rect 30196 11500 30248 11552
rect 35532 11500 35584 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 4068 11296 4120 11348
rect 8944 11296 8996 11348
rect 9312 11296 9364 11348
rect 12532 11339 12584 11348
rect 12532 11305 12541 11339
rect 12541 11305 12575 11339
rect 12575 11305 12584 11339
rect 12532 11296 12584 11305
rect 13084 11296 13136 11348
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 14464 11296 14516 11348
rect 17592 11296 17644 11348
rect 3240 11228 3292 11280
rect 1492 11160 1544 11212
rect 2872 11160 2924 11212
rect 3516 11160 3568 11212
rect 7380 11228 7432 11280
rect 10692 11271 10744 11280
rect 10692 11237 10701 11271
rect 10701 11237 10735 11271
rect 10735 11237 10744 11271
rect 10692 11228 10744 11237
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 8852 11160 8904 11212
rect 11520 11160 11572 11212
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 3240 11024 3292 11076
rect 2780 10956 2832 11008
rect 4252 10956 4304 11008
rect 4896 10956 4948 11008
rect 5448 10956 5500 11008
rect 5908 10956 5960 11008
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 8668 11135 8720 11144
rect 8668 11101 8677 11135
rect 8677 11101 8711 11135
rect 8711 11101 8720 11135
rect 8668 11092 8720 11101
rect 10324 11092 10376 11144
rect 11704 11092 11756 11144
rect 12532 11092 12584 11144
rect 12992 11160 13044 11212
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 14004 11160 14056 11212
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 16488 11160 16540 11212
rect 18972 11228 19024 11280
rect 19616 11296 19668 11348
rect 22652 11296 22704 11348
rect 22468 11228 22520 11280
rect 29184 11296 29236 11348
rect 30380 11296 30432 11348
rect 19524 11203 19576 11212
rect 19524 11169 19533 11203
rect 19533 11169 19567 11203
rect 19567 11169 19576 11203
rect 19524 11160 19576 11169
rect 19892 11160 19944 11212
rect 20536 11160 20588 11212
rect 24860 11228 24912 11280
rect 26516 11228 26568 11280
rect 29276 11228 29328 11280
rect 31392 11296 31444 11348
rect 32772 11296 32824 11348
rect 34152 11296 34204 11348
rect 34612 11296 34664 11348
rect 35532 11339 35584 11348
rect 35532 11305 35541 11339
rect 35541 11305 35575 11339
rect 35575 11305 35584 11339
rect 35532 11296 35584 11305
rect 37188 11296 37240 11348
rect 31576 11228 31628 11280
rect 33048 11228 33100 11280
rect 35348 11228 35400 11280
rect 35440 11228 35492 11280
rect 9312 11024 9364 11076
rect 9036 10956 9088 11008
rect 11888 10999 11940 11008
rect 11888 10965 11897 10999
rect 11897 10965 11931 10999
rect 11931 10965 11940 10999
rect 11888 10956 11940 10965
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 12072 10956 12124 10965
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 18328 11092 18380 11144
rect 23204 11203 23256 11212
rect 23204 11169 23213 11203
rect 23213 11169 23247 11203
rect 23247 11169 23256 11203
rect 23204 11160 23256 11169
rect 24124 11203 24176 11212
rect 24124 11169 24133 11203
rect 24133 11169 24167 11203
rect 24167 11169 24176 11203
rect 24124 11160 24176 11169
rect 26424 11160 26476 11212
rect 26608 11160 26660 11212
rect 31668 11160 31720 11212
rect 33508 11160 33560 11212
rect 35256 11160 35308 11212
rect 36084 11203 36136 11212
rect 36084 11169 36093 11203
rect 36093 11169 36127 11203
rect 36127 11169 36136 11203
rect 36084 11160 36136 11169
rect 12808 11024 12860 11076
rect 14556 11024 14608 11076
rect 15108 11024 15160 11076
rect 13176 10956 13228 11008
rect 13268 10999 13320 11008
rect 13268 10965 13293 10999
rect 13293 10965 13320 10999
rect 19432 11024 19484 11076
rect 20168 11024 20220 11076
rect 22376 11135 22428 11144
rect 22376 11101 22385 11135
rect 22385 11101 22419 11135
rect 22419 11101 22428 11135
rect 22376 11092 22428 11101
rect 23296 11092 23348 11144
rect 26332 11092 26384 11144
rect 27988 11092 28040 11144
rect 13268 10956 13320 10965
rect 18604 10956 18656 11008
rect 21088 10956 21140 11008
rect 22836 11024 22888 11076
rect 25228 11067 25280 11076
rect 25228 11033 25237 11067
rect 25237 11033 25271 11067
rect 25271 11033 25280 11067
rect 25228 11024 25280 11033
rect 29828 11067 29880 11076
rect 29828 11033 29837 11067
rect 29837 11033 29871 11067
rect 29871 11033 29880 11067
rect 29828 11024 29880 11033
rect 30472 11024 30524 11076
rect 23296 10956 23348 11008
rect 26792 10999 26844 11008
rect 26792 10965 26801 10999
rect 26801 10965 26835 10999
rect 26835 10965 26844 10999
rect 26792 10956 26844 10965
rect 27712 10999 27764 11008
rect 27712 10965 27721 10999
rect 27721 10965 27755 10999
rect 27755 10965 27764 10999
rect 27712 10956 27764 10965
rect 30564 10956 30616 11008
rect 31852 11092 31904 11144
rect 32496 11135 32548 11144
rect 32496 11101 32505 11135
rect 32505 11101 32539 11135
rect 32539 11101 32548 11135
rect 32496 11092 32548 11101
rect 32036 11024 32088 11076
rect 32772 11024 32824 11076
rect 34520 11092 34572 11144
rect 35348 11135 35400 11144
rect 35348 11101 35357 11135
rect 35357 11101 35391 11135
rect 35391 11101 35400 11135
rect 35348 11092 35400 11101
rect 35440 11135 35492 11144
rect 35440 11101 35449 11135
rect 35449 11101 35483 11135
rect 35483 11101 35492 11135
rect 35440 11092 35492 11101
rect 38384 11160 38436 11212
rect 33876 11024 33928 11076
rect 35164 11024 35216 11076
rect 37832 11135 37884 11144
rect 37832 11101 37841 11135
rect 37841 11101 37875 11135
rect 37875 11101 37884 11135
rect 37832 11092 37884 11101
rect 31944 10999 31996 11008
rect 31944 10965 31953 10999
rect 31953 10965 31987 10999
rect 31987 10965 31996 10999
rect 31944 10956 31996 10965
rect 32312 10956 32364 11008
rect 36360 10956 36412 11008
rect 37832 10956 37884 11008
rect 38292 10956 38344 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 1216 10752 1268 10804
rect 1768 10752 1820 10804
rect 3608 10752 3660 10804
rect 4804 10752 4856 10804
rect 3700 10684 3752 10736
rect 2688 10616 2740 10668
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 4528 10616 4580 10668
rect 4252 10480 4304 10532
rect 3148 10412 3200 10464
rect 4804 10548 4856 10600
rect 5632 10616 5684 10668
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 8392 10752 8444 10804
rect 8668 10752 8720 10804
rect 12808 10752 12860 10804
rect 5816 10616 5868 10625
rect 5448 10548 5500 10600
rect 6000 10591 6052 10600
rect 6000 10557 6009 10591
rect 6009 10557 6043 10591
rect 6043 10557 6052 10591
rect 6000 10548 6052 10557
rect 7104 10684 7156 10736
rect 5540 10523 5592 10532
rect 5540 10489 5549 10523
rect 5549 10489 5583 10523
rect 5583 10489 5592 10523
rect 5540 10480 5592 10489
rect 4620 10412 4672 10464
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 5264 10412 5316 10464
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 10324 10684 10376 10736
rect 13084 10684 13136 10736
rect 13728 10752 13780 10804
rect 14004 10795 14056 10804
rect 14004 10761 14013 10795
rect 14013 10761 14047 10795
rect 14047 10761 14056 10795
rect 14004 10752 14056 10761
rect 19432 10752 19484 10804
rect 22376 10752 22428 10804
rect 14464 10684 14516 10736
rect 15476 10727 15528 10736
rect 15476 10693 15485 10727
rect 15485 10693 15519 10727
rect 15519 10693 15528 10727
rect 15476 10684 15528 10693
rect 18604 10727 18656 10736
rect 18604 10693 18613 10727
rect 18613 10693 18647 10727
rect 18647 10693 18656 10727
rect 18604 10684 18656 10693
rect 7104 10548 7156 10600
rect 8208 10616 8260 10668
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 7932 10480 7984 10532
rect 8484 10480 8536 10532
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 9772 10548 9824 10600
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 12440 10548 12492 10600
rect 13268 10548 13320 10600
rect 13636 10548 13688 10600
rect 7288 10412 7340 10464
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 11428 10480 11480 10532
rect 12900 10480 12952 10532
rect 15752 10659 15804 10668
rect 15752 10625 15761 10659
rect 15761 10625 15795 10659
rect 15795 10625 15804 10659
rect 15752 10616 15804 10625
rect 20168 10616 20220 10668
rect 25228 10752 25280 10804
rect 25964 10795 26016 10804
rect 25964 10761 25973 10795
rect 25973 10761 26007 10795
rect 26007 10761 26016 10795
rect 25964 10752 26016 10761
rect 27712 10752 27764 10804
rect 28724 10795 28776 10804
rect 28724 10761 28733 10795
rect 28733 10761 28767 10795
rect 28767 10761 28776 10795
rect 28724 10752 28776 10761
rect 32496 10752 32548 10804
rect 32680 10752 32732 10804
rect 35256 10752 35308 10804
rect 36360 10752 36412 10804
rect 39120 10752 39172 10804
rect 39948 10752 40000 10804
rect 18328 10591 18380 10600
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 22192 10548 22244 10600
rect 23020 10591 23072 10600
rect 23020 10557 23029 10591
rect 23029 10557 23063 10591
rect 23063 10557 23072 10591
rect 23020 10548 23072 10557
rect 24216 10616 24268 10668
rect 26792 10684 26844 10736
rect 26884 10684 26936 10736
rect 27344 10616 27396 10668
rect 30840 10684 30892 10736
rect 33508 10684 33560 10736
rect 32312 10616 32364 10668
rect 34796 10616 34848 10668
rect 35532 10659 35584 10668
rect 35532 10625 35536 10659
rect 35536 10625 35570 10659
rect 35570 10625 35584 10659
rect 35532 10616 35584 10625
rect 38476 10684 38528 10736
rect 25136 10548 25188 10600
rect 25872 10548 25924 10600
rect 28908 10548 28960 10600
rect 29092 10548 29144 10600
rect 30196 10548 30248 10600
rect 32772 10591 32824 10600
rect 32772 10557 32781 10591
rect 32781 10557 32815 10591
rect 32815 10557 32824 10591
rect 32772 10548 32824 10557
rect 33140 10548 33192 10600
rect 34520 10591 34572 10600
rect 34520 10557 34529 10591
rect 34529 10557 34563 10591
rect 34563 10557 34572 10591
rect 34520 10548 34572 10557
rect 35348 10548 35400 10600
rect 36084 10659 36136 10668
rect 36084 10625 36093 10659
rect 36093 10625 36127 10659
rect 36127 10625 36136 10659
rect 36084 10616 36136 10625
rect 36360 10616 36412 10668
rect 36176 10548 36228 10600
rect 37372 10548 37424 10600
rect 37924 10659 37976 10668
rect 37924 10625 37933 10659
rect 37933 10625 37967 10659
rect 37967 10625 37976 10659
rect 37924 10616 37976 10625
rect 37832 10548 37884 10600
rect 38568 10548 38620 10600
rect 38936 10548 38988 10600
rect 40776 10659 40828 10668
rect 40776 10625 40785 10659
rect 40785 10625 40819 10659
rect 40819 10625 40828 10659
rect 40776 10616 40828 10625
rect 21272 10480 21324 10532
rect 26700 10480 26752 10532
rect 10048 10412 10100 10464
rect 13268 10455 13320 10464
rect 13268 10421 13277 10455
rect 13277 10421 13311 10455
rect 13311 10421 13320 10455
rect 13268 10412 13320 10421
rect 13912 10455 13964 10464
rect 13912 10421 13921 10455
rect 13921 10421 13955 10455
rect 13955 10421 13964 10455
rect 13912 10412 13964 10421
rect 20076 10455 20128 10464
rect 20076 10421 20085 10455
rect 20085 10421 20119 10455
rect 20119 10421 20128 10455
rect 20076 10412 20128 10421
rect 23756 10455 23808 10464
rect 23756 10421 23765 10455
rect 23765 10421 23799 10455
rect 23799 10421 23808 10455
rect 23756 10412 23808 10421
rect 26332 10412 26384 10464
rect 26516 10412 26568 10464
rect 30104 10412 30156 10464
rect 34336 10455 34388 10464
rect 34336 10421 34345 10455
rect 34345 10421 34379 10455
rect 34379 10421 34388 10455
rect 34336 10412 34388 10421
rect 35532 10480 35584 10532
rect 37648 10480 37700 10532
rect 37372 10412 37424 10464
rect 37464 10455 37516 10464
rect 37464 10421 37473 10455
rect 37473 10421 37507 10455
rect 37507 10421 37516 10455
rect 37464 10412 37516 10421
rect 38844 10412 38896 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2780 10208 2832 10260
rect 6000 10208 6052 10260
rect 7380 10208 7432 10260
rect 11796 10208 11848 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13728 10208 13780 10260
rect 22192 10251 22244 10260
rect 22192 10217 22201 10251
rect 22201 10217 22235 10251
rect 22235 10217 22244 10251
rect 22192 10208 22244 10217
rect 23296 10251 23348 10260
rect 23296 10217 23305 10251
rect 23305 10217 23339 10251
rect 23339 10217 23348 10251
rect 23296 10208 23348 10217
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 3424 10004 3476 10056
rect 4620 10004 4672 10056
rect 5448 10004 5500 10056
rect 6552 10140 6604 10192
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 5908 10004 5960 10056
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 11704 10072 11756 10124
rect 12072 10072 12124 10124
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 13912 10072 13964 10124
rect 21088 10072 21140 10124
rect 21364 10072 21416 10124
rect 5724 9979 5776 9988
rect 5724 9945 5733 9979
rect 5733 9945 5767 9979
rect 5767 9945 5776 9979
rect 5724 9936 5776 9945
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 6736 10004 6788 10056
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 18328 10004 18380 10056
rect 22284 10004 22336 10056
rect 22652 10047 22704 10056
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 22836 10047 22888 10056
rect 22836 10013 22845 10047
rect 22845 10013 22879 10047
rect 22879 10013 22888 10047
rect 22836 10004 22888 10013
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 23388 10004 23440 10056
rect 5356 9868 5408 9920
rect 14556 9936 14608 9988
rect 20168 9936 20220 9988
rect 21180 9936 21232 9988
rect 23664 10047 23716 10056
rect 23664 10013 23674 10047
rect 23674 10013 23708 10047
rect 23708 10013 23716 10047
rect 23664 10004 23716 10013
rect 27988 10183 28040 10192
rect 27988 10149 27997 10183
rect 27997 10149 28031 10183
rect 28031 10149 28040 10183
rect 27988 10140 28040 10149
rect 28264 10140 28316 10192
rect 24124 10072 24176 10124
rect 25044 10072 25096 10124
rect 26148 10072 26200 10124
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 6460 9911 6512 9920
rect 6460 9877 6469 9911
rect 6469 9877 6503 9911
rect 6503 9877 6512 9911
rect 6460 9868 6512 9877
rect 6644 9911 6696 9920
rect 6644 9877 6653 9911
rect 6653 9877 6687 9911
rect 6687 9877 6696 9911
rect 6644 9868 6696 9877
rect 8576 9868 8628 9920
rect 22836 9868 22888 9920
rect 25044 9936 25096 9988
rect 25504 10047 25556 10056
rect 25504 10013 25513 10047
rect 25513 10013 25547 10047
rect 25547 10013 25556 10047
rect 25504 10004 25556 10013
rect 28080 10049 28132 10056
rect 28080 10015 28089 10049
rect 28089 10015 28123 10049
rect 28123 10015 28132 10049
rect 28080 10004 28132 10015
rect 28264 10047 28316 10056
rect 28264 10013 28273 10047
rect 28273 10013 28307 10047
rect 28307 10013 28316 10047
rect 28264 10004 28316 10013
rect 28448 10208 28500 10260
rect 33140 10251 33192 10260
rect 33140 10217 33149 10251
rect 33149 10217 33183 10251
rect 33183 10217 33192 10251
rect 33140 10208 33192 10217
rect 34520 10208 34572 10260
rect 38568 10251 38620 10260
rect 38568 10217 38577 10251
rect 38577 10217 38611 10251
rect 38611 10217 38620 10251
rect 38568 10208 38620 10217
rect 30104 10115 30156 10124
rect 30104 10081 30113 10115
rect 30113 10081 30147 10115
rect 30147 10081 30156 10115
rect 30104 10072 30156 10081
rect 30196 10072 30248 10124
rect 26608 9936 26660 9988
rect 28172 9936 28224 9988
rect 27344 9868 27396 9920
rect 28540 10004 28592 10056
rect 30380 10004 30432 10056
rect 32680 10140 32732 10192
rect 31208 10115 31260 10124
rect 31208 10081 31217 10115
rect 31217 10081 31251 10115
rect 31251 10081 31260 10115
rect 31208 10072 31260 10081
rect 31760 10072 31812 10124
rect 32220 10072 32272 10124
rect 33140 10072 33192 10124
rect 34612 10072 34664 10124
rect 35348 10115 35400 10124
rect 35348 10081 35357 10115
rect 35357 10081 35391 10115
rect 35391 10081 35400 10115
rect 35348 10072 35400 10081
rect 35440 10072 35492 10124
rect 29092 9979 29144 9988
rect 29092 9945 29101 9979
rect 29101 9945 29135 9979
rect 29135 9945 29144 9979
rect 29092 9936 29144 9945
rect 29552 9911 29604 9920
rect 29552 9877 29561 9911
rect 29561 9877 29595 9911
rect 29595 9877 29604 9911
rect 29552 9868 29604 9877
rect 30472 9979 30524 9988
rect 30472 9945 30481 9979
rect 30481 9945 30515 9979
rect 30515 9945 30524 9979
rect 30472 9936 30524 9945
rect 30196 9868 30248 9920
rect 33508 10047 33560 10056
rect 33508 10013 33517 10047
rect 33517 10013 33551 10047
rect 33551 10013 33560 10047
rect 33508 10004 33560 10013
rect 36084 10047 36136 10056
rect 36084 10013 36093 10047
rect 36093 10013 36127 10047
rect 36127 10013 36136 10047
rect 36084 10004 36136 10013
rect 36452 10004 36504 10056
rect 37188 10072 37240 10124
rect 36636 10047 36688 10056
rect 36636 10013 36645 10047
rect 36645 10013 36679 10047
rect 36679 10013 36688 10047
rect 36636 10004 36688 10013
rect 37556 10047 37608 10056
rect 37556 10013 37565 10047
rect 37565 10013 37599 10047
rect 37599 10013 37608 10047
rect 37556 10004 37608 10013
rect 37648 10047 37700 10056
rect 37648 10013 37657 10047
rect 37657 10013 37691 10047
rect 37691 10013 37700 10047
rect 37648 10004 37700 10013
rect 38844 10047 38896 10056
rect 38844 10013 38853 10047
rect 38853 10013 38887 10047
rect 38887 10013 38896 10047
rect 38844 10004 38896 10013
rect 38936 10047 38988 10056
rect 38936 10013 38945 10047
rect 38945 10013 38979 10047
rect 38979 10013 38988 10047
rect 38936 10004 38988 10013
rect 40408 10047 40460 10056
rect 40408 10013 40417 10047
rect 40417 10013 40451 10047
rect 40451 10013 40460 10047
rect 40408 10004 40460 10013
rect 31944 9936 31996 9988
rect 33048 9936 33100 9988
rect 33232 9936 33284 9988
rect 37004 9936 37056 9988
rect 37464 9979 37516 9988
rect 37464 9945 37473 9979
rect 37473 9945 37507 9979
rect 37507 9945 37516 9979
rect 37464 9936 37516 9945
rect 32588 9868 32640 9920
rect 33876 9911 33928 9920
rect 33876 9877 33885 9911
rect 33885 9877 33919 9911
rect 33919 9877 33928 9911
rect 33876 9868 33928 9877
rect 37280 9868 37332 9920
rect 38660 9911 38712 9920
rect 38660 9877 38669 9911
rect 38669 9877 38703 9911
rect 38703 9877 38712 9911
rect 38660 9868 38712 9877
rect 39948 9936 40000 9988
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 5724 9664 5776 9716
rect 6828 9664 6880 9716
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 5632 9528 5684 9580
rect 5724 9528 5776 9580
rect 6184 9596 6236 9648
rect 6920 9528 6972 9580
rect 7380 9596 7432 9648
rect 23664 9664 23716 9716
rect 25504 9664 25556 9716
rect 28172 9664 28224 9716
rect 28724 9664 28776 9716
rect 31208 9707 31260 9716
rect 31208 9673 31217 9707
rect 31217 9673 31251 9707
rect 31251 9673 31260 9707
rect 31208 9664 31260 9673
rect 34796 9664 34848 9716
rect 11336 9596 11388 9648
rect 3424 9460 3476 9512
rect 4620 9460 4672 9512
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 1676 9324 1728 9376
rect 3424 9324 3476 9376
rect 6000 9392 6052 9444
rect 6276 9392 6328 9444
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 7288 9392 7340 9444
rect 5908 9324 5960 9376
rect 6368 9324 6420 9376
rect 6828 9324 6880 9376
rect 8484 9460 8536 9512
rect 8392 9392 8444 9444
rect 10140 9528 10192 9580
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 11520 9528 11572 9580
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 20076 9596 20128 9648
rect 22008 9596 22060 9648
rect 23204 9596 23256 9648
rect 23756 9596 23808 9648
rect 25688 9596 25740 9648
rect 26608 9596 26660 9648
rect 27344 9639 27396 9648
rect 27344 9605 27353 9639
rect 27353 9605 27387 9639
rect 27387 9605 27396 9639
rect 27344 9596 27396 9605
rect 28816 9596 28868 9648
rect 29552 9596 29604 9648
rect 19524 9528 19576 9580
rect 19708 9571 19760 9580
rect 19708 9537 19717 9571
rect 19717 9537 19751 9571
rect 19751 9537 19760 9571
rect 19708 9528 19760 9537
rect 19800 9571 19852 9580
rect 19800 9537 19809 9571
rect 19809 9537 19843 9571
rect 19843 9537 19852 9571
rect 19800 9528 19852 9537
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 21456 9571 21508 9580
rect 21456 9537 21465 9571
rect 21465 9537 21499 9571
rect 21499 9537 21508 9571
rect 21456 9528 21508 9537
rect 12164 9460 12216 9512
rect 21364 9460 21416 9512
rect 26700 9571 26752 9580
rect 26700 9537 26709 9571
rect 26709 9537 26743 9571
rect 26743 9537 26752 9571
rect 26700 9528 26752 9537
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 27988 9528 28040 9580
rect 30380 9528 30432 9580
rect 30840 9528 30892 9580
rect 31760 9596 31812 9648
rect 32404 9596 32456 9648
rect 33876 9639 33928 9648
rect 33876 9605 33885 9639
rect 33885 9605 33919 9639
rect 33919 9605 33928 9639
rect 33876 9596 33928 9605
rect 37648 9664 37700 9716
rect 38384 9664 38436 9716
rect 35992 9596 36044 9648
rect 36452 9639 36504 9648
rect 36452 9605 36461 9639
rect 36461 9605 36495 9639
rect 36495 9605 36504 9639
rect 36452 9596 36504 9605
rect 38660 9596 38712 9648
rect 21732 9460 21784 9512
rect 23296 9460 23348 9512
rect 23572 9503 23624 9512
rect 23572 9469 23581 9503
rect 23581 9469 23615 9503
rect 23615 9469 23624 9503
rect 23572 9460 23624 9469
rect 24584 9460 24636 9512
rect 12256 9392 12308 9444
rect 22284 9392 22336 9444
rect 25412 9392 25464 9444
rect 8024 9367 8076 9376
rect 8024 9333 8033 9367
rect 8033 9333 8067 9367
rect 8067 9333 8076 9367
rect 8024 9324 8076 9333
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10232 9367 10284 9376
rect 10232 9333 10241 9367
rect 10241 9333 10275 9367
rect 10275 9333 10284 9367
rect 10232 9324 10284 9333
rect 21640 9367 21692 9376
rect 21640 9333 21649 9367
rect 21649 9333 21683 9367
rect 21683 9333 21692 9367
rect 21640 9324 21692 9333
rect 22100 9324 22152 9376
rect 25136 9324 25188 9376
rect 28264 9392 28316 9444
rect 33048 9460 33100 9512
rect 32680 9392 32732 9444
rect 27620 9324 27672 9376
rect 29092 9324 29144 9376
rect 29828 9324 29880 9376
rect 30472 9324 30524 9376
rect 30840 9324 30892 9376
rect 33324 9324 33376 9376
rect 35532 9528 35584 9580
rect 36360 9571 36412 9580
rect 36360 9537 36369 9571
rect 36369 9537 36403 9571
rect 36403 9537 36412 9571
rect 36360 9528 36412 9537
rect 36544 9571 36596 9580
rect 36544 9537 36558 9571
rect 36558 9537 36592 9571
rect 36592 9537 36596 9571
rect 36544 9528 36596 9537
rect 36084 9460 36136 9512
rect 36176 9435 36228 9444
rect 36176 9401 36185 9435
rect 36185 9401 36219 9435
rect 36219 9401 36228 9435
rect 36176 9392 36228 9401
rect 36268 9324 36320 9376
rect 38660 9503 38712 9512
rect 38660 9469 38669 9503
rect 38669 9469 38703 9503
rect 38703 9469 38712 9503
rect 38660 9460 38712 9469
rect 40408 9503 40460 9512
rect 38568 9392 38620 9444
rect 40408 9469 40417 9503
rect 40417 9469 40451 9503
rect 40451 9469 40460 9503
rect 40408 9460 40460 9469
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2964 8984 3016 9036
rect 3148 9027 3200 9036
rect 3148 8993 3157 9027
rect 3157 8993 3191 9027
rect 3191 8993 3200 9027
rect 3976 9120 4028 9172
rect 6184 9120 6236 9172
rect 6552 9120 6604 9172
rect 7472 9120 7524 9172
rect 10232 9120 10284 9172
rect 12164 9163 12216 9172
rect 12164 9129 12173 9163
rect 12173 9129 12207 9163
rect 12207 9129 12216 9163
rect 12164 9120 12216 9129
rect 21732 9163 21784 9172
rect 21732 9129 21741 9163
rect 21741 9129 21775 9163
rect 21775 9129 21784 9163
rect 21732 9120 21784 9129
rect 3792 9052 3844 9104
rect 3148 8984 3200 8993
rect 5540 9027 5592 9036
rect 5540 8993 5549 9027
rect 5549 8993 5583 9027
rect 5583 8993 5592 9027
rect 5540 8984 5592 8993
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 6368 8984 6420 9036
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 1952 8780 2004 8832
rect 2504 8780 2556 8832
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 4712 8916 4764 8968
rect 3700 8848 3752 8900
rect 3884 8848 3936 8900
rect 5356 8916 5408 8968
rect 5816 8916 5868 8968
rect 6552 8916 6604 8968
rect 19524 9052 19576 9104
rect 22376 9120 22428 9172
rect 22744 9163 22796 9172
rect 22744 9129 22753 9163
rect 22753 9129 22787 9163
rect 22787 9129 22796 9163
rect 22744 9120 22796 9129
rect 23388 9120 23440 9172
rect 24584 9163 24636 9172
rect 24584 9129 24593 9163
rect 24593 9129 24627 9163
rect 24627 9129 24636 9163
rect 24584 9120 24636 9129
rect 32220 9163 32272 9172
rect 32220 9129 32229 9163
rect 32229 9129 32263 9163
rect 32263 9129 32272 9163
rect 32220 9120 32272 9129
rect 34336 9120 34388 9172
rect 36360 9120 36412 9172
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 8024 8984 8076 9036
rect 9312 8984 9364 9036
rect 11060 8984 11112 9036
rect 11520 8984 11572 9036
rect 11704 8984 11756 9036
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 8392 8916 8444 8968
rect 3332 8780 3384 8832
rect 6092 8848 6144 8900
rect 6736 8848 6788 8900
rect 9404 8916 9456 8968
rect 12808 8984 12860 9036
rect 10048 8848 10100 8900
rect 10324 8848 10376 8900
rect 12348 8916 12400 8968
rect 15292 8984 15344 9036
rect 15844 8984 15896 9036
rect 18328 8984 18380 9036
rect 19340 8984 19392 9036
rect 19708 8984 19760 9036
rect 22652 9052 22704 9104
rect 22928 9052 22980 9104
rect 24216 9052 24268 9104
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 19524 8959 19576 8968
rect 19524 8925 19533 8959
rect 19533 8925 19567 8959
rect 19567 8925 19576 8959
rect 19524 8916 19576 8925
rect 13176 8848 13228 8900
rect 20168 8916 20220 8968
rect 20352 8959 20404 8968
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 21640 8984 21692 9036
rect 22744 8984 22796 9036
rect 19800 8891 19852 8900
rect 19800 8857 19809 8891
rect 19809 8857 19843 8891
rect 19843 8857 19852 8891
rect 19800 8848 19852 8857
rect 19984 8848 20036 8900
rect 22008 8916 22060 8968
rect 22284 8916 22336 8968
rect 25136 9027 25188 9036
rect 25136 8993 25145 9027
rect 25145 8993 25179 9027
rect 25179 8993 25188 9027
rect 25136 8984 25188 8993
rect 25412 8984 25464 9036
rect 26424 8984 26476 9036
rect 30012 8984 30064 9036
rect 33232 9052 33284 9104
rect 33324 9052 33376 9104
rect 36728 9052 36780 9104
rect 24768 8959 24820 8968
rect 24768 8925 24777 8959
rect 24777 8925 24811 8959
rect 24811 8925 24820 8959
rect 24768 8916 24820 8925
rect 25044 8916 25096 8968
rect 5540 8780 5592 8832
rect 6552 8780 6604 8832
rect 9036 8780 9088 8832
rect 11244 8823 11296 8832
rect 11244 8789 11253 8823
rect 11253 8789 11287 8823
rect 11287 8789 11296 8823
rect 11244 8780 11296 8789
rect 11704 8780 11756 8832
rect 12992 8780 13044 8832
rect 19064 8823 19116 8832
rect 19064 8789 19073 8823
rect 19073 8789 19107 8823
rect 19107 8789 19116 8823
rect 19064 8780 19116 8789
rect 22468 8848 22520 8900
rect 23020 8848 23072 8900
rect 22100 8780 22152 8832
rect 25044 8780 25096 8832
rect 25688 8916 25740 8968
rect 29828 8959 29880 8968
rect 29828 8925 29837 8959
rect 29837 8925 29871 8959
rect 29871 8925 29880 8959
rect 29828 8916 29880 8925
rect 32956 8984 33008 9036
rect 32864 8959 32916 8968
rect 32864 8925 32873 8959
rect 32873 8925 32907 8959
rect 32907 8925 32916 8959
rect 32864 8916 32916 8925
rect 26792 8891 26844 8900
rect 26792 8857 26801 8891
rect 26801 8857 26835 8891
rect 26835 8857 26844 8891
rect 26792 8848 26844 8857
rect 26884 8848 26936 8900
rect 29920 8848 29972 8900
rect 30104 8891 30156 8900
rect 30104 8857 30113 8891
rect 30113 8857 30147 8891
rect 30147 8857 30156 8891
rect 30104 8848 30156 8857
rect 30288 8848 30340 8900
rect 31852 8848 31904 8900
rect 33232 8959 33284 8968
rect 33232 8925 33265 8959
rect 33265 8925 33284 8959
rect 33232 8916 33284 8925
rect 36176 8959 36228 8968
rect 36176 8925 36185 8959
rect 36185 8925 36219 8959
rect 36219 8925 36228 8959
rect 36176 8916 36228 8925
rect 36360 8984 36412 9036
rect 36452 8984 36504 9036
rect 37004 8984 37056 9036
rect 27160 8780 27212 8832
rect 29736 8780 29788 8832
rect 32588 8823 32640 8832
rect 32588 8789 32597 8823
rect 32597 8789 32631 8823
rect 32631 8789 32640 8823
rect 32588 8780 32640 8789
rect 37096 8959 37148 8968
rect 37096 8925 37105 8959
rect 37105 8925 37139 8959
rect 37139 8925 37148 8959
rect 37096 8916 37148 8925
rect 37280 8959 37332 8968
rect 37280 8925 37289 8959
rect 37289 8925 37323 8959
rect 37323 8925 37332 8959
rect 37280 8916 37332 8925
rect 37464 8959 37516 8968
rect 37464 8925 37473 8959
rect 37473 8925 37507 8959
rect 37507 8925 37516 8959
rect 37464 8916 37516 8925
rect 38016 8916 38068 8968
rect 38660 8959 38712 8968
rect 38660 8925 38669 8959
rect 38669 8925 38703 8959
rect 38703 8925 38712 8959
rect 38660 8916 38712 8925
rect 34244 8780 34296 8832
rect 35992 8823 36044 8832
rect 35992 8789 36001 8823
rect 36001 8789 36035 8823
rect 36035 8789 36044 8823
rect 35992 8780 36044 8789
rect 38936 8848 38988 8900
rect 37464 8780 37516 8832
rect 38476 8780 38528 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 6276 8576 6328 8628
rect 6644 8576 6696 8628
rect 3332 8508 3384 8560
rect 3700 8508 3752 8560
rect 5724 8508 5776 8560
rect 8760 8576 8812 8628
rect 9496 8576 9548 8628
rect 10140 8576 10192 8628
rect 8484 8508 8536 8560
rect 9036 8508 9088 8560
rect 10048 8508 10100 8560
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 6092 8440 6144 8492
rect 6460 8440 6512 8492
rect 7472 8440 7524 8492
rect 9312 8440 9364 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 10324 8440 10376 8492
rect 11888 8576 11940 8628
rect 13084 8576 13136 8628
rect 20352 8576 20404 8628
rect 22376 8619 22428 8628
rect 22376 8585 22385 8619
rect 22385 8585 22419 8619
rect 22419 8585 22428 8619
rect 22376 8576 22428 8585
rect 22468 8619 22520 8628
rect 22468 8585 22477 8619
rect 22477 8585 22511 8619
rect 22511 8585 22520 8619
rect 22468 8576 22520 8585
rect 22836 8576 22888 8628
rect 25136 8576 25188 8628
rect 25228 8576 25280 8628
rect 25412 8576 25464 8628
rect 26792 8576 26844 8628
rect 27160 8576 27212 8628
rect 12072 8508 12124 8560
rect 12164 8508 12216 8560
rect 12348 8508 12400 8560
rect 1952 8372 2004 8424
rect 2872 8415 2924 8424
rect 2872 8381 2881 8415
rect 2881 8381 2915 8415
rect 2915 8381 2924 8415
rect 2872 8372 2924 8381
rect 4804 8372 4856 8424
rect 8392 8372 8444 8424
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 11244 8440 11296 8492
rect 12992 8551 13044 8560
rect 12992 8517 13001 8551
rect 13001 8517 13035 8551
rect 13035 8517 13044 8551
rect 12992 8508 13044 8517
rect 14556 8508 14608 8560
rect 18144 8551 18196 8560
rect 18144 8517 18153 8551
rect 18153 8517 18187 8551
rect 18187 8517 18196 8551
rect 18144 8508 18196 8517
rect 20168 8508 20220 8560
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 23020 8440 23072 8492
rect 25136 8483 25188 8492
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 11428 8372 11480 8424
rect 11152 8304 11204 8356
rect 11336 8304 11388 8356
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 12440 8304 12492 8356
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 18420 8372 18472 8424
rect 19616 8415 19668 8424
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 19616 8372 19668 8381
rect 19984 8372 20036 8424
rect 22284 8372 22336 8424
rect 22744 8372 22796 8424
rect 24400 8372 24452 8424
rect 25228 8372 25280 8424
rect 25412 8483 25464 8492
rect 25412 8449 25421 8483
rect 25421 8449 25455 8483
rect 25455 8449 25464 8483
rect 25412 8440 25464 8449
rect 26332 8440 26384 8492
rect 26884 8440 26936 8492
rect 26976 8483 27028 8492
rect 26976 8449 26985 8483
rect 26985 8449 27019 8483
rect 27019 8449 27028 8483
rect 26976 8440 27028 8449
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 28816 8576 28868 8628
rect 29644 8576 29696 8628
rect 29736 8551 29788 8560
rect 29736 8517 29745 8551
rect 29745 8517 29779 8551
rect 29779 8517 29788 8551
rect 29736 8508 29788 8517
rect 31760 8440 31812 8492
rect 33048 8576 33100 8628
rect 34244 8551 34296 8560
rect 34244 8517 34253 8551
rect 34253 8517 34287 8551
rect 34287 8517 34296 8551
rect 34244 8508 34296 8517
rect 38016 8576 38068 8628
rect 38476 8576 38528 8628
rect 36268 8508 36320 8560
rect 38292 8508 38344 8560
rect 38936 8508 38988 8560
rect 36084 8440 36136 8492
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 4712 8279 4764 8288
rect 4712 8245 4721 8279
rect 4721 8245 4755 8279
rect 4755 8245 4764 8279
rect 4712 8236 4764 8245
rect 5356 8236 5408 8288
rect 6000 8279 6052 8288
rect 6000 8245 6009 8279
rect 6009 8245 6043 8279
rect 6043 8245 6052 8279
rect 6000 8236 6052 8245
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 6552 8236 6604 8245
rect 11244 8279 11296 8288
rect 11244 8245 11253 8279
rect 11253 8245 11287 8279
rect 11287 8245 11296 8279
rect 11244 8236 11296 8245
rect 12808 8236 12860 8288
rect 19340 8236 19392 8288
rect 24492 8304 24544 8356
rect 23756 8236 23808 8288
rect 24308 8236 24360 8288
rect 32404 8415 32456 8424
rect 32404 8381 32413 8415
rect 32413 8381 32447 8415
rect 32447 8381 32456 8415
rect 32404 8372 32456 8381
rect 33048 8372 33100 8424
rect 34336 8372 34388 8424
rect 36544 8440 36596 8492
rect 37096 8440 37148 8492
rect 37004 8372 37056 8424
rect 37464 8372 37516 8424
rect 39764 8415 39816 8424
rect 39764 8381 39773 8415
rect 39773 8381 39807 8415
rect 39807 8381 39816 8415
rect 39764 8372 39816 8381
rect 29736 8236 29788 8288
rect 30104 8279 30156 8288
rect 30104 8245 30113 8279
rect 30113 8245 30147 8279
rect 30147 8245 30156 8279
rect 30104 8236 30156 8245
rect 32864 8236 32916 8288
rect 37372 8347 37424 8356
rect 37372 8313 37381 8347
rect 37381 8313 37415 8347
rect 37415 8313 37424 8347
rect 37372 8304 37424 8313
rect 33876 8279 33928 8288
rect 33876 8245 33885 8279
rect 33885 8245 33919 8279
rect 33919 8245 33928 8279
rect 33876 8236 33928 8245
rect 35992 8279 36044 8288
rect 35992 8245 36001 8279
rect 36001 8245 36035 8279
rect 36035 8245 36044 8279
rect 35992 8236 36044 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2872 8032 2924 8084
rect 3884 8032 3936 8084
rect 4620 8032 4672 8084
rect 8300 8032 8352 8084
rect 8760 7896 8812 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 2964 7828 3016 7880
rect 3700 7828 3752 7880
rect 3884 7828 3936 7880
rect 1768 7760 1820 7812
rect 1952 7692 2004 7744
rect 3608 7803 3660 7812
rect 3608 7769 3617 7803
rect 3617 7769 3651 7803
rect 3651 7769 3660 7803
rect 4712 7828 4764 7880
rect 9680 8032 9732 8084
rect 10324 8075 10376 8084
rect 10324 8041 10333 8075
rect 10333 8041 10367 8075
rect 10367 8041 10376 8075
rect 10324 8032 10376 8041
rect 11152 8032 11204 8084
rect 11796 8032 11848 8084
rect 12164 8032 12216 8084
rect 19616 8032 19668 8084
rect 19800 8032 19852 8084
rect 9956 7964 10008 8016
rect 3608 7760 3660 7769
rect 8392 7803 8444 7812
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 8576 7803 8628 7812
rect 8576 7769 8601 7803
rect 8601 7769 8628 7803
rect 10140 7828 10192 7880
rect 11244 7964 11296 8016
rect 11888 7896 11940 7948
rect 15292 7896 15344 7948
rect 11244 7828 11296 7880
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 20352 7964 20404 8016
rect 24124 7964 24176 8016
rect 26792 8032 26844 8084
rect 26976 8075 27028 8084
rect 26976 8041 26985 8075
rect 26985 8041 27019 8075
rect 27019 8041 27028 8075
rect 26976 8032 27028 8041
rect 29828 8032 29880 8084
rect 32404 8032 32456 8084
rect 33232 8032 33284 8084
rect 38660 8032 38712 8084
rect 19064 7896 19116 7948
rect 19708 7896 19760 7948
rect 19800 7828 19852 7880
rect 22192 7896 22244 7948
rect 24400 7896 24452 7948
rect 24492 7939 24544 7948
rect 24492 7905 24501 7939
rect 24501 7905 24535 7939
rect 24535 7905 24544 7939
rect 24492 7896 24544 7905
rect 8576 7760 8628 7769
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 3792 7692 3844 7744
rect 3976 7735 4028 7744
rect 3976 7701 3985 7735
rect 3985 7701 4019 7735
rect 4019 7701 4028 7735
rect 3976 7692 4028 7701
rect 9036 7692 9088 7744
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 12808 7692 12860 7744
rect 13544 7803 13596 7812
rect 13544 7769 13553 7803
rect 13553 7769 13587 7803
rect 13587 7769 13596 7803
rect 13544 7760 13596 7769
rect 18696 7803 18748 7812
rect 18696 7769 18705 7803
rect 18705 7769 18739 7803
rect 18739 7769 18748 7803
rect 18696 7760 18748 7769
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 22928 7828 22980 7880
rect 20168 7803 20220 7812
rect 20168 7769 20177 7803
rect 20177 7769 20211 7803
rect 20211 7769 20220 7803
rect 20168 7760 20220 7769
rect 27160 7964 27212 8016
rect 25136 7896 25188 7948
rect 25320 7828 25372 7880
rect 14556 7692 14608 7744
rect 18052 7692 18104 7744
rect 20536 7735 20588 7744
rect 20536 7701 20545 7735
rect 20545 7701 20579 7735
rect 20579 7701 20588 7735
rect 20536 7692 20588 7701
rect 21272 7692 21324 7744
rect 24952 7735 25004 7744
rect 24952 7701 24961 7735
rect 24961 7701 24995 7735
rect 24995 7701 25004 7735
rect 24952 7692 25004 7701
rect 26792 7871 26844 7880
rect 26792 7837 26801 7871
rect 26801 7837 26835 7871
rect 26835 7837 26844 7871
rect 26792 7828 26844 7837
rect 29092 7939 29144 7948
rect 29092 7905 29101 7939
rect 29101 7905 29135 7939
rect 29135 7905 29144 7939
rect 29092 7896 29144 7905
rect 31668 7964 31720 8016
rect 31576 7939 31628 7948
rect 31576 7905 31585 7939
rect 31585 7905 31619 7939
rect 31619 7905 31628 7939
rect 31576 7896 31628 7905
rect 32220 7896 32272 7948
rect 26240 7760 26292 7812
rect 26424 7803 26476 7812
rect 26424 7769 26433 7803
rect 26433 7769 26467 7803
rect 26467 7769 26476 7803
rect 26424 7760 26476 7769
rect 27436 7760 27488 7812
rect 31300 7871 31352 7880
rect 31300 7837 31309 7871
rect 31309 7837 31343 7871
rect 31343 7837 31352 7871
rect 31300 7828 31352 7837
rect 29644 7760 29696 7812
rect 31024 7803 31076 7812
rect 31024 7769 31033 7803
rect 31033 7769 31067 7803
rect 31067 7769 31076 7803
rect 31024 7760 31076 7769
rect 32128 7828 32180 7880
rect 39764 7964 39816 8016
rect 33876 7939 33928 7948
rect 33876 7905 33885 7939
rect 33885 7905 33919 7939
rect 33919 7905 33928 7939
rect 33876 7896 33928 7905
rect 35348 7896 35400 7948
rect 32864 7828 32916 7880
rect 38936 7896 38988 7948
rect 38660 7871 38712 7880
rect 38660 7837 38669 7871
rect 38669 7837 38703 7871
rect 38703 7837 38712 7871
rect 38660 7828 38712 7837
rect 32772 7803 32824 7812
rect 32772 7769 32781 7803
rect 32781 7769 32815 7803
rect 32815 7769 32824 7803
rect 32772 7760 32824 7769
rect 35164 7760 35216 7812
rect 35900 7803 35952 7812
rect 35900 7769 35909 7803
rect 35909 7769 35943 7803
rect 35943 7769 35952 7803
rect 35900 7760 35952 7769
rect 36360 7760 36412 7812
rect 37372 7760 37424 7812
rect 28172 7692 28224 7744
rect 29460 7692 29512 7744
rect 32128 7692 32180 7744
rect 34888 7692 34940 7744
rect 36176 7692 36228 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 2872 7488 2924 7540
rect 3240 7488 3292 7540
rect 11244 7488 11296 7540
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 13544 7488 13596 7540
rect 18696 7488 18748 7540
rect 20168 7488 20220 7540
rect 22284 7488 22336 7540
rect 2228 7463 2280 7472
rect 2228 7429 2237 7463
rect 2237 7429 2271 7463
rect 2271 7429 2280 7463
rect 2228 7420 2280 7429
rect 12072 7420 12124 7472
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 3608 7352 3660 7404
rect 11612 7352 11664 7404
rect 12164 7352 12216 7404
rect 11888 7327 11940 7336
rect 11888 7293 11897 7327
rect 11897 7293 11931 7327
rect 11931 7293 11940 7327
rect 11888 7284 11940 7293
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 13176 7420 13228 7472
rect 19616 7420 19668 7472
rect 20352 7420 20404 7472
rect 21272 7463 21324 7472
rect 21272 7429 21281 7463
rect 21281 7429 21315 7463
rect 21315 7429 21324 7463
rect 21272 7420 21324 7429
rect 23204 7420 23256 7472
rect 23388 7420 23440 7472
rect 23756 7488 23808 7540
rect 27344 7488 27396 7540
rect 24308 7463 24360 7472
rect 24308 7429 24317 7463
rect 24317 7429 24351 7463
rect 24351 7429 24360 7463
rect 24308 7420 24360 7429
rect 24400 7463 24452 7472
rect 24400 7429 24409 7463
rect 24409 7429 24443 7463
rect 24443 7429 24452 7463
rect 24400 7420 24452 7429
rect 24768 7420 24820 7472
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24492 7395 24544 7404
rect 24492 7361 24501 7395
rect 24501 7361 24535 7395
rect 24535 7361 24544 7395
rect 24492 7352 24544 7361
rect 19984 7284 20036 7336
rect 20168 7327 20220 7336
rect 20168 7293 20177 7327
rect 20177 7293 20211 7327
rect 20211 7293 20220 7327
rect 20168 7284 20220 7293
rect 23296 7327 23348 7336
rect 23296 7293 23305 7327
rect 23305 7293 23339 7327
rect 23339 7293 23348 7327
rect 23296 7284 23348 7293
rect 23572 7327 23624 7336
rect 23572 7293 23581 7327
rect 23581 7293 23615 7327
rect 23615 7293 23624 7327
rect 23572 7284 23624 7293
rect 14556 7216 14608 7268
rect 20812 7216 20864 7268
rect 26056 7327 26108 7336
rect 26056 7293 26065 7327
rect 26065 7293 26099 7327
rect 26099 7293 26108 7327
rect 26056 7284 26108 7293
rect 27160 7420 27212 7472
rect 26240 7395 26292 7404
rect 26240 7361 26249 7395
rect 26249 7361 26283 7395
rect 26283 7361 26292 7395
rect 26240 7352 26292 7361
rect 27344 7352 27396 7404
rect 27804 7352 27856 7404
rect 28172 7463 28224 7472
rect 28172 7429 28181 7463
rect 28181 7429 28215 7463
rect 28215 7429 28224 7463
rect 28172 7420 28224 7429
rect 30472 7488 30524 7540
rect 31024 7488 31076 7540
rect 32404 7488 32456 7540
rect 32680 7488 32732 7540
rect 29092 7420 29144 7472
rect 31392 7420 31444 7472
rect 31576 7420 31628 7472
rect 34704 7531 34756 7540
rect 34704 7497 34713 7531
rect 34713 7497 34747 7531
rect 34747 7497 34756 7531
rect 34704 7488 34756 7497
rect 34980 7488 35032 7540
rect 35440 7488 35492 7540
rect 18696 7148 18748 7200
rect 21824 7191 21876 7200
rect 21824 7157 21833 7191
rect 21833 7157 21867 7191
rect 21867 7157 21876 7191
rect 21824 7148 21876 7157
rect 25412 7191 25464 7200
rect 25412 7157 25421 7191
rect 25421 7157 25455 7191
rect 25455 7157 25464 7191
rect 25412 7148 25464 7157
rect 26976 7191 27028 7200
rect 26976 7157 26985 7191
rect 26985 7157 27019 7191
rect 27019 7157 27028 7191
rect 26976 7148 27028 7157
rect 27620 7327 27672 7336
rect 27620 7293 27629 7327
rect 27629 7293 27663 7327
rect 27663 7293 27672 7327
rect 27620 7284 27672 7293
rect 27436 7216 27488 7268
rect 28908 7284 28960 7336
rect 29276 7327 29328 7336
rect 29276 7293 29285 7327
rect 29285 7293 29319 7327
rect 29319 7293 29328 7327
rect 29276 7284 29328 7293
rect 28448 7216 28500 7268
rect 29092 7148 29144 7200
rect 29460 7352 29512 7404
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 29736 7395 29788 7404
rect 29736 7361 29745 7395
rect 29745 7361 29779 7395
rect 29779 7361 29788 7395
rect 29736 7352 29788 7361
rect 30656 7352 30708 7404
rect 30932 7395 30984 7404
rect 30932 7361 30941 7395
rect 30941 7361 30975 7395
rect 30975 7361 30984 7395
rect 30932 7352 30984 7361
rect 31760 7352 31812 7404
rect 31024 7284 31076 7336
rect 31300 7327 31352 7336
rect 31300 7293 31309 7327
rect 31309 7293 31343 7327
rect 31343 7293 31352 7327
rect 31300 7284 31352 7293
rect 31392 7327 31444 7336
rect 31392 7293 31401 7327
rect 31401 7293 31435 7327
rect 31435 7293 31444 7327
rect 31392 7284 31444 7293
rect 34152 7395 34204 7404
rect 34152 7361 34161 7395
rect 34161 7361 34195 7395
rect 34195 7361 34204 7395
rect 34796 7420 34848 7472
rect 34152 7352 34204 7361
rect 34888 7395 34940 7404
rect 34888 7361 34897 7395
rect 34897 7361 34931 7395
rect 34931 7361 34940 7395
rect 34888 7352 34940 7361
rect 34980 7395 35032 7404
rect 34980 7361 34989 7395
rect 34989 7361 35023 7395
rect 35023 7361 35032 7395
rect 34980 7352 35032 7361
rect 35164 7352 35216 7404
rect 34336 7284 34388 7336
rect 35992 7463 36044 7472
rect 35992 7429 36001 7463
rect 36001 7429 36035 7463
rect 36035 7429 36044 7463
rect 35992 7420 36044 7429
rect 36544 7420 36596 7472
rect 37648 7488 37700 7540
rect 38936 7488 38988 7540
rect 41420 7488 41472 7540
rect 36360 7352 36412 7404
rect 36452 7395 36504 7404
rect 36452 7361 36461 7395
rect 36461 7361 36495 7395
rect 36495 7361 36504 7395
rect 36452 7352 36504 7361
rect 36544 7284 36596 7336
rect 36728 7395 36780 7404
rect 36728 7361 36737 7395
rect 36737 7361 36771 7395
rect 36771 7361 36780 7395
rect 36728 7352 36780 7361
rect 36820 7395 36872 7404
rect 36820 7361 36829 7395
rect 36829 7361 36863 7395
rect 36863 7361 36872 7395
rect 36820 7352 36872 7361
rect 37188 7352 37240 7404
rect 38200 7463 38252 7472
rect 38200 7429 38209 7463
rect 38209 7429 38243 7463
rect 38243 7429 38252 7463
rect 38200 7420 38252 7429
rect 38660 7463 38712 7472
rect 38660 7429 38669 7463
rect 38669 7429 38703 7463
rect 38703 7429 38712 7463
rect 38660 7420 38712 7429
rect 37004 7284 37056 7336
rect 31024 7148 31076 7200
rect 34336 7148 34388 7200
rect 36084 7216 36136 7268
rect 38752 7395 38804 7404
rect 38752 7361 38761 7395
rect 38761 7361 38795 7395
rect 38795 7361 38804 7395
rect 38752 7352 38804 7361
rect 39672 7352 39724 7404
rect 38844 7216 38896 7268
rect 35992 7148 36044 7200
rect 36636 7148 36688 7200
rect 37372 7148 37424 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2964 6944 3016 6996
rect 4436 6944 4488 6996
rect 5540 6944 5592 6996
rect 6092 6944 6144 6996
rect 8576 6987 8628 6996
rect 8576 6953 8585 6987
rect 8585 6953 8619 6987
rect 8619 6953 8628 6987
rect 8576 6944 8628 6953
rect 8760 6987 8812 6996
rect 8760 6953 8769 6987
rect 8769 6953 8803 6987
rect 8803 6953 8812 6987
rect 8760 6944 8812 6953
rect 3056 6876 3108 6928
rect 3792 6876 3844 6928
rect 2872 6783 2924 6792
rect 2872 6749 2881 6783
rect 2881 6749 2915 6783
rect 2915 6749 2924 6783
rect 2872 6740 2924 6749
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3240 6740 3292 6792
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 1676 6604 1728 6656
rect 3332 6604 3384 6656
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 6000 6876 6052 6928
rect 10876 6944 10928 6996
rect 11888 6987 11940 6996
rect 11888 6953 11897 6987
rect 11897 6953 11931 6987
rect 11931 6953 11940 6987
rect 11888 6944 11940 6953
rect 19616 6987 19668 6996
rect 19616 6953 19625 6987
rect 19625 6953 19659 6987
rect 19659 6953 19668 6987
rect 19616 6944 19668 6953
rect 20536 6944 20588 6996
rect 24124 6944 24176 6996
rect 25412 6944 25464 6996
rect 26976 6944 27028 6996
rect 27804 6944 27856 6996
rect 5908 6808 5960 6860
rect 6552 6808 6604 6860
rect 5724 6740 5776 6792
rect 6000 6672 6052 6724
rect 8392 6808 8444 6860
rect 9036 6851 9088 6860
rect 9036 6817 9045 6851
rect 9045 6817 9079 6851
rect 9079 6817 9088 6851
rect 9036 6808 9088 6817
rect 11060 6808 11112 6860
rect 18420 6808 18472 6860
rect 23572 6808 23624 6860
rect 26240 6851 26292 6860
rect 26240 6817 26249 6851
rect 26249 6817 26283 6851
rect 26283 6817 26292 6851
rect 26240 6808 26292 6817
rect 28724 6808 28776 6860
rect 7104 6740 7156 6792
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 9128 6740 9180 6792
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 5540 6604 5592 6656
rect 5724 6604 5776 6656
rect 6368 6604 6420 6656
rect 9312 6672 9364 6724
rect 10324 6672 10376 6724
rect 21180 6672 21232 6724
rect 21732 6715 21784 6724
rect 21732 6681 21741 6715
rect 21741 6681 21775 6715
rect 21775 6681 21784 6715
rect 21732 6672 21784 6681
rect 23388 6672 23440 6724
rect 7380 6604 7432 6656
rect 9404 6647 9456 6656
rect 9404 6613 9413 6647
rect 9413 6613 9447 6647
rect 9447 6613 9456 6647
rect 9404 6604 9456 6613
rect 22468 6604 22520 6656
rect 23020 6604 23072 6656
rect 23480 6604 23532 6656
rect 24492 6740 24544 6792
rect 24216 6715 24268 6724
rect 24216 6681 24225 6715
rect 24225 6681 24259 6715
rect 24259 6681 24268 6715
rect 24216 6672 24268 6681
rect 25596 6672 25648 6724
rect 27804 6672 27856 6724
rect 24952 6604 25004 6656
rect 29276 6944 29328 6996
rect 29644 6944 29696 6996
rect 30840 6944 30892 6996
rect 29460 6876 29512 6928
rect 30288 6876 30340 6928
rect 31760 6944 31812 6996
rect 32772 6944 32824 6996
rect 34704 6944 34756 6996
rect 36452 6987 36504 6996
rect 36452 6953 36461 6987
rect 36461 6953 36495 6987
rect 36495 6953 36504 6987
rect 36452 6944 36504 6953
rect 36820 6944 36872 6996
rect 31576 6919 31628 6928
rect 31576 6885 31585 6919
rect 31585 6885 31619 6919
rect 31619 6885 31628 6919
rect 31576 6876 31628 6885
rect 29000 6808 29052 6860
rect 29920 6783 29972 6792
rect 29920 6749 29929 6783
rect 29929 6749 29963 6783
rect 29963 6749 29972 6783
rect 29920 6740 29972 6749
rect 30472 6851 30524 6860
rect 30472 6817 30481 6851
rect 30481 6817 30515 6851
rect 30515 6817 30524 6851
rect 30472 6808 30524 6817
rect 30932 6808 30984 6860
rect 31208 6808 31260 6860
rect 31300 6740 31352 6792
rect 31392 6783 31444 6792
rect 31392 6749 31401 6783
rect 31401 6749 31435 6783
rect 31435 6749 31444 6783
rect 31392 6740 31444 6749
rect 34612 6740 34664 6792
rect 36728 6876 36780 6928
rect 36176 6808 36228 6860
rect 35992 6783 36044 6792
rect 35992 6749 36001 6783
rect 36001 6749 36035 6783
rect 36035 6749 36044 6783
rect 35992 6740 36044 6749
rect 36360 6783 36412 6792
rect 36360 6749 36369 6783
rect 36369 6749 36403 6783
rect 36403 6749 36412 6783
rect 36360 6740 36412 6749
rect 37004 6783 37056 6792
rect 37004 6749 37013 6783
rect 37013 6749 37047 6783
rect 37047 6749 37056 6783
rect 37004 6740 37056 6749
rect 37740 6783 37792 6792
rect 37740 6749 37749 6783
rect 37749 6749 37783 6783
rect 37783 6749 37792 6783
rect 37740 6740 37792 6749
rect 38844 6783 38896 6792
rect 38844 6749 38853 6783
rect 38853 6749 38887 6783
rect 38887 6749 38896 6783
rect 38844 6740 38896 6749
rect 29368 6672 29420 6724
rect 31024 6672 31076 6724
rect 34336 6672 34388 6724
rect 35440 6672 35492 6724
rect 30196 6647 30248 6656
rect 30196 6613 30205 6647
rect 30205 6613 30239 6647
rect 30239 6613 30248 6647
rect 30196 6604 30248 6613
rect 31300 6647 31352 6656
rect 31300 6613 31309 6647
rect 31309 6613 31343 6647
rect 31343 6613 31352 6647
rect 31300 6604 31352 6613
rect 34796 6604 34848 6656
rect 36268 6672 36320 6724
rect 38292 6715 38344 6724
rect 38292 6681 38301 6715
rect 38301 6681 38335 6715
rect 38335 6681 38344 6715
rect 38292 6672 38344 6681
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 1400 6400 1452 6452
rect 1676 6375 1728 6384
rect 1676 6341 1685 6375
rect 1685 6341 1719 6375
rect 1719 6341 1728 6375
rect 1676 6332 1728 6341
rect 2964 6332 3016 6384
rect 3240 6332 3292 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 3792 6332 3844 6384
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4620 6400 4672 6452
rect 8392 6400 8444 6452
rect 8852 6400 8904 6452
rect 10324 6400 10376 6452
rect 4436 6332 4488 6384
rect 4712 6332 4764 6384
rect 6368 6375 6420 6384
rect 6368 6341 6377 6375
rect 6377 6341 6411 6375
rect 6411 6341 6420 6375
rect 6368 6332 6420 6341
rect 6552 6375 6604 6384
rect 6552 6341 6593 6375
rect 6593 6341 6604 6375
rect 6552 6332 6604 6341
rect 7012 6332 7064 6384
rect 7380 6332 7432 6384
rect 8484 6332 8536 6384
rect 10508 6375 10560 6384
rect 10508 6341 10517 6375
rect 10517 6341 10551 6375
rect 10551 6341 10560 6375
rect 10508 6332 10560 6341
rect 10784 6332 10836 6384
rect 20168 6443 20220 6452
rect 20168 6409 20177 6443
rect 20177 6409 20211 6443
rect 20211 6409 20220 6443
rect 20168 6400 20220 6409
rect 23388 6400 23440 6452
rect 18696 6375 18748 6384
rect 18696 6341 18705 6375
rect 18705 6341 18739 6375
rect 18739 6341 18748 6375
rect 18696 6332 18748 6341
rect 20812 6375 20864 6384
rect 20812 6341 20821 6375
rect 20821 6341 20855 6375
rect 20855 6341 20864 6375
rect 20812 6332 20864 6341
rect 21180 6375 21232 6384
rect 21180 6341 21189 6375
rect 21189 6341 21223 6375
rect 21223 6341 21232 6375
rect 21180 6332 21232 6341
rect 9404 6264 9456 6316
rect 17960 6264 18012 6316
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 21824 6264 21876 6316
rect 23572 6332 23624 6384
rect 26056 6400 26108 6452
rect 27436 6400 27488 6452
rect 27804 6400 27856 6452
rect 25596 6332 25648 6384
rect 29552 6400 29604 6452
rect 28448 6375 28500 6384
rect 28448 6341 28457 6375
rect 28457 6341 28491 6375
rect 28491 6341 28500 6375
rect 28448 6332 28500 6341
rect 30196 6332 30248 6384
rect 30656 6332 30708 6384
rect 31852 6400 31904 6452
rect 33048 6400 33100 6452
rect 34336 6400 34388 6452
rect 32680 6375 32732 6384
rect 5908 6196 5960 6248
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 8944 6239 8996 6248
rect 8944 6205 8953 6239
rect 8953 6205 8987 6239
rect 8987 6205 8996 6239
rect 8944 6196 8996 6205
rect 23480 6239 23532 6248
rect 23480 6205 23489 6239
rect 23489 6205 23523 6239
rect 23523 6205 23532 6239
rect 23480 6196 23532 6205
rect 30840 6307 30892 6316
rect 30840 6273 30849 6307
rect 30849 6273 30883 6307
rect 30883 6273 30892 6307
rect 30840 6264 30892 6273
rect 31300 6264 31352 6316
rect 32680 6341 32689 6375
rect 32689 6341 32723 6375
rect 32723 6341 32732 6375
rect 32680 6332 32732 6341
rect 31668 6307 31720 6316
rect 31668 6273 31677 6307
rect 31677 6273 31711 6307
rect 31711 6273 31720 6307
rect 31668 6264 31720 6273
rect 31852 6264 31904 6316
rect 31944 6307 31996 6316
rect 31944 6273 31953 6307
rect 31953 6273 31987 6307
rect 31987 6273 31996 6307
rect 31944 6264 31996 6273
rect 32404 6307 32456 6316
rect 32404 6273 32413 6307
rect 32413 6273 32447 6307
rect 32447 6273 32456 6307
rect 32404 6264 32456 6273
rect 32588 6264 32640 6316
rect 35348 6332 35400 6384
rect 35440 6375 35492 6384
rect 35440 6341 35449 6375
rect 35449 6341 35483 6375
rect 35483 6341 35492 6375
rect 35440 6332 35492 6341
rect 36268 6400 36320 6452
rect 37740 6400 37792 6452
rect 3424 6060 3476 6112
rect 3516 6103 3568 6112
rect 3516 6069 3525 6103
rect 3525 6069 3559 6103
rect 3559 6069 3568 6103
rect 3516 6060 3568 6069
rect 3976 6060 4028 6112
rect 4068 6060 4120 6112
rect 10784 6128 10836 6180
rect 28724 6239 28776 6248
rect 28724 6205 28733 6239
rect 28733 6205 28767 6239
rect 28767 6205 28776 6239
rect 28724 6196 28776 6205
rect 29460 6239 29512 6248
rect 29460 6205 29469 6239
rect 29469 6205 29503 6239
rect 29503 6205 29512 6239
rect 29460 6196 29512 6205
rect 29920 6239 29972 6248
rect 29920 6205 29929 6239
rect 29929 6205 29963 6239
rect 29963 6205 29972 6239
rect 29920 6196 29972 6205
rect 30012 6196 30064 6248
rect 34704 6239 34756 6248
rect 34704 6205 34713 6239
rect 34713 6205 34747 6239
rect 34747 6205 34756 6239
rect 34704 6196 34756 6205
rect 5816 6060 5868 6112
rect 7472 6060 7524 6112
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 22652 6103 22704 6112
rect 22652 6069 22661 6103
rect 22661 6069 22695 6103
rect 22695 6069 22704 6103
rect 22652 6060 22704 6069
rect 28448 6060 28500 6112
rect 29092 6128 29144 6180
rect 31484 6128 31536 6180
rect 30472 6060 30524 6112
rect 30564 6103 30616 6112
rect 30564 6069 30573 6103
rect 30573 6069 30607 6103
rect 30607 6069 30616 6103
rect 30564 6060 30616 6069
rect 30748 6060 30800 6112
rect 32128 6103 32180 6112
rect 32128 6069 32137 6103
rect 32137 6069 32171 6103
rect 32171 6069 32180 6103
rect 32128 6060 32180 6069
rect 33232 6103 33284 6112
rect 33232 6069 33241 6103
rect 33241 6069 33275 6103
rect 33275 6069 33284 6103
rect 33232 6060 33284 6069
rect 41972 6264 42024 6316
rect 37464 6171 37516 6180
rect 37464 6137 37473 6171
rect 37473 6137 37507 6171
rect 37507 6137 37516 6171
rect 37464 6128 37516 6137
rect 38752 6128 38804 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 4068 5856 4120 5908
rect 4712 5856 4764 5908
rect 3884 5788 3936 5840
rect 1400 5720 1452 5772
rect 3240 5720 3292 5772
rect 3424 5720 3476 5772
rect 3056 5652 3108 5704
rect 4344 5720 4396 5772
rect 4620 5763 4672 5772
rect 4620 5729 4629 5763
rect 4629 5729 4663 5763
rect 4663 5729 4672 5763
rect 4620 5720 4672 5729
rect 6828 5720 6880 5772
rect 8944 5856 8996 5908
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 21732 5856 21784 5908
rect 23296 5856 23348 5908
rect 31300 5899 31352 5908
rect 31300 5865 31309 5899
rect 31309 5865 31343 5899
rect 31343 5865 31352 5899
rect 31300 5856 31352 5865
rect 32680 5856 32732 5908
rect 37004 5856 37056 5908
rect 41972 5899 42024 5908
rect 41972 5865 41981 5899
rect 41981 5865 42015 5899
rect 42015 5865 42024 5899
rect 41972 5856 42024 5865
rect 4804 5652 4856 5704
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 7196 5652 7248 5704
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 6184 5627 6236 5636
rect 6184 5593 6193 5627
rect 6193 5593 6227 5627
rect 6227 5593 6236 5627
rect 6184 5584 6236 5593
rect 10416 5720 10468 5772
rect 10784 5763 10836 5772
rect 10784 5729 10793 5763
rect 10793 5729 10827 5763
rect 10827 5729 10836 5763
rect 10784 5720 10836 5729
rect 11060 5763 11112 5772
rect 11060 5729 11069 5763
rect 11069 5729 11103 5763
rect 11103 5729 11112 5763
rect 11060 5720 11112 5729
rect 23756 5720 23808 5772
rect 28724 5720 28776 5772
rect 30564 5720 30616 5772
rect 32128 5720 32180 5772
rect 37372 5763 37424 5772
rect 37372 5729 37381 5763
rect 37381 5729 37415 5763
rect 37415 5729 37424 5763
rect 37372 5720 37424 5729
rect 37648 5763 37700 5772
rect 37648 5729 37657 5763
rect 37657 5729 37691 5763
rect 37691 5729 37700 5763
rect 37648 5720 37700 5729
rect 8852 5652 8904 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 22376 5695 22428 5704
rect 22376 5661 22385 5695
rect 22385 5661 22419 5695
rect 22419 5661 22428 5695
rect 22376 5652 22428 5661
rect 22836 5695 22888 5704
rect 22836 5661 22845 5695
rect 22845 5661 22879 5695
rect 22879 5661 22888 5695
rect 22836 5652 22888 5661
rect 24216 5652 24268 5704
rect 31208 5652 31260 5704
rect 33232 5652 33284 5704
rect 34152 5652 34204 5704
rect 10324 5584 10376 5636
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 8392 5516 8444 5568
rect 9496 5516 9548 5568
rect 22100 5584 22152 5636
rect 22652 5584 22704 5636
rect 29552 5584 29604 5636
rect 33048 5584 33100 5636
rect 38292 5584 38344 5636
rect 42064 5627 42116 5636
rect 42064 5593 42073 5627
rect 42073 5593 42107 5627
rect 42107 5593 42116 5627
rect 42064 5584 42116 5593
rect 22928 5516 22980 5568
rect 30748 5516 30800 5568
rect 30840 5516 30892 5568
rect 31668 5516 31720 5568
rect 34612 5516 34664 5568
rect 35256 5516 35308 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 5540 5355 5592 5364
rect 5540 5321 5549 5355
rect 5549 5321 5583 5355
rect 5583 5321 5592 5355
rect 5540 5312 5592 5321
rect 6000 5312 6052 5364
rect 9128 5312 9180 5364
rect 29920 5355 29972 5364
rect 29920 5321 29929 5355
rect 29929 5321 29963 5355
rect 29963 5321 29972 5355
rect 29920 5312 29972 5321
rect 31944 5312 31996 5364
rect 34704 5355 34756 5364
rect 34704 5321 34713 5355
rect 34713 5321 34747 5355
rect 34747 5321 34756 5355
rect 34704 5312 34756 5321
rect 3424 5244 3476 5296
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 4344 5244 4396 5296
rect 4712 5244 4764 5296
rect 9496 5244 9548 5296
rect 22192 5287 22244 5296
rect 22192 5253 22201 5287
rect 22201 5253 22235 5287
rect 22235 5253 22244 5287
rect 22192 5244 22244 5253
rect 22284 5287 22336 5296
rect 22284 5253 22293 5287
rect 22293 5253 22327 5287
rect 22327 5253 22336 5287
rect 22284 5244 22336 5253
rect 6828 5176 6880 5228
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 22468 5219 22520 5228
rect 22468 5185 22477 5219
rect 22477 5185 22511 5219
rect 22511 5185 22520 5219
rect 22468 5176 22520 5185
rect 28724 5244 28776 5296
rect 30656 5287 30708 5296
rect 30656 5253 30665 5287
rect 30665 5253 30699 5287
rect 30699 5253 30708 5287
rect 30656 5244 30708 5253
rect 29552 5176 29604 5228
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 6184 5151 6236 5160
rect 6184 5117 6193 5151
rect 6193 5117 6227 5151
rect 6227 5117 6236 5151
rect 6184 5108 6236 5117
rect 6368 5108 6420 5160
rect 6644 5108 6696 5160
rect 7656 5108 7708 5160
rect 8116 5151 8168 5160
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 28448 5151 28500 5160
rect 28448 5117 28457 5151
rect 28457 5117 28491 5151
rect 28491 5117 28500 5151
rect 28448 5108 28500 5117
rect 32772 5151 32824 5160
rect 32772 5117 32781 5151
rect 32781 5117 32815 5151
rect 32815 5117 32824 5151
rect 32772 5108 32824 5117
rect 32956 5108 33008 5160
rect 34612 5244 34664 5296
rect 36544 5244 36596 5296
rect 34796 5176 34848 5228
rect 35256 5219 35308 5228
rect 35256 5185 35265 5219
rect 35265 5185 35299 5219
rect 35299 5185 35308 5219
rect 35256 5176 35308 5185
rect 37464 5108 37516 5160
rect 22376 5040 22428 5092
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4804 4768 4856 4820
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 8116 4768 8168 4820
rect 32956 4811 33008 4820
rect 32956 4777 32965 4811
rect 32965 4777 32999 4811
rect 32999 4777 33008 4811
rect 32956 4768 33008 4777
rect 6000 4700 6052 4752
rect 8852 4632 8904 4684
rect 31208 4675 31260 4684
rect 31208 4641 31217 4675
rect 31217 4641 31251 4675
rect 31251 4641 31260 4675
rect 31208 4632 31260 4641
rect 31484 4675 31536 4684
rect 31484 4641 31493 4675
rect 31493 4641 31527 4675
rect 31527 4641 31536 4675
rect 31484 4632 31536 4641
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 6644 4564 6696 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 6092 4496 6144 4548
rect 10508 4496 10560 4548
rect 33048 4496 33100 4548
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 11428 2388 11480 2440
rect 11612 2252 11664 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 19982 45098 20038 45757
rect 20626 45098 20682 45757
rect 19982 45070 20300 45098
rect 19982 44957 20038 45070
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 20272 43450 20300 45070
rect 20548 45070 20682 45098
rect 20548 43450 20576 45070
rect 20626 44957 20682 45070
rect 21270 45098 21326 45757
rect 22558 45098 22614 45757
rect 23846 45098 23902 45757
rect 21270 45070 21588 45098
rect 21270 44957 21326 45070
rect 21560 43450 21588 45070
rect 22558 45070 22784 45098
rect 22558 44957 22614 45070
rect 22756 43450 22784 45070
rect 23846 45070 24072 45098
rect 23846 44957 23902 45070
rect 24044 43450 24072 45070
rect 35594 43548 35902 43557
rect 35594 43546 35600 43548
rect 35656 43546 35680 43548
rect 35736 43546 35760 43548
rect 35816 43546 35840 43548
rect 35896 43546 35902 43548
rect 35656 43494 35658 43546
rect 35838 43494 35840 43546
rect 35594 43492 35600 43494
rect 35656 43492 35680 43494
rect 35736 43492 35760 43494
rect 35816 43492 35840 43494
rect 35896 43492 35902 43494
rect 35594 43483 35902 43492
rect 20260 43444 20312 43450
rect 20260 43386 20312 43392
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 21548 43444 21600 43450
rect 21548 43386 21600 43392
rect 22744 43444 22796 43450
rect 22744 43386 22796 43392
rect 24032 43444 24084 43450
rect 24032 43386 24084 43392
rect 21640 43376 21692 43382
rect 21640 43318 21692 43324
rect 19892 43308 19944 43314
rect 19892 43250 19944 43256
rect 20904 43308 20956 43314
rect 20904 43250 20956 43256
rect 21088 43308 21140 43314
rect 21088 43250 21140 43256
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 17868 42832 17920 42838
rect 17868 42774 17920 42780
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 110 41984 166 41993
rect 110 41919 166 41928
rect 124 23186 152 41919
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 17132 41540 17184 41546
rect 17132 41482 17184 41488
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 17144 41274 17172 41482
rect 17132 41268 17184 41274
rect 17132 41210 17184 41216
rect 17224 41200 17276 41206
rect 17224 41142 17276 41148
rect 16856 41064 16908 41070
rect 16856 41006 16908 41012
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 16868 40730 16896 41006
rect 17040 40928 17092 40934
rect 17040 40870 17092 40876
rect 16856 40724 16908 40730
rect 16856 40666 16908 40672
rect 14740 40520 14792 40526
rect 14740 40462 14792 40468
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 14752 38962 14780 40462
rect 15660 40452 15712 40458
rect 15660 40394 15712 40400
rect 16120 40452 16172 40458
rect 16120 40394 16172 40400
rect 15672 40186 15700 40394
rect 15660 40180 15712 40186
rect 15660 40122 15712 40128
rect 16132 38962 16160 40394
rect 17052 40186 17080 40870
rect 17040 40180 17092 40186
rect 17040 40122 17092 40128
rect 17236 39098 17264 41142
rect 17776 41064 17828 41070
rect 17776 41006 17828 41012
rect 17880 41018 17908 42774
rect 19432 42628 19484 42634
rect 19432 42570 19484 42576
rect 19444 42226 19472 42570
rect 19524 42560 19576 42566
rect 19524 42502 19576 42508
rect 19616 42560 19668 42566
rect 19616 42502 19668 42508
rect 19800 42560 19852 42566
rect 19800 42502 19852 42508
rect 19432 42220 19484 42226
rect 19432 42162 19484 42168
rect 19444 41546 19472 42162
rect 19536 41682 19564 42502
rect 19628 41818 19656 42502
rect 19812 42294 19840 42502
rect 19800 42288 19852 42294
rect 19800 42230 19852 42236
rect 19616 41812 19668 41818
rect 19616 41754 19668 41760
rect 19524 41676 19576 41682
rect 19524 41618 19576 41624
rect 19432 41540 19484 41546
rect 19432 41482 19484 41488
rect 18604 41472 18656 41478
rect 18604 41414 18656 41420
rect 18616 41138 18644 41414
rect 18604 41132 18656 41138
rect 18604 41074 18656 41080
rect 18788 41132 18840 41138
rect 18788 41074 18840 41080
rect 18052 41064 18104 41070
rect 17880 41012 18052 41018
rect 17880 41006 18104 41012
rect 17788 40730 17816 41006
rect 17880 40990 18092 41006
rect 17776 40724 17828 40730
rect 17776 40666 17828 40672
rect 17408 40588 17460 40594
rect 17408 40530 17460 40536
rect 17316 39976 17368 39982
rect 17316 39918 17368 39924
rect 17224 39092 17276 39098
rect 17224 39034 17276 39040
rect 16580 39024 16632 39030
rect 16580 38966 16632 38972
rect 14740 38956 14792 38962
rect 14740 38898 14792 38904
rect 16120 38956 16172 38962
rect 16120 38898 16172 38904
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 14752 38654 14780 38898
rect 14752 38626 14872 38654
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 14844 38350 14872 38626
rect 14832 38344 14884 38350
rect 14832 38286 14884 38292
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 13360 37800 13412 37806
rect 13360 37742 13412 37748
rect 13636 37800 13688 37806
rect 13636 37742 13688 37748
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 13372 37262 13400 37742
rect 12900 37256 12952 37262
rect 12900 37198 12952 37204
rect 13360 37256 13412 37262
rect 13360 37198 13412 37204
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 5448 36848 5500 36854
rect 5448 36790 5500 36796
rect 7288 36848 7340 36854
rect 7288 36790 7340 36796
rect 3240 36712 3292 36718
rect 3240 36654 3292 36660
rect 4068 36712 4120 36718
rect 4068 36654 4120 36660
rect 3252 35766 3280 36654
rect 4080 36378 4108 36654
rect 4804 36576 4856 36582
rect 4804 36518 4856 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4068 36372 4120 36378
rect 4068 36314 4120 36320
rect 4620 36304 4672 36310
rect 4620 36246 4672 36252
rect 3976 36236 4028 36242
rect 3976 36178 4028 36184
rect 3884 36168 3936 36174
rect 3884 36110 3936 36116
rect 3896 35834 3924 36110
rect 3884 35828 3936 35834
rect 3884 35770 3936 35776
rect 3240 35760 3292 35766
rect 3240 35702 3292 35708
rect 2964 35624 3016 35630
rect 2964 35566 3016 35572
rect 2976 35290 3004 35566
rect 3332 35488 3384 35494
rect 3332 35430 3384 35436
rect 2964 35284 3016 35290
rect 2964 35226 3016 35232
rect 3344 35086 3372 35430
rect 3896 35086 3924 35770
rect 3332 35080 3384 35086
rect 3332 35022 3384 35028
rect 3516 35080 3568 35086
rect 3516 35022 3568 35028
rect 3884 35080 3936 35086
rect 3884 35022 3936 35028
rect 3528 34746 3556 35022
rect 3516 34740 3568 34746
rect 3516 34682 3568 34688
rect 3988 34542 4016 36178
rect 4252 36100 4304 36106
rect 4252 36042 4304 36048
rect 4264 35476 4292 36042
rect 4632 35766 4660 36246
rect 4712 36168 4764 36174
rect 4712 36110 4764 36116
rect 4620 35760 4672 35766
rect 4620 35702 4672 35708
rect 4724 35698 4752 36110
rect 4816 36038 4844 36518
rect 5460 36310 5488 36790
rect 7300 36310 7328 36790
rect 8116 36780 8168 36786
rect 8116 36722 8168 36728
rect 5448 36304 5500 36310
rect 5448 36246 5500 36252
rect 7288 36304 7340 36310
rect 7288 36246 7340 36252
rect 4804 36032 4856 36038
rect 4804 35974 4856 35980
rect 5356 36032 5408 36038
rect 5356 35974 5408 35980
rect 4816 35766 4844 35974
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4804 35760 4856 35766
rect 4804 35702 4856 35708
rect 4712 35692 4764 35698
rect 4712 35634 4764 35640
rect 4620 35624 4672 35630
rect 4620 35566 4672 35572
rect 4080 35448 4292 35476
rect 4080 35290 4108 35448
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 35284 4120 35290
rect 4068 35226 4120 35232
rect 4632 35170 4660 35566
rect 4540 35142 4660 35170
rect 4068 35080 4120 35086
rect 4540 35034 4568 35142
rect 4068 35022 4120 35028
rect 3240 34536 3292 34542
rect 3240 34478 3292 34484
rect 3976 34536 4028 34542
rect 3976 34478 4028 34484
rect 3252 33658 3280 34478
rect 3240 33652 3292 33658
rect 3240 33594 3292 33600
rect 3148 33584 3200 33590
rect 3148 33526 3200 33532
rect 1860 33516 1912 33522
rect 1860 33458 1912 33464
rect 2136 33516 2188 33522
rect 2136 33458 2188 33464
rect 1400 31136 1452 31142
rect 1400 31078 1452 31084
rect 1412 28626 1440 31078
rect 1872 30666 1900 33458
rect 2148 32774 2176 33458
rect 2228 33312 2280 33318
rect 2228 33254 2280 33260
rect 2412 33312 2464 33318
rect 2412 33254 2464 33260
rect 2136 32768 2188 32774
rect 2136 32710 2188 32716
rect 2240 32434 2268 33254
rect 2320 32836 2372 32842
rect 2320 32778 2372 32784
rect 2228 32428 2280 32434
rect 2228 32370 2280 32376
rect 2332 31396 2360 32778
rect 2424 32502 2452 33254
rect 3160 33017 3188 33526
rect 3146 33008 3202 33017
rect 2780 32972 2832 32978
rect 3146 32943 3202 32952
rect 2780 32914 2832 32920
rect 2504 32768 2556 32774
rect 2504 32710 2556 32716
rect 2412 32496 2464 32502
rect 2412 32438 2464 32444
rect 2516 32434 2544 32710
rect 2504 32428 2556 32434
rect 2504 32370 2556 32376
rect 2412 31408 2464 31414
rect 2332 31376 2412 31396
rect 2464 31376 2466 31385
rect 2332 31368 2410 31376
rect 2410 31311 2466 31320
rect 2044 31272 2096 31278
rect 2044 31214 2096 31220
rect 2056 30802 2084 31214
rect 2044 30796 2096 30802
rect 2044 30738 2096 30744
rect 1584 30660 1636 30666
rect 1584 30602 1636 30608
rect 1860 30660 1912 30666
rect 1860 30602 1912 30608
rect 2412 30660 2464 30666
rect 2412 30602 2464 30608
rect 1596 30190 1624 30602
rect 1872 30326 1900 30602
rect 2424 30394 2452 30602
rect 2412 30388 2464 30394
rect 2412 30330 2464 30336
rect 1860 30320 1912 30326
rect 1860 30262 1912 30268
rect 2516 30190 2544 32370
rect 2792 31736 2820 32914
rect 2872 32836 2924 32842
rect 2872 32778 2924 32784
rect 2884 32570 2912 32778
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 3160 32434 3188 32943
rect 3252 32570 3280 33594
rect 3608 33584 3660 33590
rect 3608 33526 3660 33532
rect 3332 33312 3384 33318
rect 3332 33254 3384 33260
rect 3344 32910 3372 33254
rect 3332 32904 3384 32910
rect 3332 32846 3384 32852
rect 3240 32564 3292 32570
rect 3240 32506 3292 32512
rect 3148 32428 3200 32434
rect 3148 32370 3200 32376
rect 3424 32428 3476 32434
rect 3424 32370 3476 32376
rect 3332 32292 3384 32298
rect 3332 32234 3384 32240
rect 3344 31890 3372 32234
rect 3332 31884 3384 31890
rect 3332 31826 3384 31832
rect 2872 31816 2924 31822
rect 2872 31758 2924 31764
rect 2700 31708 2820 31736
rect 2700 31142 2728 31708
rect 2778 31376 2834 31385
rect 2778 31311 2834 31320
rect 2688 31136 2740 31142
rect 2688 31078 2740 31084
rect 2596 30864 2648 30870
rect 2596 30806 2648 30812
rect 2608 30258 2636 30806
rect 2596 30252 2648 30258
rect 2596 30194 2648 30200
rect 1584 30184 1636 30190
rect 1584 30126 1636 30132
rect 2504 30184 2556 30190
rect 2504 30126 2556 30132
rect 2608 30122 2636 30194
rect 2596 30116 2648 30122
rect 2596 30058 2648 30064
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1780 29170 1808 29582
rect 1952 29572 2004 29578
rect 1952 29514 2004 29520
rect 1964 29170 1992 29514
rect 2412 29504 2464 29510
rect 2412 29446 2464 29452
rect 2424 29238 2452 29446
rect 2412 29232 2464 29238
rect 2412 29174 2464 29180
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1952 29164 2004 29170
rect 1952 29106 2004 29112
rect 2044 28960 2096 28966
rect 2044 28902 2096 28908
rect 2056 28626 2084 28902
rect 1400 28620 1452 28626
rect 1400 28562 1452 28568
rect 2044 28620 2096 28626
rect 2044 28562 2096 28568
rect 1412 28014 1440 28562
rect 2792 28558 2820 31311
rect 2884 30938 2912 31758
rect 3344 31754 3372 31826
rect 3160 31726 3372 31754
rect 3056 31340 3108 31346
rect 3056 31282 3108 31288
rect 2964 31136 3016 31142
rect 2964 31078 3016 31084
rect 2872 30932 2924 30938
rect 2872 30874 2924 30880
rect 2884 29646 2912 30874
rect 2976 30802 3004 31078
rect 3068 30802 3096 31282
rect 2964 30796 3016 30802
rect 2964 30738 3016 30744
rect 3056 30796 3108 30802
rect 3056 30738 3108 30744
rect 2964 30660 3016 30666
rect 3160 30648 3188 31726
rect 3332 31680 3384 31686
rect 3332 31622 3384 31628
rect 3240 31272 3292 31278
rect 3240 31214 3292 31220
rect 3252 30734 3280 31214
rect 3240 30728 3292 30734
rect 3240 30670 3292 30676
rect 3016 30620 3188 30648
rect 2964 30602 3016 30608
rect 3068 29646 3096 30620
rect 3252 30326 3280 30670
rect 3344 30598 3372 31622
rect 3436 30802 3464 32370
rect 3620 31754 3648 33526
rect 4080 32858 4108 35022
rect 4448 35006 4568 35034
rect 4724 35018 4752 35634
rect 4816 35578 4844 35702
rect 5368 35698 5396 35974
rect 4988 35692 5040 35698
rect 4988 35634 5040 35640
rect 5356 35692 5408 35698
rect 5356 35634 5408 35640
rect 4816 35550 4936 35578
rect 4908 35290 4936 35550
rect 5000 35494 5028 35634
rect 5460 35562 5488 36246
rect 6736 36168 6788 36174
rect 6736 36110 6788 36116
rect 7012 36168 7064 36174
rect 7012 36110 7064 36116
rect 5540 36100 5592 36106
rect 5540 36042 5592 36048
rect 5552 35766 5580 36042
rect 5540 35760 5592 35766
rect 5540 35702 5592 35708
rect 6748 35612 6776 36110
rect 6828 36032 6880 36038
rect 6828 35974 6880 35980
rect 6920 36032 6972 36038
rect 6920 35974 6972 35980
rect 6840 35766 6868 35974
rect 6828 35760 6880 35766
rect 6828 35702 6880 35708
rect 6828 35624 6880 35630
rect 6748 35584 6828 35612
rect 6828 35566 6880 35572
rect 5356 35556 5408 35562
rect 5356 35498 5408 35504
rect 5448 35556 5500 35562
rect 5448 35498 5500 35504
rect 4988 35488 5040 35494
rect 4988 35430 5040 35436
rect 5368 35442 5396 35498
rect 5540 35488 5592 35494
rect 4896 35284 4948 35290
rect 4896 35226 4948 35232
rect 5000 35018 5028 35430
rect 5368 35414 5488 35442
rect 5540 35430 5592 35436
rect 5356 35284 5408 35290
rect 5356 35226 5408 35232
rect 5264 35080 5316 35086
rect 5264 35022 5316 35028
rect 4712 35012 4764 35018
rect 4448 34950 4476 35006
rect 4712 34954 4764 34960
rect 4804 35012 4856 35018
rect 4804 34954 4856 34960
rect 4988 35012 5040 35018
rect 4988 34954 5040 34960
rect 4436 34944 4488 34950
rect 4436 34886 4488 34892
rect 4528 34944 4580 34950
rect 4528 34886 4580 34892
rect 4540 34678 4568 34886
rect 4528 34672 4580 34678
rect 4528 34614 4580 34620
rect 4540 34490 4568 34614
rect 4540 34462 4752 34490
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 33114 4660 33390
rect 4724 33130 4752 34462
rect 4816 34406 4844 34954
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4804 34400 4856 34406
rect 4804 34342 4856 34348
rect 5276 34066 5304 35022
rect 5368 34610 5396 35226
rect 5356 34604 5408 34610
rect 5356 34546 5408 34552
rect 5356 34468 5408 34474
rect 5356 34410 5408 34416
rect 5264 34060 5316 34066
rect 5264 34002 5316 34008
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 5276 33590 5304 34002
rect 5264 33584 5316 33590
rect 5264 33526 5316 33532
rect 5368 33522 5396 34410
rect 5460 33522 5488 35414
rect 5552 35154 5580 35430
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 6840 34950 6868 35566
rect 6932 35086 6960 35974
rect 7024 35222 7052 36110
rect 7104 36032 7156 36038
rect 7104 35974 7156 35980
rect 7116 35562 7144 35974
rect 7300 35698 7328 36246
rect 7288 35692 7340 35698
rect 7288 35634 7340 35640
rect 7380 35692 7432 35698
rect 7380 35634 7432 35640
rect 7104 35556 7156 35562
rect 7104 35498 7156 35504
rect 7012 35216 7064 35222
rect 7012 35158 7064 35164
rect 6920 35080 6972 35086
rect 6920 35022 6972 35028
rect 7116 35018 7144 35498
rect 7392 35290 7420 35634
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 7104 35012 7156 35018
rect 7104 34954 7156 34960
rect 7748 35012 7800 35018
rect 7748 34954 7800 34960
rect 6828 34944 6880 34950
rect 6828 34886 6880 34892
rect 6840 34610 6868 34886
rect 6828 34604 6880 34610
rect 6828 34546 6880 34552
rect 5632 34400 5684 34406
rect 5632 34342 5684 34348
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 5644 34202 5672 34342
rect 5632 34196 5684 34202
rect 5632 34138 5684 34144
rect 5908 33992 5960 33998
rect 5908 33934 5960 33940
rect 5724 33856 5776 33862
rect 5724 33798 5776 33804
rect 5356 33516 5408 33522
rect 5356 33458 5408 33464
rect 5448 33516 5500 33522
rect 5448 33458 5500 33464
rect 5540 33516 5592 33522
rect 5540 33458 5592 33464
rect 5172 33448 5224 33454
rect 5172 33390 5224 33396
rect 5264 33448 5316 33454
rect 5264 33390 5316 33396
rect 4988 33312 5040 33318
rect 4988 33254 5040 33260
rect 4620 33108 4672 33114
rect 4724 33102 4844 33130
rect 4620 33050 4672 33056
rect 4816 33046 4844 33102
rect 4804 33040 4856 33046
rect 4804 32982 4856 32988
rect 4712 32904 4764 32910
rect 3988 32842 4200 32858
rect 4448 32852 4712 32858
rect 4448 32846 4764 32852
rect 3988 32836 4212 32842
rect 3988 32830 4160 32836
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3712 31958 3740 32302
rect 3700 31952 3752 31958
rect 3700 31894 3752 31900
rect 3528 31726 3648 31754
rect 3424 30796 3476 30802
rect 3424 30738 3476 30744
rect 3332 30592 3384 30598
rect 3332 30534 3384 30540
rect 3240 30320 3292 30326
rect 3240 30262 3292 30268
rect 3252 30122 3280 30262
rect 3240 30116 3292 30122
rect 3240 30058 3292 30064
rect 3436 29782 3464 30738
rect 3424 29776 3476 29782
rect 3424 29718 3476 29724
rect 2872 29640 2924 29646
rect 2872 29582 2924 29588
rect 3056 29640 3108 29646
rect 3056 29582 3108 29588
rect 2872 29504 2924 29510
rect 2872 29446 2924 29452
rect 2780 28552 2832 28558
rect 2780 28494 2832 28500
rect 2792 28150 2820 28494
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 1400 28008 1452 28014
rect 1400 27950 1452 27956
rect 848 27872 900 27878
rect 846 27840 848 27849
rect 900 27840 902 27849
rect 846 27775 902 27784
rect 2792 27402 2820 28086
rect 2884 28014 2912 29446
rect 3068 29238 3096 29582
rect 3148 29572 3200 29578
rect 3148 29514 3200 29520
rect 3160 29238 3188 29514
rect 3056 29232 3108 29238
rect 3056 29174 3108 29180
rect 3148 29232 3200 29238
rect 3148 29174 3200 29180
rect 3068 28694 3096 29174
rect 3424 29028 3476 29034
rect 3424 28970 3476 28976
rect 3056 28688 3108 28694
rect 3056 28630 3108 28636
rect 3436 28626 3464 28970
rect 3424 28620 3476 28626
rect 3424 28562 3476 28568
rect 3528 28150 3556 31726
rect 3712 31346 3740 31894
rect 3988 31890 4016 32830
rect 4160 32778 4212 32784
rect 4448 32830 4752 32846
rect 4448 32774 4476 32830
rect 4436 32768 4488 32774
rect 4436 32710 4488 32716
rect 4528 32768 4580 32774
rect 4528 32710 4580 32716
rect 4540 32570 4568 32710
rect 4528 32564 4580 32570
rect 4528 32506 4580 32512
rect 4540 32314 4568 32506
rect 4724 32366 4752 32830
rect 4816 32434 4844 32982
rect 5000 32978 5028 33254
rect 5080 33108 5132 33114
rect 5080 33050 5132 33056
rect 4988 32972 5040 32978
rect 4988 32914 5040 32920
rect 5092 32842 5120 33050
rect 5080 32836 5132 32842
rect 5080 32778 5132 32784
rect 5184 32756 5212 33390
rect 5276 32824 5304 33390
rect 5368 32978 5396 33458
rect 5460 33114 5488 33458
rect 5448 33108 5500 33114
rect 5448 33050 5500 33056
rect 5460 33017 5488 33050
rect 5446 33008 5502 33017
rect 5356 32972 5408 32978
rect 5446 32943 5502 32952
rect 5356 32914 5408 32920
rect 5448 32836 5500 32842
rect 5276 32796 5396 32824
rect 5184 32728 5304 32756
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4988 32564 5040 32570
rect 4988 32506 5040 32512
rect 5000 32434 5028 32506
rect 4804 32428 4856 32434
rect 4804 32370 4856 32376
rect 4988 32428 5040 32434
rect 4988 32370 5040 32376
rect 4712 32360 4764 32366
rect 4540 32286 4660 32314
rect 4712 32302 4764 32308
rect 4068 32224 4120 32230
rect 4068 32166 4120 32172
rect 3976 31884 4028 31890
rect 3976 31826 4028 31832
rect 4080 31482 4108 32166
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 32026 4660 32286
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4068 31476 4120 31482
rect 4068 31418 4120 31424
rect 3700 31340 3752 31346
rect 3700 31282 3752 31288
rect 3608 30184 3660 30190
rect 3608 30126 3660 30132
rect 3620 29782 3648 30126
rect 3608 29776 3660 29782
rect 3608 29718 3660 29724
rect 3712 29730 3740 31282
rect 3884 30660 3936 30666
rect 3884 30602 3936 30608
rect 3896 30054 3924 30602
rect 4080 30394 4108 31418
rect 4724 31362 4752 32166
rect 4816 31822 4844 32370
rect 5000 32230 5028 32370
rect 5080 32360 5132 32366
rect 5276 32314 5304 32728
rect 5368 32502 5396 32796
rect 5448 32778 5500 32784
rect 5356 32496 5408 32502
rect 5356 32438 5408 32444
rect 5080 32302 5132 32308
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 5092 31822 5120 32302
rect 5184 32286 5304 32314
rect 5184 32026 5212 32286
rect 5264 32224 5316 32230
rect 5264 32166 5316 32172
rect 5172 32020 5224 32026
rect 5172 31962 5224 31968
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 5080 31816 5132 31822
rect 5080 31758 5132 31764
rect 5184 31686 5212 31962
rect 5276 31754 5304 32166
rect 5368 32026 5396 32438
rect 5460 32434 5488 32778
rect 5552 32774 5580 33458
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5540 32768 5592 32774
rect 5540 32710 5592 32716
rect 5448 32428 5500 32434
rect 5448 32370 5500 32376
rect 5540 32292 5592 32298
rect 5540 32234 5592 32240
rect 5356 32020 5408 32026
rect 5356 31962 5408 31968
rect 5356 31816 5408 31822
rect 5356 31758 5408 31764
rect 5264 31748 5316 31754
rect 5264 31690 5316 31696
rect 5172 31680 5224 31686
rect 5172 31622 5224 31628
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4724 31334 4844 31362
rect 4712 31272 4764 31278
rect 4712 31214 4764 31220
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30734 4660 31078
rect 4724 30938 4752 31214
rect 4712 30932 4764 30938
rect 4712 30874 4764 30880
rect 4816 30802 4844 31334
rect 5172 30932 5224 30938
rect 5172 30874 5224 30880
rect 4804 30796 4856 30802
rect 4804 30738 4856 30744
rect 5184 30734 5212 30874
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 5172 30728 5224 30734
rect 5224 30688 5304 30716
rect 5172 30670 5224 30676
rect 4068 30388 4120 30394
rect 4068 30330 4120 30336
rect 4632 30326 4660 30670
rect 4712 30660 4764 30666
rect 4712 30602 4764 30608
rect 4160 30320 4212 30326
rect 4160 30262 4212 30268
rect 4620 30320 4672 30326
rect 4620 30262 4672 30268
rect 4172 30138 4200 30262
rect 4080 30110 4200 30138
rect 4620 30116 4672 30122
rect 3884 30048 3936 30054
rect 3884 29990 3936 29996
rect 3620 29510 3648 29718
rect 3712 29702 3832 29730
rect 3804 29646 3832 29702
rect 3700 29640 3752 29646
rect 3700 29582 3752 29588
rect 3792 29640 3844 29646
rect 3792 29582 3844 29588
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 3620 29170 3648 29446
rect 3608 29164 3660 29170
rect 3608 29106 3660 29112
rect 3620 28762 3648 29106
rect 3608 28756 3660 28762
rect 3608 28698 3660 28704
rect 3712 28694 3740 29582
rect 3896 29578 3924 29990
rect 4080 29730 4108 30110
rect 4620 30058 4672 30064
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4080 29702 4200 29730
rect 3976 29640 4028 29646
rect 3976 29582 4028 29588
rect 3884 29572 3936 29578
rect 3884 29514 3936 29520
rect 3988 29510 4016 29582
rect 3792 29504 3844 29510
rect 3792 29446 3844 29452
rect 3976 29504 4028 29510
rect 3976 29446 4028 29452
rect 3804 29306 3832 29446
rect 3792 29300 3844 29306
rect 3792 29242 3844 29248
rect 3988 29034 4016 29446
rect 4172 29170 4200 29702
rect 4436 29708 4488 29714
rect 4436 29650 4488 29656
rect 4344 29640 4396 29646
rect 4344 29582 4396 29588
rect 4160 29164 4212 29170
rect 4160 29106 4212 29112
rect 4172 29050 4200 29106
rect 3976 29028 4028 29034
rect 3976 28970 4028 28976
rect 4080 29022 4200 29050
rect 3700 28688 3752 28694
rect 4080 28676 4108 29022
rect 4356 28966 4384 29582
rect 4448 29238 4476 29650
rect 4436 29232 4488 29238
rect 4436 29174 4488 29180
rect 4344 28960 4396 28966
rect 4344 28902 4396 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4080 28648 4200 28676
rect 3700 28630 3752 28636
rect 4172 28558 4200 28648
rect 4632 28558 4660 30058
rect 4724 29306 4752 30602
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5276 30376 5304 30688
rect 5184 30348 5304 30376
rect 5184 30122 5212 30348
rect 5262 30288 5318 30297
rect 5262 30223 5264 30232
rect 5316 30223 5318 30232
rect 5264 30194 5316 30200
rect 5172 30116 5224 30122
rect 5172 30058 5224 30064
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 4712 29096 4764 29102
rect 4712 29038 4764 29044
rect 4724 28642 4752 29038
rect 4816 28762 4844 29514
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5172 29164 5224 29170
rect 5092 29124 5172 29152
rect 5092 28966 5120 29124
rect 5172 29106 5224 29112
rect 5172 29028 5224 29034
rect 5172 28970 5224 28976
rect 5080 28960 5132 28966
rect 5080 28902 5132 28908
rect 4804 28756 4856 28762
rect 4804 28698 4856 28704
rect 5092 28694 5120 28902
rect 5080 28688 5132 28694
rect 4724 28626 4844 28642
rect 5080 28630 5132 28636
rect 4724 28620 4856 28626
rect 4724 28614 4804 28620
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 3608 28416 3660 28422
rect 3608 28358 3660 28364
rect 3620 28218 3648 28358
rect 4172 28218 4200 28494
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 4160 28212 4212 28218
rect 4160 28154 4212 28160
rect 3516 28144 3568 28150
rect 3516 28086 3568 28092
rect 2872 28008 2924 28014
rect 2872 27950 2924 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4160 27668 4212 27674
rect 4160 27610 4212 27616
rect 3608 27464 3660 27470
rect 3608 27406 3660 27412
rect 2780 27396 2832 27402
rect 2780 27338 2832 27344
rect 2792 27010 2820 27338
rect 2792 26982 3004 27010
rect 2780 26920 2832 26926
rect 2780 26862 2832 26868
rect 2792 26450 2820 26862
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 846 26072 902 26081
rect 846 26007 848 26016
rect 900 26007 902 26016
rect 848 25978 900 25984
rect 2792 25906 2820 26386
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 1306 25256 1362 25265
rect 1306 25191 1362 25200
rect 1320 24682 1348 25191
rect 1400 25152 1452 25158
rect 1400 25094 1452 25100
rect 1412 24818 1440 25094
rect 2700 24818 2728 25842
rect 2884 25362 2912 26726
rect 2976 26314 3004 26982
rect 3424 26852 3476 26858
rect 3424 26794 3476 26800
rect 3436 26586 3464 26794
rect 3424 26580 3476 26586
rect 3424 26522 3476 26528
rect 3516 26376 3568 26382
rect 3516 26318 3568 26324
rect 2964 26308 3016 26314
rect 2964 26250 3016 26256
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2976 25226 3004 26250
rect 3528 25362 3556 26318
rect 3620 25838 3648 27406
rect 4172 26994 4200 27610
rect 4632 27606 4660 28358
rect 4724 28014 4752 28614
rect 4804 28562 4856 28568
rect 5184 28558 5212 28970
rect 5172 28552 5224 28558
rect 5172 28494 5224 28500
rect 4804 28484 4856 28490
rect 4804 28426 4856 28432
rect 4816 28218 4844 28426
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4804 28212 4856 28218
rect 4804 28154 4856 28160
rect 5080 28212 5132 28218
rect 5080 28154 5132 28160
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4712 28008 4764 28014
rect 4712 27950 4764 27956
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4526 27432 4582 27441
rect 4526 27367 4528 27376
rect 4580 27367 4582 27376
rect 4528 27338 4580 27344
rect 4632 27282 4660 27542
rect 4540 27254 4660 27282
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4172 26874 4200 26930
rect 4080 26846 4200 26874
rect 4080 26466 4108 26846
rect 4540 26790 4568 27254
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 4528 26784 4580 26790
rect 4528 26726 4580 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4436 26580 4488 26586
rect 4436 26522 4488 26528
rect 4080 26438 4200 26466
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 3988 25906 4016 26318
rect 4172 26246 4200 26438
rect 4160 26240 4212 26246
rect 4160 26182 4212 26188
rect 4448 25906 4476 26522
rect 4528 26240 4580 26246
rect 4528 26182 4580 26188
rect 3792 25900 3844 25906
rect 3976 25900 4028 25906
rect 3844 25860 3976 25888
rect 3792 25842 3844 25848
rect 3976 25842 4028 25848
rect 4436 25900 4488 25906
rect 4436 25842 4488 25848
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3516 25356 3568 25362
rect 3516 25298 3568 25304
rect 2964 25220 3016 25226
rect 2964 25162 3016 25168
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 1308 24676 1360 24682
rect 1308 24618 1360 24624
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2136 24132 2188 24138
rect 2136 24074 2188 24080
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 23322 1440 23666
rect 2148 23594 2176 24074
rect 2516 23798 2544 24550
rect 2700 23798 2728 24754
rect 2976 24206 3004 25162
rect 3528 24274 3556 25298
rect 3804 24800 3832 25842
rect 4540 25770 4568 26182
rect 4632 25838 4660 27066
rect 4724 26858 4752 27950
rect 4816 27334 4844 28018
rect 5092 27878 5120 28154
rect 5172 27940 5224 27946
rect 5172 27882 5224 27888
rect 4988 27872 5040 27878
rect 4988 27814 5040 27820
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 5000 27674 5028 27814
rect 4988 27668 5040 27674
rect 4988 27610 5040 27616
rect 5184 27402 5212 27882
rect 5172 27396 5224 27402
rect 5172 27338 5224 27344
rect 4804 27328 4856 27334
rect 4804 27270 4856 27276
rect 4712 26852 4764 26858
rect 4712 26794 4764 26800
rect 4710 26616 4766 26625
rect 4710 26551 4712 26560
rect 4764 26551 4766 26560
rect 4712 26522 4764 26528
rect 4710 26344 4766 26353
rect 4816 26314 4844 27270
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4896 27124 4948 27130
rect 4896 27066 4948 27072
rect 4908 26382 4936 27066
rect 4988 26988 5040 26994
rect 4988 26930 5040 26936
rect 5000 26790 5028 26930
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 4896 26376 4948 26382
rect 5080 26376 5132 26382
rect 4896 26318 4948 26324
rect 5078 26344 5080 26353
rect 5132 26344 5134 26353
rect 4710 26279 4766 26288
rect 4804 26308 4856 26314
rect 4724 26042 4752 26279
rect 5078 26279 5134 26288
rect 4804 26250 4856 26256
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4712 25900 4764 25906
rect 4712 25842 4764 25848
rect 4620 25832 4672 25838
rect 4620 25774 4672 25780
rect 4528 25764 4580 25770
rect 4528 25706 4580 25712
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4436 25424 4488 25430
rect 4436 25366 4488 25372
rect 4448 24818 4476 25366
rect 4528 25288 4580 25294
rect 4528 25230 4580 25236
rect 4540 24818 4568 25230
rect 4632 24818 4660 25774
rect 4724 25702 4752 25842
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4724 24954 4752 25638
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 3884 24812 3936 24818
rect 3804 24772 3884 24800
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3804 24206 3832 24772
rect 3884 24754 3936 24760
rect 4436 24812 4488 24818
rect 4436 24754 4488 24760
rect 4528 24812 4580 24818
rect 4528 24754 4580 24760
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 3792 24200 3844 24206
rect 3792 24142 3844 24148
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2504 23792 2556 23798
rect 2504 23734 2556 23740
rect 2688 23792 2740 23798
rect 2688 23734 2740 23740
rect 2136 23588 2188 23594
rect 2136 23530 2188 23536
rect 1584 23520 1636 23526
rect 1584 23462 1636 23468
rect 2700 23474 2728 23734
rect 2792 23730 2820 24006
rect 3804 23730 3832 24142
rect 3988 23866 4016 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 2792 23610 2820 23666
rect 2792 23582 2912 23610
rect 4172 23594 4200 24006
rect 4264 23662 4292 24074
rect 4632 23798 4660 24074
rect 4724 24070 4752 24890
rect 4816 24206 4844 25774
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5276 24818 5304 30194
rect 5368 28762 5396 31758
rect 5552 31124 5580 32234
rect 5644 32026 5672 32846
rect 5632 32020 5684 32026
rect 5632 31962 5684 31968
rect 5632 31136 5684 31142
rect 5552 31096 5632 31124
rect 5632 31078 5684 31084
rect 5448 30864 5500 30870
rect 5448 30806 5500 30812
rect 5460 30326 5488 30806
rect 5644 30682 5672 31078
rect 5736 30870 5764 33798
rect 5920 33590 5948 33934
rect 6932 33930 6960 34342
rect 6920 33924 6972 33930
rect 6920 33866 6972 33872
rect 7012 33924 7064 33930
rect 7012 33866 7064 33872
rect 5908 33584 5960 33590
rect 5908 33526 5960 33532
rect 5816 33312 5868 33318
rect 5816 33254 5868 33260
rect 5828 32570 5856 33254
rect 5920 33046 5948 33526
rect 7024 33114 7052 33866
rect 7656 33584 7708 33590
rect 7656 33526 7708 33532
rect 6552 33108 6604 33114
rect 6552 33050 6604 33056
rect 7012 33108 7064 33114
rect 7012 33050 7064 33056
rect 5908 33040 5960 33046
rect 5960 33000 6040 33028
rect 5908 32982 5960 32988
rect 5908 32836 5960 32842
rect 5908 32778 5960 32784
rect 5816 32564 5868 32570
rect 5816 32506 5868 32512
rect 5920 31414 5948 32778
rect 6012 32366 6040 33000
rect 6276 32428 6328 32434
rect 6276 32370 6328 32376
rect 6460 32428 6512 32434
rect 6460 32370 6512 32376
rect 6000 32360 6052 32366
rect 6000 32302 6052 32308
rect 6092 32360 6144 32366
rect 6092 32302 6144 32308
rect 5908 31408 5960 31414
rect 5906 31376 5908 31385
rect 5960 31376 5962 31385
rect 5906 31311 5962 31320
rect 5816 30932 5868 30938
rect 5816 30874 5868 30880
rect 5724 30864 5776 30870
rect 5724 30806 5776 30812
rect 5828 30734 5856 30874
rect 5724 30728 5776 30734
rect 5644 30676 5724 30682
rect 5644 30670 5776 30676
rect 5816 30728 5868 30734
rect 5816 30670 5868 30676
rect 5644 30654 5764 30670
rect 5448 30320 5500 30326
rect 5448 30262 5500 30268
rect 5736 30190 5764 30654
rect 5816 30592 5868 30598
rect 5816 30534 5868 30540
rect 5828 30394 5856 30534
rect 5816 30388 5868 30394
rect 5816 30330 5868 30336
rect 6104 30274 6132 32302
rect 6288 31890 6316 32370
rect 6276 31884 6328 31890
rect 6276 31826 6328 31832
rect 6184 31476 6236 31482
rect 6184 31418 6236 31424
rect 6196 30734 6224 31418
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 5920 30246 6132 30274
rect 5540 30184 5592 30190
rect 5540 30126 5592 30132
rect 5632 30184 5684 30190
rect 5632 30126 5684 30132
rect 5724 30184 5776 30190
rect 5920 30138 5948 30246
rect 6288 30190 6316 31826
rect 6472 31822 6500 32370
rect 6564 32298 6592 33050
rect 7196 32836 7248 32842
rect 7196 32778 7248 32784
rect 7208 32570 7236 32778
rect 7196 32564 7248 32570
rect 7196 32506 7248 32512
rect 6552 32292 6604 32298
rect 6552 32234 6604 32240
rect 7668 32026 7696 33526
rect 7760 32910 7788 34954
rect 8128 33590 8156 36722
rect 12912 36242 12940 37198
rect 11060 36236 11112 36242
rect 11060 36178 11112 36184
rect 12900 36236 12952 36242
rect 12900 36178 12952 36184
rect 8668 36168 8720 36174
rect 8668 36110 8720 36116
rect 8392 36100 8444 36106
rect 8392 36042 8444 36048
rect 8404 35834 8432 36042
rect 8392 35828 8444 35834
rect 8392 35770 8444 35776
rect 8680 34626 8708 36110
rect 10324 36100 10376 36106
rect 10324 36042 10376 36048
rect 10416 36100 10468 36106
rect 10416 36042 10468 36048
rect 8944 36032 8996 36038
rect 8944 35974 8996 35980
rect 8760 35760 8812 35766
rect 8760 35702 8812 35708
rect 8772 35494 8800 35702
rect 8956 35630 8984 35974
rect 9036 35692 9088 35698
rect 9036 35634 9088 35640
rect 9956 35692 10008 35698
rect 9956 35634 10008 35640
rect 8944 35624 8996 35630
rect 8944 35566 8996 35572
rect 8760 35488 8812 35494
rect 8760 35430 8812 35436
rect 8956 35222 8984 35566
rect 9048 35222 9076 35634
rect 8944 35216 8996 35222
rect 8944 35158 8996 35164
rect 9036 35216 9088 35222
rect 9036 35158 9088 35164
rect 8956 34678 8984 35158
rect 9048 35018 9076 35158
rect 9036 35012 9088 35018
rect 9036 34954 9088 34960
rect 8312 34610 8708 34626
rect 8944 34672 8996 34678
rect 8944 34614 8996 34620
rect 8300 34604 8708 34610
rect 8352 34598 8708 34604
rect 8300 34546 8352 34552
rect 8312 34066 8340 34546
rect 9048 34542 9076 34954
rect 9312 34944 9364 34950
rect 9312 34886 9364 34892
rect 9324 34610 9352 34886
rect 9128 34604 9180 34610
rect 9128 34546 9180 34552
rect 9312 34604 9364 34610
rect 9312 34546 9364 34552
rect 9036 34536 9088 34542
rect 9036 34478 9088 34484
rect 8576 34468 8628 34474
rect 8576 34410 8628 34416
rect 8588 34202 8616 34410
rect 8576 34196 8628 34202
rect 8576 34138 8628 34144
rect 8588 34066 8616 34138
rect 9140 34134 9168 34546
rect 9588 34536 9640 34542
rect 9588 34478 9640 34484
rect 9128 34128 9180 34134
rect 9128 34070 9180 34076
rect 8300 34060 8352 34066
rect 8300 34002 8352 34008
rect 8576 34060 8628 34066
rect 8576 34002 8628 34008
rect 8312 33590 8340 34002
rect 8116 33584 8168 33590
rect 8116 33526 8168 33532
rect 8300 33584 8352 33590
rect 8300 33526 8352 33532
rect 8312 32978 8340 33526
rect 8588 33522 8616 34002
rect 8668 33924 8720 33930
rect 8668 33866 8720 33872
rect 8576 33516 8628 33522
rect 8576 33458 8628 33464
rect 8680 33454 8708 33866
rect 8944 33856 8996 33862
rect 8944 33798 8996 33804
rect 8668 33448 8720 33454
rect 8668 33390 8720 33396
rect 8300 32972 8352 32978
rect 8300 32914 8352 32920
rect 7748 32904 7800 32910
rect 7748 32846 7800 32852
rect 8116 32836 8168 32842
rect 8116 32778 8168 32784
rect 8128 32570 8156 32778
rect 8116 32564 8168 32570
rect 8116 32506 8168 32512
rect 7656 32020 7708 32026
rect 7656 31962 7708 31968
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6656 30802 6684 31758
rect 7012 31748 7064 31754
rect 7012 31690 7064 31696
rect 7024 31482 7052 31690
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 6644 30796 6696 30802
rect 6644 30738 6696 30744
rect 6552 30592 6604 30598
rect 6552 30534 6604 30540
rect 6564 30258 6592 30534
rect 6552 30252 6604 30258
rect 6552 30194 6604 30200
rect 5724 30126 5776 30132
rect 5448 30116 5500 30122
rect 5448 30058 5500 30064
rect 5460 29646 5488 30058
rect 5448 29640 5500 29646
rect 5448 29582 5500 29588
rect 5356 28756 5408 28762
rect 5356 28698 5408 28704
rect 5356 28484 5408 28490
rect 5356 28426 5408 28432
rect 5368 28218 5396 28426
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 5356 27396 5408 27402
rect 5356 27338 5408 27344
rect 5368 26586 5396 27338
rect 5460 27130 5488 29582
rect 5552 29306 5580 30126
rect 5644 29850 5672 30126
rect 5632 29844 5684 29850
rect 5632 29786 5684 29792
rect 5736 29782 5764 30126
rect 5828 30110 5948 30138
rect 6000 30184 6052 30190
rect 6000 30126 6052 30132
rect 6184 30184 6236 30190
rect 6184 30126 6236 30132
rect 6276 30184 6328 30190
rect 6276 30126 6328 30132
rect 5828 30054 5856 30110
rect 5816 30048 5868 30054
rect 5816 29990 5868 29996
rect 5908 30048 5960 30054
rect 5908 29990 5960 29996
rect 5724 29776 5776 29782
rect 5724 29718 5776 29724
rect 5920 29714 5948 29990
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5540 29300 5592 29306
rect 5540 29242 5592 29248
rect 5644 29186 5672 29582
rect 5724 29504 5776 29510
rect 5724 29446 5776 29452
rect 5736 29306 5764 29446
rect 5724 29300 5776 29306
rect 5724 29242 5776 29248
rect 5644 29170 5764 29186
rect 5828 29170 5856 29582
rect 5644 29164 5776 29170
rect 5644 29158 5724 29164
rect 5724 29106 5776 29112
rect 5816 29164 5868 29170
rect 5816 29106 5868 29112
rect 5736 29034 5764 29106
rect 5724 29028 5776 29034
rect 5724 28970 5776 28976
rect 5632 28960 5684 28966
rect 5632 28902 5684 28908
rect 5540 28688 5592 28694
rect 5540 28630 5592 28636
rect 5552 28558 5580 28630
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5552 27946 5580 28494
rect 5644 28218 5672 28902
rect 6012 28762 6040 30126
rect 6092 29776 6144 29782
rect 6092 29718 6144 29724
rect 6000 28756 6052 28762
rect 6000 28698 6052 28704
rect 5632 28212 5684 28218
rect 5632 28154 5684 28160
rect 5724 28144 5776 28150
rect 5724 28086 5776 28092
rect 5540 27940 5592 27946
rect 5540 27882 5592 27888
rect 5736 27674 5764 28086
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5724 27668 5776 27674
rect 5724 27610 5776 27616
rect 5736 27554 5764 27610
rect 5552 27526 5764 27554
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5552 26858 5580 27526
rect 5722 27432 5778 27441
rect 5722 27367 5724 27376
rect 5776 27367 5778 27376
rect 5724 27338 5776 27344
rect 5736 27130 5764 27338
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 5632 26920 5684 26926
rect 5632 26862 5684 26868
rect 5540 26852 5592 26858
rect 5540 26794 5592 26800
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 5354 26480 5410 26489
rect 5354 26415 5410 26424
rect 5368 25906 5396 26415
rect 5460 26330 5488 26726
rect 5540 26376 5592 26382
rect 5460 26324 5540 26330
rect 5460 26318 5592 26324
rect 5460 26302 5580 26318
rect 5448 26240 5500 26246
rect 5448 26182 5500 26188
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 5368 24886 5396 25842
rect 5460 25430 5488 26182
rect 5644 25770 5672 26862
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 5736 26382 5764 26794
rect 5828 26489 5856 27814
rect 6012 26625 6040 28698
rect 6104 28150 6132 29718
rect 6092 28144 6144 28150
rect 6092 28086 6144 28092
rect 6196 27878 6224 30126
rect 6460 30048 6512 30054
rect 6460 29990 6512 29996
rect 6472 29714 6500 29990
rect 6564 29782 6592 30194
rect 6552 29776 6604 29782
rect 6552 29718 6604 29724
rect 6656 29714 6684 30738
rect 7668 30297 7696 31962
rect 8128 31414 8156 32506
rect 8312 31890 8340 32914
rect 8680 32366 8708 33390
rect 8760 33312 8812 33318
rect 8760 33254 8812 33260
rect 8772 32910 8800 33254
rect 8760 32904 8812 32910
rect 8760 32846 8812 32852
rect 8956 32842 8984 33798
rect 9140 33454 9168 34070
rect 9600 33590 9628 34478
rect 9680 34400 9732 34406
rect 9680 34342 9732 34348
rect 9692 34202 9720 34342
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 9784 33998 9812 34138
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9864 33992 9916 33998
rect 9968 33980 9996 35634
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 10048 34400 10100 34406
rect 10048 34342 10100 34348
rect 10060 34066 10088 34342
rect 10048 34060 10100 34066
rect 10048 34002 10100 34008
rect 9916 33952 9996 33980
rect 9864 33934 9916 33940
rect 9588 33584 9640 33590
rect 9588 33526 9640 33532
rect 9128 33448 9180 33454
rect 9128 33390 9180 33396
rect 9496 33448 9548 33454
rect 9496 33390 9548 33396
rect 9508 33114 9536 33390
rect 9600 33114 9628 33526
rect 9496 33108 9548 33114
rect 9496 33050 9548 33056
rect 9588 33108 9640 33114
rect 9588 33050 9640 33056
rect 9968 32910 9996 33952
rect 10140 33856 10192 33862
rect 10140 33798 10192 33804
rect 10152 32910 10180 33798
rect 10244 32978 10272 35430
rect 10336 34898 10364 36042
rect 10428 35834 10456 36042
rect 10416 35828 10468 35834
rect 10416 35770 10468 35776
rect 11072 35766 11100 36178
rect 11060 35760 11112 35766
rect 11060 35702 11112 35708
rect 10416 35692 10468 35698
rect 10416 35634 10468 35640
rect 10508 35692 10560 35698
rect 10508 35634 10560 35640
rect 10784 35692 10836 35698
rect 10784 35634 10836 35640
rect 10876 35692 10928 35698
rect 10876 35634 10928 35640
rect 10428 35494 10456 35634
rect 10416 35488 10468 35494
rect 10416 35430 10468 35436
rect 10520 35290 10548 35634
rect 10600 35488 10652 35494
rect 10600 35430 10652 35436
rect 10508 35284 10560 35290
rect 10508 35226 10560 35232
rect 10612 35086 10640 35430
rect 10796 35222 10824 35634
rect 10784 35216 10836 35222
rect 10784 35158 10836 35164
rect 10600 35080 10652 35086
rect 10600 35022 10652 35028
rect 10888 34950 10916 35634
rect 12256 35624 12308 35630
rect 12256 35566 12308 35572
rect 12440 35624 12492 35630
rect 12440 35566 12492 35572
rect 12268 35290 12296 35566
rect 12256 35284 12308 35290
rect 12256 35226 12308 35232
rect 12452 35086 12480 35566
rect 12624 35488 12676 35494
rect 12544 35448 12624 35476
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 10876 34944 10928 34950
rect 10336 34870 10640 34898
rect 10876 34886 10928 34892
rect 10612 34678 10640 34870
rect 11428 34740 11480 34746
rect 11428 34682 11480 34688
rect 10600 34672 10652 34678
rect 10600 34614 10652 34620
rect 10612 34202 10640 34614
rect 11440 34542 11468 34682
rect 11428 34536 11480 34542
rect 11428 34478 11480 34484
rect 11440 34202 11468 34478
rect 10600 34196 10652 34202
rect 10600 34138 10652 34144
rect 11152 34196 11204 34202
rect 11152 34138 11204 34144
rect 11428 34196 11480 34202
rect 11428 34138 11480 34144
rect 10612 33522 10640 34138
rect 10968 34060 11020 34066
rect 10968 34002 11020 34008
rect 10980 33658 11008 34002
rect 11060 33992 11112 33998
rect 11060 33934 11112 33940
rect 10968 33652 11020 33658
rect 10968 33594 11020 33600
rect 10600 33516 10652 33522
rect 10600 33458 10652 33464
rect 10980 33318 11008 33594
rect 11072 33386 11100 33934
rect 11164 33522 11192 34138
rect 11336 33856 11388 33862
rect 11336 33798 11388 33804
rect 11348 33522 11376 33798
rect 12452 33658 12480 35022
rect 12544 33930 12572 35448
rect 12624 35430 12676 35436
rect 12912 34542 12940 36178
rect 13452 36168 13504 36174
rect 13452 36110 13504 36116
rect 13464 35766 13492 36110
rect 13452 35760 13504 35766
rect 13452 35702 13504 35708
rect 13360 35692 13412 35698
rect 13360 35634 13412 35640
rect 13372 35562 13400 35634
rect 13360 35556 13412 35562
rect 13360 35498 13412 35504
rect 13176 35284 13228 35290
rect 13176 35226 13228 35232
rect 13188 35018 13216 35226
rect 13372 35018 13400 35498
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 13360 35012 13412 35018
rect 13360 34954 13412 34960
rect 13464 34678 13492 35702
rect 13648 35290 13676 37742
rect 14844 37262 14872 38286
rect 16132 38282 16160 38898
rect 16488 38888 16540 38894
rect 16488 38830 16540 38836
rect 16500 38554 16528 38830
rect 16488 38548 16540 38554
rect 16488 38490 16540 38496
rect 16592 38486 16620 38966
rect 16580 38480 16632 38486
rect 16580 38422 16632 38428
rect 15108 38276 15160 38282
rect 15108 38218 15160 38224
rect 16120 38276 16172 38282
rect 16120 38218 16172 38224
rect 15120 38010 15148 38218
rect 15108 38004 15160 38010
rect 15108 37946 15160 37952
rect 15752 37868 15804 37874
rect 15752 37810 15804 37816
rect 16028 37868 16080 37874
rect 16132 37856 16160 38218
rect 16080 37828 16160 37856
rect 16212 37868 16264 37874
rect 16028 37810 16080 37816
rect 16212 37810 16264 37816
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 15108 37188 15160 37194
rect 15108 37130 15160 37136
rect 15016 36576 15068 36582
rect 15016 36518 15068 36524
rect 13912 36372 13964 36378
rect 13912 36314 13964 36320
rect 13728 36032 13780 36038
rect 13728 35974 13780 35980
rect 13740 35766 13768 35974
rect 13728 35760 13780 35766
rect 13728 35702 13780 35708
rect 13636 35284 13688 35290
rect 13636 35226 13688 35232
rect 13820 35148 13872 35154
rect 13820 35090 13872 35096
rect 13452 34672 13504 34678
rect 13452 34614 13504 34620
rect 12900 34536 12952 34542
rect 12900 34478 12952 34484
rect 12912 34066 12940 34478
rect 13464 34066 13492 34614
rect 13832 34202 13860 35090
rect 13924 35018 13952 36314
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 14464 36168 14516 36174
rect 14464 36110 14516 36116
rect 14108 35834 14136 36110
rect 14188 36032 14240 36038
rect 14188 35974 14240 35980
rect 14096 35828 14148 35834
rect 14096 35770 14148 35776
rect 14200 35698 14228 35974
rect 14476 35834 14504 36110
rect 14464 35828 14516 35834
rect 14464 35770 14516 35776
rect 14476 35698 14504 35770
rect 15028 35766 15056 36518
rect 15016 35760 15068 35766
rect 15016 35702 15068 35708
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 14188 35692 14240 35698
rect 14188 35634 14240 35640
rect 14464 35692 14516 35698
rect 14464 35634 14516 35640
rect 13912 35012 13964 35018
rect 13912 34954 13964 34960
rect 14108 34950 14136 35634
rect 14200 35222 14228 35634
rect 15120 35630 15148 37130
rect 15568 36712 15620 36718
rect 15568 36654 15620 36660
rect 15292 36576 15344 36582
rect 15292 36518 15344 36524
rect 15304 36106 15332 36518
rect 15292 36100 15344 36106
rect 15292 36042 15344 36048
rect 15108 35624 15160 35630
rect 15108 35566 15160 35572
rect 15580 35290 15608 36654
rect 15764 36106 15792 37810
rect 16224 37466 16252 37810
rect 16592 37806 16620 38422
rect 17132 38208 17184 38214
rect 17132 38150 17184 38156
rect 16856 37936 16908 37942
rect 16856 37878 16908 37884
rect 16580 37800 16632 37806
rect 16580 37742 16632 37748
rect 16212 37460 16264 37466
rect 16212 37402 16264 37408
rect 16580 37256 16632 37262
rect 16580 37198 16632 37204
rect 16028 37120 16080 37126
rect 16028 37062 16080 37068
rect 15936 36780 15988 36786
rect 15936 36722 15988 36728
rect 15752 36100 15804 36106
rect 15752 36042 15804 36048
rect 15764 35766 15792 36042
rect 15948 36038 15976 36722
rect 15936 36032 15988 36038
rect 15936 35974 15988 35980
rect 15752 35760 15804 35766
rect 15752 35702 15804 35708
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 14188 35216 14240 35222
rect 14188 35158 14240 35164
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14096 34944 14148 34950
rect 14096 34886 14148 34892
rect 14464 34944 14516 34950
rect 14464 34886 14516 34892
rect 13912 34400 13964 34406
rect 13912 34342 13964 34348
rect 13924 34202 13952 34342
rect 13820 34196 13872 34202
rect 13820 34138 13872 34144
rect 13912 34196 13964 34202
rect 13912 34138 13964 34144
rect 12900 34060 12952 34066
rect 12900 34002 12952 34008
rect 13452 34060 13504 34066
rect 13452 34002 13504 34008
rect 14476 33998 14504 34886
rect 14556 34536 14608 34542
rect 14556 34478 14608 34484
rect 14568 33998 14596 34478
rect 14660 34066 14688 35022
rect 15764 34678 15792 35702
rect 15948 35154 15976 35974
rect 15936 35148 15988 35154
rect 15936 35090 15988 35096
rect 16040 35086 16068 37062
rect 16488 36304 16540 36310
rect 16488 36246 16540 36252
rect 16028 35080 16080 35086
rect 16028 35022 16080 35028
rect 15844 34944 15896 34950
rect 15844 34886 15896 34892
rect 15752 34672 15804 34678
rect 15752 34614 15804 34620
rect 14648 34060 14700 34066
rect 14648 34002 14700 34008
rect 15856 33998 15884 34886
rect 16040 34746 16068 35022
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 16396 34604 16448 34610
rect 16396 34546 16448 34552
rect 16408 34202 16436 34546
rect 16396 34196 16448 34202
rect 16396 34138 16448 34144
rect 16500 34066 16528 36246
rect 16488 34060 16540 34066
rect 16488 34002 16540 34008
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14556 33992 14608 33998
rect 14556 33934 14608 33940
rect 15660 33992 15712 33998
rect 15660 33934 15712 33940
rect 15844 33992 15896 33998
rect 15844 33934 15896 33940
rect 12532 33924 12584 33930
rect 12532 33866 12584 33872
rect 12440 33652 12492 33658
rect 12440 33594 12492 33600
rect 12452 33522 12480 33594
rect 13176 33584 13228 33590
rect 13176 33526 13228 33532
rect 11152 33516 11204 33522
rect 11152 33458 11204 33464
rect 11336 33516 11388 33522
rect 11336 33458 11388 33464
rect 12440 33516 12492 33522
rect 12440 33458 12492 33464
rect 11060 33380 11112 33386
rect 11060 33322 11112 33328
rect 10692 33312 10744 33318
rect 10692 33254 10744 33260
rect 10968 33312 11020 33318
rect 10968 33254 11020 33260
rect 10232 32972 10284 32978
rect 10232 32914 10284 32920
rect 10704 32910 10732 33254
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 10140 32904 10192 32910
rect 10140 32846 10192 32852
rect 10692 32904 10744 32910
rect 10692 32846 10744 32852
rect 8944 32836 8996 32842
rect 8944 32778 8996 32784
rect 9968 32570 9996 32846
rect 11348 32842 11376 33458
rect 11428 33448 11480 33454
rect 11428 33390 11480 33396
rect 12348 33448 12400 33454
rect 12348 33390 12400 33396
rect 13084 33448 13136 33454
rect 13084 33390 13136 33396
rect 10600 32836 10652 32842
rect 10600 32778 10652 32784
rect 11336 32836 11388 32842
rect 11336 32778 11388 32784
rect 9956 32564 10008 32570
rect 9956 32506 10008 32512
rect 9864 32428 9916 32434
rect 9864 32370 9916 32376
rect 8668 32360 8720 32366
rect 8668 32302 8720 32308
rect 8300 31884 8352 31890
rect 8300 31826 8352 31832
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 8116 31408 8168 31414
rect 8116 31350 8168 31356
rect 8208 31408 8260 31414
rect 8208 31350 8260 31356
rect 7840 31272 7892 31278
rect 7840 31214 7892 31220
rect 7852 30938 7880 31214
rect 7840 30932 7892 30938
rect 7840 30874 7892 30880
rect 8220 30666 8248 31350
rect 8496 31210 8524 31622
rect 8680 31482 8708 32302
rect 9588 32224 9640 32230
rect 9588 32166 9640 32172
rect 9404 31748 9456 31754
rect 9404 31690 9456 31696
rect 9416 31482 9444 31690
rect 8668 31476 8720 31482
rect 8668 31418 8720 31424
rect 9128 31476 9180 31482
rect 9128 31418 9180 31424
rect 9404 31476 9456 31482
rect 9404 31418 9456 31424
rect 8760 31408 8812 31414
rect 8760 31350 8812 31356
rect 8484 31204 8536 31210
rect 8484 31146 8536 31152
rect 8496 30734 8524 31146
rect 8772 30938 8800 31350
rect 9140 31278 9168 31418
rect 9600 31414 9628 32166
rect 9588 31408 9640 31414
rect 9876 31362 9904 32370
rect 9968 31414 9996 32506
rect 10612 32434 10640 32778
rect 10600 32428 10652 32434
rect 10600 32370 10652 32376
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10416 31680 10468 31686
rect 10416 31622 10468 31628
rect 9588 31350 9640 31356
rect 9496 31340 9548 31346
rect 9496 31282 9548 31288
rect 9784 31334 9904 31362
rect 9956 31408 10008 31414
rect 9956 31350 10008 31356
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 8760 30932 8812 30938
rect 8760 30874 8812 30880
rect 8772 30734 8800 30874
rect 8484 30728 8536 30734
rect 8484 30670 8536 30676
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 8208 30660 8260 30666
rect 8208 30602 8260 30608
rect 7654 30288 7710 30297
rect 6828 30252 6880 30258
rect 7654 30223 7710 30232
rect 6828 30194 6880 30200
rect 6460 29708 6512 29714
rect 6460 29650 6512 29656
rect 6644 29708 6696 29714
rect 6644 29650 6696 29656
rect 6472 29306 6500 29650
rect 6460 29300 6512 29306
rect 6460 29242 6512 29248
rect 6276 29164 6328 29170
rect 6276 29106 6328 29112
rect 6288 28558 6316 29106
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 6276 28552 6328 28558
rect 6276 28494 6328 28500
rect 6564 28082 6592 29038
rect 6552 28076 6604 28082
rect 6552 28018 6604 28024
rect 6184 27872 6236 27878
rect 6184 27814 6236 27820
rect 6564 27418 6592 28018
rect 6656 27538 6684 29650
rect 6840 28762 6868 30194
rect 8220 29510 8248 30602
rect 8668 30592 8720 30598
rect 8668 30534 8720 30540
rect 8680 30326 8708 30534
rect 8668 30320 8720 30326
rect 8668 30262 8720 30268
rect 9036 30252 9088 30258
rect 9140 30240 9168 31214
rect 9508 31090 9536 31282
rect 9784 31210 9812 31334
rect 10428 31278 10456 31622
rect 10232 31272 10284 31278
rect 10232 31214 10284 31220
rect 10416 31272 10468 31278
rect 10416 31214 10468 31220
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9864 31204 9916 31210
rect 9864 31146 9916 31152
rect 10140 31204 10192 31210
rect 10140 31146 10192 31152
rect 9876 31090 9904 31146
rect 9508 31062 9904 31090
rect 9220 30660 9272 30666
rect 9220 30602 9272 30608
rect 9232 30394 9260 30602
rect 10152 30598 10180 31146
rect 10244 30938 10272 31214
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10140 30592 10192 30598
rect 10140 30534 10192 30540
rect 9220 30388 9272 30394
rect 9220 30330 9272 30336
rect 10244 30258 10272 30874
rect 9220 30252 9272 30258
rect 9140 30212 9220 30240
rect 9036 30194 9088 30200
rect 9220 30194 9272 30200
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 9048 29850 9076 30194
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 10244 29714 10272 30194
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 10428 29578 10456 31214
rect 10520 30666 10548 31758
rect 11440 31754 11468 33390
rect 11520 33312 11572 33318
rect 11520 33254 11572 33260
rect 11532 32910 11560 33254
rect 12360 33114 12388 33390
rect 12716 33380 12768 33386
rect 12716 33322 12768 33328
rect 12348 33108 12400 33114
rect 12348 33050 12400 33056
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 12164 32496 12216 32502
rect 12164 32438 12216 32444
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 11348 31726 11468 31754
rect 11532 31770 11560 31962
rect 12176 31822 12204 32438
rect 11612 31816 11664 31822
rect 11532 31764 11612 31770
rect 11532 31758 11664 31764
rect 12164 31816 12216 31822
rect 12164 31758 12216 31764
rect 11532 31742 11652 31758
rect 10876 31680 10928 31686
rect 10876 31622 10928 31628
rect 10968 31680 11020 31686
rect 10968 31622 11020 31628
rect 10888 31278 10916 31622
rect 10980 31346 11008 31622
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 10876 31272 10928 31278
rect 10876 31214 10928 31220
rect 10508 30660 10560 30666
rect 10508 30602 10560 30608
rect 10968 30660 11020 30666
rect 10968 30602 11020 30608
rect 10980 29782 11008 30602
rect 10968 29776 11020 29782
rect 10968 29718 11020 29724
rect 10416 29572 10468 29578
rect 10416 29514 10468 29520
rect 8208 29504 8260 29510
rect 8208 29446 8260 29452
rect 8220 29170 8248 29446
rect 8208 29164 8260 29170
rect 8208 29106 8260 29112
rect 10980 29102 11008 29718
rect 9496 29096 9548 29102
rect 9496 29038 9548 29044
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 10968 29096 11020 29102
rect 10968 29038 11020 29044
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 7472 28756 7524 28762
rect 7472 28698 7524 28704
rect 6644 27532 6696 27538
rect 6644 27474 6696 27480
rect 7484 27470 7512 28698
rect 9508 28626 9536 29038
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 7656 28552 7708 28558
rect 7656 28494 7708 28500
rect 7668 27878 7696 28494
rect 9508 28150 9536 28562
rect 9784 28218 9812 29038
rect 10876 28756 10928 28762
rect 10876 28698 10928 28704
rect 10888 28218 10916 28698
rect 10980 28490 11008 29038
rect 11244 29028 11296 29034
rect 11244 28970 11296 28976
rect 10968 28484 11020 28490
rect 10968 28426 11020 28432
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 10876 28212 10928 28218
rect 10876 28154 10928 28160
rect 9496 28144 9548 28150
rect 9496 28086 9548 28092
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 7656 27872 7708 27878
rect 7656 27814 7708 27820
rect 7104 27464 7156 27470
rect 6564 27390 6684 27418
rect 7104 27406 7156 27412
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 5998 26616 6054 26625
rect 5998 26551 6054 26560
rect 5814 26480 5870 26489
rect 5814 26415 5870 26424
rect 6012 26382 6040 26551
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 6000 26376 6052 26382
rect 6184 26376 6236 26382
rect 6000 26318 6052 26324
rect 6182 26344 6184 26353
rect 6236 26344 6238 26353
rect 5736 26042 5764 26318
rect 5724 26036 5776 26042
rect 5724 25978 5776 25984
rect 6012 25906 6040 26318
rect 6182 26279 6238 26288
rect 6092 26036 6144 26042
rect 6092 25978 6144 25984
rect 6104 25906 6132 25978
rect 5816 25900 5868 25906
rect 5816 25842 5868 25848
rect 6000 25900 6052 25906
rect 6000 25842 6052 25848
rect 6092 25900 6144 25906
rect 6092 25842 6144 25848
rect 5632 25764 5684 25770
rect 5632 25706 5684 25712
rect 5724 25696 5776 25702
rect 5724 25638 5776 25644
rect 5448 25424 5500 25430
rect 5448 25366 5500 25372
rect 5736 25158 5764 25638
rect 5828 25430 5856 25842
rect 5908 25764 5960 25770
rect 5908 25706 5960 25712
rect 5816 25424 5868 25430
rect 5816 25366 5868 25372
rect 5724 25152 5776 25158
rect 5724 25094 5776 25100
rect 5356 24880 5408 24886
rect 5356 24822 5408 24828
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 5092 24070 5120 24754
rect 5172 24200 5224 24206
rect 5224 24160 5580 24188
rect 5172 24142 5224 24148
rect 4712 24064 4764 24070
rect 4712 24006 4764 24012
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 5448 24064 5500 24070
rect 5448 24006 5500 24012
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4252 23656 4304 23662
rect 4252 23598 4304 23604
rect 1400 23316 1452 23322
rect 1400 23258 1452 23264
rect 1596 23225 1624 23462
rect 2700 23446 2820 23474
rect 1582 23216 1638 23225
rect 112 23180 164 23186
rect 1582 23151 1638 23160
rect 112 23122 164 23128
rect 2412 23044 2464 23050
rect 2412 22986 2464 22992
rect 2424 22710 2452 22986
rect 2412 22704 2464 22710
rect 2412 22646 2464 22652
rect 2792 22574 2820 23446
rect 2884 23050 2912 23582
rect 4160 23588 4212 23594
rect 4160 23530 4212 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5460 23322 5488 24006
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5552 23202 5580 24160
rect 5632 24132 5684 24138
rect 5632 24074 5684 24080
rect 5644 23322 5672 24074
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5552 23174 5672 23202
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 2872 23044 2924 23050
rect 2872 22986 2924 22992
rect 3252 22574 3280 23054
rect 5356 23044 5408 23050
rect 5408 23004 5488 23032
rect 5356 22986 5408 22992
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 2780 22568 2832 22574
rect 1306 22536 1362 22545
rect 2780 22510 2832 22516
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 1306 22471 1362 22480
rect 1320 21894 1348 22471
rect 1400 22432 1452 22438
rect 1400 22374 1452 22380
rect 1412 22030 1440 22374
rect 3252 22098 3280 22510
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1308 21888 1360 21894
rect 1308 21830 1360 21836
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2608 20942 2636 21286
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 1688 20466 1716 20878
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1688 19854 1716 20402
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1398 17776 1454 17785
rect 1596 17746 1624 18022
rect 1398 17711 1454 17720
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1688 17678 1716 19790
rect 1872 19514 1900 20402
rect 3068 20262 3096 20878
rect 3160 20602 3188 21422
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3056 20256 3108 20262
rect 3056 20198 3108 20204
rect 3252 19854 3280 22034
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4264 21622 4292 21966
rect 4724 21690 4752 22510
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4252 21616 4304 21622
rect 4252 21558 4304 21564
rect 4816 21554 4844 22374
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5276 21418 5304 21490
rect 5264 21412 5316 21418
rect 5264 21354 5316 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4620 21072 4672 21078
rect 4620 21014 4672 21020
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3344 20398 3372 20742
rect 3436 20466 3464 20742
rect 3424 20460 3476 20466
rect 3424 20402 3476 20408
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 3056 19780 3108 19786
rect 3056 19722 3108 19728
rect 3068 19514 3096 19722
rect 1860 19508 1912 19514
rect 1860 19450 1912 19456
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3252 19446 3280 19790
rect 3240 19440 3292 19446
rect 3240 19382 3292 19388
rect 3344 19310 3372 20334
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3712 19854 3740 20198
rect 3896 20058 3924 20334
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 3712 18766 3740 19790
rect 3700 18760 3752 18766
rect 3896 18748 3924 19994
rect 3988 18902 4016 20878
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 4528 20868 4580 20874
rect 4528 20810 4580 20816
rect 4172 20346 4200 20810
rect 4540 20602 4568 20810
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4632 20466 4660 21014
rect 5276 21010 5304 21354
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4080 20318 4200 20346
rect 4080 19938 4108 20318
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4724 20058 4752 20742
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4080 19910 4200 19938
rect 4172 19854 4200 19910
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4172 19446 4200 19790
rect 4344 19780 4396 19786
rect 4344 19722 4396 19728
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4356 19310 4384 19722
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4632 19310 4660 19654
rect 4724 19378 4752 19994
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4724 18970 4752 19314
rect 4816 19242 4844 20878
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5276 20466 5304 20946
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4896 19440 4948 19446
rect 4896 19382 4948 19388
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 3976 18896 4028 18902
rect 3976 18838 4028 18844
rect 4816 18766 4844 19178
rect 3976 18760 4028 18766
rect 3896 18720 3976 18748
rect 3700 18702 3752 18708
rect 3976 18702 4028 18708
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 18086 4844 18702
rect 4908 18630 4936 19382
rect 5276 19378 5304 20198
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 1676 17672 1728 17678
rect 1728 17620 1808 17626
rect 1676 17614 1808 17620
rect 1688 17598 1808 17614
rect 846 17232 902 17241
rect 846 17167 848 17176
rect 900 17167 902 17176
rect 848 17138 900 17144
rect 1780 17134 1808 17598
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16658 1624 16934
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1676 16584 1728 16590
rect 1780 16538 1808 17070
rect 1728 16532 1808 16538
rect 1676 16526 1808 16532
rect 1688 16510 1808 16526
rect 2792 16522 2820 17546
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 3068 17202 3096 17478
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3988 16522 4016 17138
rect 4632 16998 4660 17750
rect 5184 17678 5212 17750
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4724 17218 4752 17614
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4816 17338 4844 17546
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 5264 17332 5316 17338
rect 5368 17320 5396 20878
rect 5460 17898 5488 23004
rect 5644 22710 5672 23174
rect 5736 22778 5764 23666
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5540 22704 5592 22710
rect 5540 22646 5592 22652
rect 5632 22704 5684 22710
rect 5632 22646 5684 22652
rect 5552 22234 5580 22646
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5644 22094 5672 22646
rect 5552 22066 5672 22094
rect 5552 21554 5580 22066
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5828 21842 5856 23462
rect 5920 21962 5948 25706
rect 6368 25696 6420 25702
rect 6368 25638 6420 25644
rect 6092 25356 6144 25362
rect 6092 25298 6144 25304
rect 6104 24750 6132 25298
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 6092 24744 6144 24750
rect 6092 24686 6144 24692
rect 6104 24206 6132 24686
rect 6196 24274 6224 24754
rect 6184 24268 6236 24274
rect 6184 24210 6236 24216
rect 6092 24200 6144 24206
rect 6090 24168 6092 24177
rect 6144 24168 6146 24177
rect 6090 24103 6146 24112
rect 6000 23656 6052 23662
rect 6104 23644 6132 24103
rect 6052 23616 6132 23644
rect 6000 23598 6052 23604
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 6012 22001 6040 22918
rect 5998 21992 6054 22001
rect 5908 21956 5960 21962
rect 5998 21927 6054 21936
rect 5908 21898 5960 21904
rect 5736 21622 5764 21830
rect 5828 21814 5948 21842
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5644 21146 5672 21490
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5736 18970 5764 19246
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5460 17870 5672 17898
rect 5828 17882 5856 21626
rect 5920 19718 5948 21814
rect 6012 21350 6040 21927
rect 6196 21894 6224 24210
rect 6380 22030 6408 25638
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6472 24206 6500 25094
rect 6564 24410 6592 26930
rect 6656 26382 6684 27390
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6932 26382 6960 27270
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 6644 26376 6696 26382
rect 6644 26318 6696 26324
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 6552 24404 6604 24410
rect 6552 24346 6604 24352
rect 6460 24200 6512 24206
rect 6460 24142 6512 24148
rect 6472 23610 6500 24142
rect 6564 23730 6592 24346
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6472 23582 6592 23610
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 5920 19446 5948 19654
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5316 17292 5396 17320
rect 5264 17274 5316 17280
rect 4988 17264 5040 17270
rect 4894 17232 4950 17241
rect 4724 17190 4844 17218
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 860 15881 888 16050
rect 1780 16046 1808 16510
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2976 16114 3004 16390
rect 3988 16182 4016 16458
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1676 15904 1728 15910
rect 846 15872 902 15881
rect 1676 15846 1728 15852
rect 846 15807 902 15816
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12782 1440 13262
rect 1504 13025 1532 13670
rect 1596 13394 1624 15302
rect 1688 14414 1716 15846
rect 1780 15570 1808 15982
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 2240 14074 2268 15438
rect 3988 15434 4016 16118
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 3988 15094 4016 15370
rect 4632 15162 4660 16934
rect 4816 16590 4844 17190
rect 5460 17218 5488 17682
rect 5552 17241 5580 17682
rect 4988 17206 5040 17212
rect 4894 17167 4896 17176
rect 4948 17167 4950 17176
rect 4896 17138 4948 17144
rect 5000 16969 5028 17206
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5368 17190 5488 17218
rect 5538 17232 5594 17241
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 4986 16960 5042 16969
rect 4986 16895 5042 16904
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 15706 4844 16526
rect 4908 16522 4936 16662
rect 5184 16522 5212 17070
rect 5276 16658 5304 17138
rect 5368 17105 5396 17190
rect 5644 17218 5672 17870
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 6012 17814 6040 21286
rect 6196 20942 6224 21286
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6288 20602 6316 21422
rect 6380 20874 6408 21966
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6368 20868 6420 20874
rect 6368 20810 6420 20816
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 19310 6132 19858
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 5908 17808 5960 17814
rect 5908 17750 5960 17756
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5644 17190 5764 17218
rect 5538 17167 5594 17176
rect 5354 17096 5410 17105
rect 5354 17031 5410 17040
rect 5368 16658 5396 17031
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16658 5488 16934
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5368 16114 5396 16594
rect 5552 16182 5580 17167
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5644 16794 5672 17070
rect 5632 16788 5684 16794
rect 5632 16730 5684 16736
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 5368 15570 5396 15914
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 2700 14482 2728 14894
rect 3804 14618 3832 14894
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 3988 14346 4016 15030
rect 5184 14940 5212 15098
rect 5276 15094 5304 15438
rect 5552 15162 5580 16118
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 5184 14912 5396 14940
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4908 14618 4936 14758
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 2792 13258 2820 14282
rect 4632 14006 4660 14282
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4712 14000 4764 14006
rect 4712 13942 4764 13948
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 2976 13530 3004 13806
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 1490 13016 1546 13025
rect 1490 12951 1546 12960
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 12442 1808 12718
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 2688 12368 2740 12374
rect 1214 12336 1270 12345
rect 2688 12310 2740 12316
rect 1214 12271 1270 12280
rect 1228 10810 1256 12271
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1504 11218 1532 11630
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1780 10810 1808 11630
rect 1216 10804 1268 10810
rect 1216 10746 1268 10752
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 2700 10674 2728 12310
rect 2792 12170 2820 12582
rect 2884 12238 2912 12650
rect 3068 12646 3096 13806
rect 3344 13530 3372 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 4632 13002 4660 13942
rect 4724 13190 4752 13942
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 3804 12974 4660 13002
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11642 2820 12106
rect 3252 11762 3280 12854
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3436 12238 3464 12650
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 2792 11614 2912 11642
rect 2884 11218 2912 11614
rect 3252 11286 3280 11698
rect 3344 11665 3372 12038
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3330 11656 3386 11665
rect 3330 11591 3386 11600
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2792 10266 2820 10950
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 8906 1716 9318
rect 1676 8900 1728 8906
rect 1676 8842 1728 8848
rect 2516 8838 2544 9522
rect 2884 9024 2912 11154
rect 3252 11082 3280 11222
rect 3436 11150 3464 11562
rect 3528 11218 3556 11698
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3620 11150 3648 12174
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3620 10810 3648 11086
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3712 10742 3740 12582
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3160 10062 3188 10406
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3160 9042 3188 9522
rect 3436 9518 3464 9998
rect 3804 9738 3832 12974
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3988 11898 4016 12718
rect 4080 12238 4108 12786
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12238 4660 12786
rect 4724 12646 4752 13126
rect 4816 12986 4844 14010
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12238 5212 12582
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3988 10674 4016 11834
rect 4172 11830 4200 12174
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4540 11694 4568 12106
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 11354 4108 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11348 4120 11354
rect 4120 11308 4200 11336
rect 4068 11290 4120 11296
rect 4172 10674 4200 11308
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4264 10538 4292 10950
rect 4528 10668 4580 10674
rect 4632 10656 4660 12174
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4712 11892 4764 11898
rect 4816 11880 4844 12038
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4816 11852 4936 11880
rect 4712 11834 4764 11840
rect 4580 10628 4660 10656
rect 4528 10610 4580 10616
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 4724 10470 4752 11834
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4816 10810 4844 11698
rect 4908 11014 4936 11852
rect 5276 11762 5304 14758
rect 5368 14006 5396 14912
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5356 14000 5408 14006
rect 5356 13942 5408 13948
rect 5368 13462 5396 13942
rect 5460 13870 5488 14758
rect 5644 14074 5672 16390
rect 5736 15706 5764 17190
rect 5920 16998 5948 17750
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6012 17338 6040 17614
rect 6104 17542 6132 19246
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5920 16726 5948 16934
rect 6012 16794 6040 17138
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 6012 16114 6040 16730
rect 6104 16114 6132 17138
rect 6196 16658 6224 17614
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5736 15178 5764 15642
rect 5736 15150 5856 15178
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5736 14890 5764 15030
rect 5828 14958 5856 15150
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5632 14068 5684 14074
rect 5552 14028 5632 14056
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 13734 5488 13806
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5368 13190 5396 13398
rect 5460 13258 5488 13670
rect 5552 13394 5580 14028
rect 5632 14010 5684 14016
rect 5632 13932 5684 13938
rect 5736 13920 5764 14826
rect 5684 13892 5764 13920
rect 5632 13874 5684 13880
rect 5920 13870 5948 14962
rect 6012 14278 6040 16050
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6012 14006 6040 14214
rect 6104 14006 6132 16050
rect 6288 14822 6316 20334
rect 6472 20058 6500 21898
rect 6564 20466 6592 23582
rect 6656 22094 6684 26318
rect 7024 25752 7052 26386
rect 7116 26042 7144 27406
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 7104 25764 7156 25770
rect 7024 25724 7104 25752
rect 7104 25706 7156 25712
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6828 24676 6880 24682
rect 6828 24618 6880 24624
rect 6840 24206 6868 24618
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6840 23594 6868 24142
rect 6932 24070 6960 24754
rect 7116 24750 7144 25706
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 7024 24313 7052 24550
rect 7010 24304 7066 24313
rect 7116 24290 7144 24686
rect 7208 24614 7236 26318
rect 7668 25906 7696 27814
rect 8312 27606 8340 28018
rect 9036 27872 9088 27878
rect 9036 27814 9088 27820
rect 8300 27600 8352 27606
rect 8036 27538 8248 27554
rect 8300 27542 8352 27548
rect 9048 27538 9076 27814
rect 9692 27606 9720 28018
rect 10876 27872 10928 27878
rect 10876 27814 10928 27820
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 10888 27538 10916 27814
rect 10980 27674 11008 28426
rect 11256 28218 11284 28970
rect 11244 28212 11296 28218
rect 11244 28154 11296 28160
rect 11152 28076 11204 28082
rect 11072 28036 11152 28064
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 8024 27532 8248 27538
rect 8076 27526 8248 27532
rect 8024 27474 8076 27480
rect 8220 27452 8248 27526
rect 9036 27532 9088 27538
rect 9036 27474 9088 27480
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 8220 27424 8524 27452
rect 8116 27396 8168 27402
rect 8116 27338 8168 27344
rect 7932 27328 7984 27334
rect 7932 27270 7984 27276
rect 7944 26518 7972 27270
rect 7932 26512 7984 26518
rect 7932 26454 7984 26460
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 7300 24954 7328 25842
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 7392 24886 7420 25842
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7380 24880 7432 24886
rect 7380 24822 7432 24828
rect 7576 24750 7604 25230
rect 7472 24744 7524 24750
rect 7472 24686 7524 24692
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7288 24404 7340 24410
rect 7288 24346 7340 24352
rect 7116 24262 7236 24290
rect 7010 24239 7066 24248
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7116 24070 7144 24142
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 7208 23730 7236 24262
rect 7300 23798 7328 24346
rect 7380 24336 7432 24342
rect 7380 24278 7432 24284
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 6828 23588 6880 23594
rect 6828 23530 6880 23536
rect 6840 22438 6868 23530
rect 7208 23526 7236 23666
rect 7300 23610 7328 23734
rect 7392 23730 7420 24278
rect 7484 24206 7512 24686
rect 7576 24274 7604 24686
rect 7760 24682 7788 25230
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 7748 24676 7800 24682
rect 7748 24618 7800 24624
rect 7564 24268 7616 24274
rect 7564 24210 7616 24216
rect 7656 24268 7708 24274
rect 7656 24210 7708 24216
rect 7472 24200 7524 24206
rect 7668 24177 7696 24210
rect 7472 24142 7524 24148
rect 7654 24168 7710 24177
rect 7380 23724 7432 23730
rect 7380 23666 7432 23672
rect 7300 23582 7420 23610
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7288 23520 7340 23526
rect 7288 23462 7340 23468
rect 7208 23118 7236 23462
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 7116 22778 7144 23054
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 7104 22160 7156 22166
rect 7104 22102 7156 22108
rect 6656 22066 6776 22094
rect 6748 21570 6776 22066
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6840 21690 6868 21966
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6748 21542 6868 21570
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6656 21010 6684 21422
rect 6748 21146 6776 21422
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6656 19990 6684 20946
rect 6840 20262 6868 21542
rect 6932 20874 6960 21830
rect 6920 20868 6972 20874
rect 6920 20810 6972 20816
rect 7024 20806 7052 21830
rect 7116 21622 7144 22102
rect 7300 22030 7328 23462
rect 7392 23254 7420 23582
rect 7380 23248 7432 23254
rect 7380 23190 7432 23196
rect 7484 23118 7512 24142
rect 7852 24138 7880 25094
rect 7944 24954 7972 25842
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 7944 24290 7972 24550
rect 8036 24410 8064 25774
rect 8128 24954 8156 27338
rect 8496 26586 8524 27424
rect 9048 27062 9076 27474
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 9324 27130 9352 27270
rect 9312 27124 9364 27130
rect 9312 27066 9364 27072
rect 9036 27056 9088 27062
rect 9036 26998 9088 27004
rect 9416 26790 9444 27406
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 9496 26988 9548 26994
rect 9496 26930 9548 26936
rect 8668 26784 8720 26790
rect 8668 26726 8720 26732
rect 9404 26784 9456 26790
rect 9404 26726 9456 26732
rect 8484 26580 8536 26586
rect 8484 26522 8536 26528
rect 8496 26382 8524 26522
rect 8300 26376 8352 26382
rect 8300 26318 8352 26324
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 8312 26042 8340 26318
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 8680 25974 8708 26726
rect 9508 26586 9536 26930
rect 10152 26790 10180 27270
rect 10888 26994 10916 27474
rect 11072 27402 11100 28036
rect 11152 28018 11204 28024
rect 11060 27396 11112 27402
rect 11060 27338 11112 27344
rect 11152 27396 11204 27402
rect 11152 27338 11204 27344
rect 11164 27130 11192 27338
rect 11152 27124 11204 27130
rect 11152 27066 11204 27072
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10140 26784 10192 26790
rect 10140 26726 10192 26732
rect 9220 26580 9272 26586
rect 9220 26522 9272 26528
rect 9496 26580 9548 26586
rect 9496 26522 9548 26528
rect 9588 26580 9640 26586
rect 9588 26522 9640 26528
rect 9232 26466 9260 26522
rect 9600 26466 9628 26522
rect 9232 26438 9628 26466
rect 10152 26450 10180 26726
rect 10232 26512 10284 26518
rect 10232 26454 10284 26460
rect 10140 26444 10192 26450
rect 9232 26382 9260 26438
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 9220 26376 9272 26382
rect 9220 26318 9272 26324
rect 8956 26042 8984 26318
rect 8944 26036 8996 26042
rect 8944 25978 8996 25984
rect 8668 25968 8720 25974
rect 8668 25910 8720 25916
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8852 25900 8904 25906
rect 8852 25842 8904 25848
rect 8300 25220 8352 25226
rect 8300 25162 8352 25168
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 8312 24818 8340 25162
rect 8404 24954 8432 25842
rect 8588 25770 8616 25842
rect 8576 25764 8628 25770
rect 8576 25706 8628 25712
rect 8392 24948 8444 24954
rect 8392 24890 8444 24896
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8024 24404 8076 24410
rect 8024 24346 8076 24352
rect 8220 24342 8248 24754
rect 8864 24750 8892 25842
rect 9508 24970 9536 26438
rect 10140 26386 10192 26392
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9600 26042 9628 26318
rect 9588 26036 9640 26042
rect 9588 25978 9640 25984
rect 10244 25974 10272 26454
rect 10704 26450 10732 26930
rect 11348 26586 11376 31726
rect 11532 28558 11560 31742
rect 11612 31272 11664 31278
rect 11612 31214 11664 31220
rect 12624 31272 12676 31278
rect 12624 31214 12676 31220
rect 11624 30258 11652 31214
rect 12636 30938 12664 31214
rect 12624 30932 12676 30938
rect 12624 30874 12676 30880
rect 11612 30252 11664 30258
rect 11612 30194 11664 30200
rect 11624 29714 11652 30194
rect 11612 29708 11664 29714
rect 11612 29650 11664 29656
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11624 28490 11652 29650
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11808 29306 11836 29514
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 11980 28688 12032 28694
rect 11980 28630 12032 28636
rect 11612 28484 11664 28490
rect 11612 28426 11664 28432
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11532 28218 11560 28358
rect 11520 28212 11572 28218
rect 11520 28154 11572 28160
rect 11624 27878 11652 28426
rect 11992 28218 12020 28630
rect 12348 28484 12400 28490
rect 12348 28426 12400 28432
rect 11980 28212 12032 28218
rect 11980 28154 12032 28160
rect 12360 28014 12388 28426
rect 12544 28150 12572 29038
rect 12728 28694 12756 33322
rect 13096 33114 13124 33390
rect 13084 33108 13136 33114
rect 13084 33050 13136 33056
rect 13188 32298 13216 33526
rect 13636 33312 13688 33318
rect 13636 33254 13688 33260
rect 13176 32292 13228 32298
rect 13176 32234 13228 32240
rect 13188 31890 13216 32234
rect 13648 31890 13676 33254
rect 13820 32904 13872 32910
rect 13820 32846 13872 32852
rect 13176 31884 13228 31890
rect 13176 31826 13228 31832
rect 13636 31884 13688 31890
rect 13636 31826 13688 31832
rect 13832 31822 13860 32846
rect 13912 32836 13964 32842
rect 13912 32778 13964 32784
rect 13924 32434 13952 32778
rect 13912 32428 13964 32434
rect 13912 32370 13964 32376
rect 14464 32360 14516 32366
rect 14464 32302 14516 32308
rect 14476 32026 14504 32302
rect 14464 32020 14516 32026
rect 14464 31962 14516 31968
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 14464 31748 14516 31754
rect 14464 31690 14516 31696
rect 13452 31680 13504 31686
rect 13452 31622 13504 31628
rect 12900 31408 12952 31414
rect 12900 31350 12952 31356
rect 12912 30240 12940 31350
rect 13464 31346 13492 31622
rect 14476 31482 14504 31690
rect 14464 31476 14516 31482
rect 14464 31418 14516 31424
rect 13452 31340 13504 31346
rect 13452 31282 13504 31288
rect 12992 31204 13044 31210
rect 12992 31146 13044 31152
rect 13004 30734 13032 31146
rect 13360 30796 13412 30802
rect 13360 30738 13412 30744
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 13176 30592 13228 30598
rect 13176 30534 13228 30540
rect 12992 30252 13044 30258
rect 12912 30212 12992 30240
rect 12992 30194 13044 30200
rect 13004 29578 13032 30194
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 13096 29850 13124 30126
rect 13084 29844 13136 29850
rect 13084 29786 13136 29792
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 13188 28994 13216 30534
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 13280 29102 13308 29582
rect 13372 29306 13400 30738
rect 13464 30734 13492 31282
rect 13452 30728 13504 30734
rect 13452 30670 13504 30676
rect 13544 30728 13596 30734
rect 13544 30670 13596 30676
rect 13556 30258 13584 30670
rect 13544 30252 13596 30258
rect 13544 30194 13596 30200
rect 13912 30252 13964 30258
rect 13912 30194 13964 30200
rect 13556 29782 13584 30194
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 13544 29776 13596 29782
rect 13464 29736 13544 29764
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 13268 29096 13320 29102
rect 13268 29038 13320 29044
rect 13188 28966 13308 28994
rect 12900 28960 12952 28966
rect 12900 28902 12952 28908
rect 12992 28960 13044 28966
rect 12992 28902 13044 28908
rect 12716 28688 12768 28694
rect 12716 28630 12768 28636
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12532 28144 12584 28150
rect 12532 28086 12584 28092
rect 12636 28082 12664 28358
rect 12440 28076 12492 28082
rect 12440 28018 12492 28024
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 12348 28008 12400 28014
rect 12348 27950 12400 27956
rect 11612 27872 11664 27878
rect 11612 27814 11664 27820
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11992 27130 12020 27270
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 12084 26926 12112 27950
rect 12072 26920 12124 26926
rect 12072 26862 12124 26868
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 10692 26444 10744 26450
rect 10744 26404 10824 26432
rect 10692 26386 10744 26392
rect 10692 26240 10744 26246
rect 10692 26182 10744 26188
rect 10704 25974 10732 26182
rect 10232 25968 10284 25974
rect 10232 25910 10284 25916
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10796 25906 10824 26404
rect 11978 26344 12034 26353
rect 11978 26279 12034 26288
rect 11992 26246 12020 26279
rect 11520 26240 11572 26246
rect 11520 26182 11572 26188
rect 11980 26240 12032 26246
rect 11980 26182 12032 26188
rect 11532 26042 11560 26182
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 11992 25702 12020 26182
rect 12084 25922 12112 26862
rect 12164 26580 12216 26586
rect 12164 26522 12216 26528
rect 12176 26042 12204 26522
rect 12164 26036 12216 26042
rect 12164 25978 12216 25984
rect 12084 25894 12204 25922
rect 12452 25906 12480 28018
rect 12636 26858 12664 28018
rect 12728 27470 12756 28630
rect 12808 28552 12860 28558
rect 12912 28529 12940 28902
rect 12808 28494 12860 28500
rect 12898 28520 12954 28529
rect 12716 27464 12768 27470
rect 12716 27406 12768 27412
rect 12728 27062 12756 27406
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12820 25906 12848 28494
rect 12898 28455 12900 28464
rect 12952 28455 12954 28464
rect 12900 28426 12952 28432
rect 13004 26586 13032 28902
rect 12992 26580 13044 26586
rect 12992 26522 13044 26528
rect 13176 26444 13228 26450
rect 13176 26386 13228 26392
rect 13188 26314 13216 26386
rect 13176 26308 13228 26314
rect 13176 26250 13228 26256
rect 12176 25838 12204 25894
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12164 25832 12216 25838
rect 12164 25774 12216 25780
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 9140 24942 9628 24970
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8852 24744 8904 24750
rect 8852 24686 8904 24692
rect 8404 24410 8432 24686
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8208 24336 8260 24342
rect 7944 24262 8064 24290
rect 8208 24278 8260 24284
rect 8036 24138 8064 24262
rect 8220 24206 8248 24278
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 7654 24103 7710 24112
rect 7748 24132 7800 24138
rect 7748 24074 7800 24080
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 8024 24132 8076 24138
rect 8024 24074 8076 24080
rect 7564 24064 7616 24070
rect 7616 24012 7696 24018
rect 7564 24006 7696 24012
rect 7576 23990 7696 24006
rect 7668 23730 7696 23990
rect 7760 23866 7788 24074
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 7668 23118 7696 23666
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7472 23112 7524 23118
rect 7656 23112 7708 23118
rect 7524 23060 7604 23066
rect 7472 23054 7604 23060
rect 7656 23054 7708 23060
rect 7288 22024 7340 22030
rect 7392 22012 7420 23054
rect 7484 23038 7604 23054
rect 7472 22024 7524 22030
rect 7392 21992 7472 22012
rect 7524 21992 7526 22001
rect 7392 21984 7470 21992
rect 7288 21966 7340 21972
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7116 21026 7144 21558
rect 7300 21486 7328 21966
rect 7470 21927 7526 21936
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 7576 21350 7604 23038
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 22642 7788 22918
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7668 22234 7696 22510
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7760 22030 7788 22374
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7944 21894 7972 22714
rect 8036 22710 8064 24074
rect 8864 23746 8892 24686
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 8956 23866 8984 24142
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 8864 23718 8984 23746
rect 9048 23730 9076 24754
rect 9140 24138 9168 24942
rect 9600 24886 9628 24942
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9232 24313 9260 24754
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9218 24304 9274 24313
rect 9218 24239 9274 24248
rect 9232 24206 9260 24239
rect 9324 24206 9352 24346
rect 9508 24206 9536 24754
rect 10324 24744 10376 24750
rect 10324 24686 10376 24692
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 9588 24676 9640 24682
rect 9588 24618 9640 24624
rect 9600 24206 9628 24618
rect 10232 24608 10284 24614
rect 10232 24550 10284 24556
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 9312 24200 9364 24206
rect 9496 24200 9548 24206
rect 9312 24142 9364 24148
rect 9416 24160 9496 24188
rect 9128 24132 9180 24138
rect 9128 24074 9180 24080
rect 9416 24070 9444 24160
rect 9496 24142 9548 24148
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9416 23730 9444 24006
rect 9968 23730 9996 24142
rect 10244 23798 10272 24550
rect 10232 23792 10284 23798
rect 10232 23734 10284 23740
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 8864 21486 8892 21966
rect 8956 21486 8984 23718
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9876 22778 9904 23598
rect 10336 23526 10364 24686
rect 11348 24410 11376 24686
rect 11336 24404 11388 24410
rect 11336 24346 11388 24352
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10244 23118 10272 23462
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 10152 22710 10180 23054
rect 10140 22704 10192 22710
rect 10140 22646 10192 22652
rect 11152 22704 11204 22710
rect 11152 22646 11204 22652
rect 10152 22098 10180 22646
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 9036 21956 9088 21962
rect 9036 21898 9088 21904
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9048 21554 9076 21898
rect 9416 21690 9444 21898
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 8864 21146 8892 21422
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 7116 20998 7236 21026
rect 7012 20800 7064 20806
rect 7064 20748 7144 20754
rect 7012 20742 7144 20748
rect 7024 20726 7144 20742
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6380 18970 6408 19722
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6380 18154 6408 18906
rect 6368 18148 6420 18154
rect 6368 18090 6420 18096
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6380 16250 6408 17070
rect 6472 16969 6500 19654
rect 6656 19378 6684 19926
rect 6840 19922 6868 20198
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 19786 6868 19858
rect 7116 19786 7144 20726
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18970 6868 19110
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6932 18902 6960 19314
rect 7024 18902 7052 19654
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 7012 18896 7064 18902
rect 7012 18838 7064 18844
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6564 17202 6592 17546
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6748 17105 6776 17138
rect 6734 17096 6790 17105
rect 6734 17031 6790 17040
rect 6552 16992 6604 16998
rect 6458 16960 6514 16969
rect 6552 16934 6604 16940
rect 6458 16895 6514 16904
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6472 15706 6500 16895
rect 6564 16794 6592 16934
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6472 15450 6500 15642
rect 6472 15434 6684 15450
rect 6472 15428 6696 15434
rect 6472 15422 6644 15428
rect 6644 15370 6696 15376
rect 7116 15162 7144 19722
rect 7208 19718 7236 20998
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8404 20534 8432 20878
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8404 19990 8432 20470
rect 8956 20466 8984 21422
rect 10152 20942 10180 22034
rect 11164 21962 11192 22646
rect 11440 22642 11468 25162
rect 12072 24744 12124 24750
rect 12072 24686 12124 24692
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11808 23730 11836 24142
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 12084 22710 12112 24686
rect 12176 23186 12204 25774
rect 12452 23254 12480 25842
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12728 24857 12756 25638
rect 12714 24848 12770 24857
rect 12714 24783 12716 24792
rect 12768 24783 12770 24792
rect 12716 24754 12768 24760
rect 12820 24682 12848 25842
rect 13280 25276 13308 28966
rect 13372 27402 13400 29242
rect 13464 29170 13492 29736
rect 13544 29718 13596 29724
rect 13544 29504 13596 29510
rect 13544 29446 13596 29452
rect 13556 29170 13584 29446
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13544 29164 13596 29170
rect 13544 29106 13596 29112
rect 13556 29034 13584 29106
rect 13544 29028 13596 29034
rect 13544 28970 13596 28976
rect 13556 28762 13584 28970
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 13740 26314 13768 28154
rect 13728 26308 13780 26314
rect 13728 26250 13780 26256
rect 13452 25288 13504 25294
rect 13280 25256 13452 25276
rect 13504 25256 13506 25265
rect 13280 25248 13450 25256
rect 12808 24676 12860 24682
rect 12808 24618 12860 24624
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 12544 24206 12572 24550
rect 13004 24410 13032 24550
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 13096 23866 13124 24550
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 13004 23526 13032 23802
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12072 22704 12124 22710
rect 12072 22646 12124 22652
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 12452 22506 12480 23190
rect 13188 23118 13216 24550
rect 13280 23594 13308 25248
rect 13450 25191 13506 25200
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13648 24954 13676 25094
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 13648 23118 13676 24890
rect 13832 24818 13860 30126
rect 13924 29578 13952 30194
rect 14004 30048 14056 30054
rect 14004 29990 14056 29996
rect 14016 29714 14044 29990
rect 14004 29708 14056 29714
rect 14004 29650 14056 29656
rect 13912 29572 13964 29578
rect 13912 29514 13964 29520
rect 13924 28762 13952 29514
rect 13912 28756 13964 28762
rect 13912 28698 13964 28704
rect 14568 28558 14596 33934
rect 15672 33046 15700 33934
rect 15660 33040 15712 33046
rect 15660 32982 15712 32988
rect 15856 32978 15884 33934
rect 16592 33658 16620 37198
rect 16764 36780 16816 36786
rect 16764 36722 16816 36728
rect 16672 36576 16724 36582
rect 16672 36518 16724 36524
rect 16684 35222 16712 36518
rect 16776 36378 16804 36722
rect 16868 36718 16896 37878
rect 17144 37466 17172 38150
rect 17132 37460 17184 37466
rect 17132 37402 17184 37408
rect 17132 37256 17184 37262
rect 17132 37198 17184 37204
rect 16856 36712 16908 36718
rect 16856 36654 16908 36660
rect 17040 36712 17092 36718
rect 17040 36654 17092 36660
rect 16764 36372 16816 36378
rect 16764 36314 16816 36320
rect 16868 36258 16896 36654
rect 16868 36230 16988 36258
rect 16960 36174 16988 36230
rect 16948 36168 17000 36174
rect 16948 36110 17000 36116
rect 17052 35834 17080 36654
rect 17144 36174 17172 37198
rect 17236 36582 17264 39034
rect 17328 38418 17356 39918
rect 17420 39914 17448 40530
rect 17776 40384 17828 40390
rect 17776 40326 17828 40332
rect 17788 40118 17816 40326
rect 17776 40112 17828 40118
rect 17776 40054 17828 40060
rect 17408 39908 17460 39914
rect 17408 39850 17460 39856
rect 17420 38554 17448 39850
rect 17592 38752 17644 38758
rect 17592 38694 17644 38700
rect 17408 38548 17460 38554
rect 17408 38490 17460 38496
rect 17316 38412 17368 38418
rect 17316 38354 17368 38360
rect 17328 37942 17356 38354
rect 17420 37942 17448 38490
rect 17500 38344 17552 38350
rect 17500 38286 17552 38292
rect 17316 37936 17368 37942
rect 17316 37878 17368 37884
rect 17408 37936 17460 37942
rect 17408 37878 17460 37884
rect 17420 37466 17448 37878
rect 17408 37460 17460 37466
rect 17408 37402 17460 37408
rect 17224 36576 17276 36582
rect 17224 36518 17276 36524
rect 17132 36168 17184 36174
rect 17132 36110 17184 36116
rect 17040 35828 17092 35834
rect 17040 35770 17092 35776
rect 17144 35766 17172 36110
rect 17132 35760 17184 35766
rect 17132 35702 17184 35708
rect 17040 35624 17092 35630
rect 17040 35566 17092 35572
rect 16856 35556 16908 35562
rect 16856 35498 16908 35504
rect 16672 35216 16724 35222
rect 16672 35158 16724 35164
rect 16672 34944 16724 34950
rect 16672 34886 16724 34892
rect 16684 34066 16712 34886
rect 16672 34060 16724 34066
rect 16672 34002 16724 34008
rect 16580 33652 16632 33658
rect 16580 33594 16632 33600
rect 16764 33380 16816 33386
rect 16764 33322 16816 33328
rect 16776 32978 16804 33322
rect 15844 32972 15896 32978
rect 15844 32914 15896 32920
rect 16580 32972 16632 32978
rect 16580 32914 16632 32920
rect 16764 32972 16816 32978
rect 16764 32914 16816 32920
rect 15476 32836 15528 32842
rect 15476 32778 15528 32784
rect 15200 32768 15252 32774
rect 15200 32710 15252 32716
rect 15108 32224 15160 32230
rect 15212 32212 15240 32710
rect 15160 32184 15240 32212
rect 15108 32166 15160 32172
rect 15488 32026 15516 32778
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 15568 32428 15620 32434
rect 15568 32370 15620 32376
rect 15580 32026 15608 32370
rect 15476 32020 15528 32026
rect 15476 31962 15528 31968
rect 15568 32020 15620 32026
rect 15568 31962 15620 31968
rect 15384 31408 15436 31414
rect 15384 31350 15436 31356
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 14924 30320 14976 30326
rect 14924 30262 14976 30268
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 14648 28688 14700 28694
rect 14648 28630 14700 28636
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14464 28416 14516 28422
rect 14464 28358 14516 28364
rect 14476 28150 14504 28358
rect 14464 28144 14516 28150
rect 14464 28086 14516 28092
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 13912 27532 13964 27538
rect 14016 27520 14044 27814
rect 14476 27606 14504 27950
rect 14464 27600 14516 27606
rect 14464 27542 14516 27548
rect 13964 27492 14044 27520
rect 13912 27474 13964 27480
rect 13924 26450 13952 27474
rect 14370 27432 14426 27441
rect 14370 27367 14426 27376
rect 14384 27334 14412 27367
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14464 27328 14516 27334
rect 14464 27270 14516 27276
rect 13912 26444 13964 26450
rect 13912 26386 13964 26392
rect 14476 26217 14504 27270
rect 14568 27062 14596 28494
rect 14660 27470 14688 28630
rect 14752 28218 14780 29446
rect 14936 28626 14964 30262
rect 15212 29646 15240 30534
rect 15396 30054 15424 31350
rect 15488 31346 15516 31962
rect 16040 31822 16068 32710
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 16120 32224 16172 32230
rect 16120 32166 16172 32172
rect 16132 31822 16160 32166
rect 16408 32026 16436 32370
rect 16396 32020 16448 32026
rect 16396 31962 16448 31968
rect 16408 31890 16436 31962
rect 16396 31884 16448 31890
rect 16396 31826 16448 31832
rect 16028 31816 16080 31822
rect 16028 31758 16080 31764
rect 16120 31816 16172 31822
rect 16120 31758 16172 31764
rect 16592 31754 16620 32914
rect 16868 32502 16896 35498
rect 17052 34066 17080 35566
rect 17144 35154 17172 35702
rect 17316 35488 17368 35494
rect 17316 35430 17368 35436
rect 17328 35290 17356 35430
rect 17316 35284 17368 35290
rect 17316 35226 17368 35232
rect 17132 35148 17184 35154
rect 17132 35090 17184 35096
rect 17144 34542 17172 35090
rect 17224 35012 17276 35018
rect 17224 34954 17276 34960
rect 17236 34746 17264 34954
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 17132 34536 17184 34542
rect 17132 34478 17184 34484
rect 17512 34134 17540 38286
rect 17604 38282 17632 38694
rect 17592 38276 17644 38282
rect 17592 38218 17644 38224
rect 17684 38208 17736 38214
rect 17684 38150 17736 38156
rect 17696 38010 17724 38150
rect 17684 38004 17736 38010
rect 17684 37946 17736 37952
rect 17592 37664 17644 37670
rect 17592 37606 17644 37612
rect 17604 37330 17632 37606
rect 17592 37324 17644 37330
rect 17592 37266 17644 37272
rect 17592 35692 17644 35698
rect 17592 35634 17644 35640
rect 17500 34128 17552 34134
rect 17500 34070 17552 34076
rect 17040 34060 17092 34066
rect 17040 34002 17092 34008
rect 17052 33046 17080 34002
rect 17316 33856 17368 33862
rect 17316 33798 17368 33804
rect 17224 33516 17276 33522
rect 17224 33458 17276 33464
rect 17236 33114 17264 33458
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17040 33040 17092 33046
rect 17040 32982 17092 32988
rect 16856 32496 16908 32502
rect 16854 32464 16856 32473
rect 16908 32464 16910 32473
rect 16854 32399 16910 32408
rect 16580 31748 16632 31754
rect 16580 31690 16632 31696
rect 16672 31748 16724 31754
rect 16672 31690 16724 31696
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 15948 31482 15976 31622
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 16488 31476 16540 31482
rect 16488 31418 16540 31424
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 16500 30394 16528 31418
rect 16592 31278 16620 31690
rect 16580 31272 16632 31278
rect 16580 31214 16632 31220
rect 16580 31136 16632 31142
rect 16580 31078 16632 31084
rect 16488 30388 16540 30394
rect 16488 30330 16540 30336
rect 16304 30184 16356 30190
rect 16304 30126 16356 30132
rect 15384 30048 15436 30054
rect 15384 29990 15436 29996
rect 16316 29850 16344 30126
rect 16304 29844 16356 29850
rect 16304 29786 16356 29792
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 16212 29504 16264 29510
rect 16212 29446 16264 29452
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 15568 28620 15620 28626
rect 15568 28562 15620 28568
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14740 28212 14792 28218
rect 14740 28154 14792 28160
rect 14844 27878 14872 28358
rect 14832 27872 14884 27878
rect 14832 27814 14884 27820
rect 14936 27538 14964 28562
rect 15200 28484 15252 28490
rect 15200 28426 15252 28432
rect 15212 28218 15240 28426
rect 15200 28212 15252 28218
rect 15200 28154 15252 28160
rect 15016 28076 15068 28082
rect 15016 28018 15068 28024
rect 14924 27532 14976 27538
rect 14924 27474 14976 27480
rect 15028 27470 15056 28018
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 15120 27878 15148 27950
rect 15108 27872 15160 27878
rect 15108 27814 15160 27820
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 15016 27464 15068 27470
rect 15016 27406 15068 27412
rect 14832 27396 14884 27402
rect 14832 27338 14884 27344
rect 14924 27396 14976 27402
rect 14924 27338 14976 27344
rect 14556 27056 14608 27062
rect 14556 26998 14608 27004
rect 14844 26790 14872 27338
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 14936 26586 14964 27338
rect 15028 27130 15056 27406
rect 15120 27334 15148 27814
rect 15396 27690 15424 27814
rect 15212 27662 15424 27690
rect 15212 27606 15240 27662
rect 15200 27600 15252 27606
rect 15200 27542 15252 27548
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15108 27328 15160 27334
rect 15108 27270 15160 27276
rect 15016 27124 15068 27130
rect 15016 27066 15068 27072
rect 15014 27024 15070 27033
rect 15014 26959 15070 26968
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 14924 26444 14976 26450
rect 14924 26386 14976 26392
rect 14556 26240 14608 26246
rect 14462 26208 14518 26217
rect 14556 26182 14608 26188
rect 14462 26143 14518 26152
rect 14372 25900 14424 25906
rect 14372 25842 14424 25848
rect 14384 25226 14412 25842
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 14372 24812 14424 24818
rect 14476 24800 14504 26143
rect 14568 25906 14596 26182
rect 14738 26072 14794 26081
rect 14936 26042 14964 26386
rect 14738 26007 14740 26016
rect 14792 26007 14794 26016
rect 14924 26036 14976 26042
rect 14740 25978 14792 25984
rect 14924 25978 14976 25984
rect 15028 25906 15056 26959
rect 15304 26790 15332 27542
rect 15396 26926 15424 27662
rect 15580 27402 15608 28562
rect 16118 27568 16174 27577
rect 16118 27503 16174 27512
rect 15568 27396 15620 27402
rect 15568 27338 15620 27344
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15384 26920 15436 26926
rect 15384 26862 15436 26868
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15304 25906 15332 26726
rect 15474 26480 15530 26489
rect 15474 26415 15476 26424
rect 15528 26415 15530 26424
rect 15476 26386 15528 26392
rect 15580 25974 15608 27338
rect 15672 27130 15700 27338
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 15752 26852 15804 26858
rect 15752 26794 15804 26800
rect 15764 26382 15792 26794
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15856 26382 15884 26726
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15844 26376 15896 26382
rect 15844 26318 15896 26324
rect 15948 26364 15976 26998
rect 16028 26376 16080 26382
rect 15948 26336 16028 26364
rect 15568 25968 15620 25974
rect 15568 25910 15620 25916
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15476 25900 15528 25906
rect 15476 25842 15528 25848
rect 14568 25226 14596 25842
rect 14844 25702 14872 25842
rect 14924 25832 14976 25838
rect 14924 25774 14976 25780
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14936 25650 14964 25774
rect 15108 25764 15160 25770
rect 15108 25706 15160 25712
rect 14844 25498 14872 25638
rect 14936 25622 15056 25650
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 14936 25242 14964 25434
rect 15028 25294 15056 25622
rect 15120 25362 15148 25706
rect 15488 25702 15516 25842
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15580 25378 15608 25910
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 15488 25350 15608 25378
rect 14556 25220 14608 25226
rect 14556 25162 14608 25168
rect 14844 25214 14964 25242
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 14424 24772 14504 24800
rect 14372 24754 14424 24760
rect 13832 23526 13860 24754
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14016 24342 14044 24550
rect 14004 24336 14056 24342
rect 14004 24278 14056 24284
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14108 24154 14136 24210
rect 14016 24126 14136 24154
rect 14016 23662 14044 24126
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 14004 23656 14056 23662
rect 14004 23598 14056 23604
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13924 23186 13952 23598
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13636 23112 13688 23118
rect 13636 23054 13688 23060
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12636 22778 12664 22918
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12440 22500 12492 22506
rect 12440 22442 12492 22448
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11164 21622 11192 21898
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11624 21554 11652 21966
rect 12268 21622 12296 22374
rect 12820 22030 12848 22374
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 13004 21690 13032 23054
rect 13728 23044 13780 23050
rect 13728 22986 13780 22992
rect 13740 22710 13768 22986
rect 13728 22704 13780 22710
rect 13728 22646 13780 22652
rect 14016 22574 14044 23598
rect 14200 23186 14228 24550
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14188 22976 14240 22982
rect 14188 22918 14240 22924
rect 14200 22710 14228 22918
rect 14188 22704 14240 22710
rect 14188 22646 14240 22652
rect 14292 22642 14320 23734
rect 14568 23186 14596 25162
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14752 24410 14780 24754
rect 14740 24404 14792 24410
rect 14740 24346 14792 24352
rect 14844 24206 14872 25214
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14936 24818 14964 25094
rect 15028 24886 15056 25230
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 14924 24812 14976 24818
rect 14924 24754 14976 24760
rect 15488 24682 15516 25350
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15476 24676 15528 24682
rect 15476 24618 15528 24624
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14844 23118 14872 24142
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 14476 22778 14504 23054
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 14476 22234 14504 22714
rect 15120 22234 15148 23054
rect 15304 22778 15332 23054
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 15396 22094 15424 24550
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15488 22098 15516 23190
rect 15580 23118 15608 25230
rect 15672 24818 15700 26318
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15764 26081 15792 26182
rect 15750 26072 15806 26081
rect 15750 26007 15806 26016
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15856 25362 15884 25638
rect 15844 25356 15896 25362
rect 15844 25298 15896 25304
rect 15948 24818 15976 26336
rect 16028 26318 16080 26324
rect 16132 26314 16160 27503
rect 16120 26308 16172 26314
rect 16120 26250 16172 26256
rect 16028 25832 16080 25838
rect 16132 25820 16160 26250
rect 16080 25792 16160 25820
rect 16028 25774 16080 25780
rect 16132 24954 16160 25792
rect 16120 24948 16172 24954
rect 16120 24890 16172 24896
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 15672 24682 15700 24754
rect 15660 24676 15712 24682
rect 15660 24618 15712 24624
rect 15948 24614 15976 24754
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15580 22574 15608 23054
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15304 22066 15424 22094
rect 15476 22092 15528 22098
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 15028 21554 15056 21830
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9784 20602 9812 20810
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8496 19854 8524 20334
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 9140 19802 9168 20402
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9772 19848 9824 19854
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 19446 7236 19654
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 8128 19378 8156 19790
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7392 17202 7420 18022
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7484 17338 7512 17546
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7668 17134 7696 17614
rect 7656 17128 7708 17134
rect 7576 17088 7656 17116
rect 7576 15502 7604 17088
rect 7656 17070 7708 17076
rect 7760 15978 7788 18634
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 7944 17202 7972 18566
rect 8128 18154 8156 19110
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 8128 16794 8156 17138
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 8220 15706 8248 16118
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8220 15502 8248 15642
rect 7564 15496 7616 15502
rect 8208 15496 8260 15502
rect 7564 15438 7616 15444
rect 8128 15456 8208 15484
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 11898 5396 13126
rect 5460 12850 5488 13194
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5460 12306 5488 12786
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5644 12442 5672 12718
rect 5736 12442 5764 13330
rect 5828 13326 5856 13670
rect 5816 13320 5868 13326
rect 6012 13308 6040 13942
rect 6564 13530 6592 13942
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 5816 13262 5868 13268
rect 5920 13280 6040 13308
rect 6736 13320 6788 13326
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5736 12306 5764 12378
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5920 12238 5948 13280
rect 6736 13262 6788 13268
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6012 12986 6040 13126
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6472 12646 6500 13126
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 5908 12232 5960 12238
rect 5906 12200 5908 12209
rect 5960 12200 5962 12209
rect 5906 12135 5962 12144
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5828 11830 5856 12038
rect 6564 11898 6592 12718
rect 6748 12306 6776 13262
rect 6840 12850 6868 14962
rect 7576 14958 7604 15438
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 7944 15162 7972 15370
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 8128 14958 8156 15456
rect 8208 15438 8260 15444
rect 8312 15094 8340 19450
rect 8680 19446 8708 19790
rect 9140 19786 9352 19802
rect 9772 19790 9824 19796
rect 9140 19780 9364 19786
rect 9140 19774 9312 19780
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8864 19446 8892 19654
rect 9140 19514 9168 19774
rect 9312 19722 9364 19728
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 8668 19440 8720 19446
rect 8668 19382 8720 19388
rect 8852 19440 8904 19446
rect 8852 19382 8904 19388
rect 9692 19378 9720 19654
rect 9784 19378 9812 19790
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8404 18426 8432 18702
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8496 18290 8524 18770
rect 9232 18766 9260 19246
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8496 16590 8524 18226
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8496 16250 8524 16526
rect 8680 16522 8708 18634
rect 9416 18630 9444 19246
rect 9692 18902 9720 19314
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9692 18290 9720 18838
rect 9968 18698 9996 19110
rect 10060 18850 10088 19994
rect 10508 19984 10560 19990
rect 10508 19926 10560 19932
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10152 18970 10180 19790
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10428 19446 10456 19654
rect 10520 19514 10548 19926
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10416 19440 10468 19446
rect 10416 19382 10468 19388
rect 10796 18970 10824 20946
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 20466 11008 20742
rect 11624 20466 11652 21490
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11624 19990 11652 20402
rect 11808 20058 11836 20946
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12268 20534 12296 20742
rect 13188 20602 13216 20878
rect 14384 20874 14412 21286
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 13176 20596 13228 20602
rect 13096 20556 13176 20584
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11612 19984 11664 19990
rect 11612 19926 11664 19932
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10060 18822 10180 18850
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9876 18358 9904 18566
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 10060 18290 10088 18702
rect 10152 18426 10180 18822
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 8864 17542 8892 18158
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 9232 16998 9260 18226
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17610 9812 18022
rect 10152 17678 10180 18362
rect 10244 17746 10272 18566
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10520 17678 10548 18770
rect 10796 18698 10824 18906
rect 10888 18766 10916 19450
rect 10980 19446 11008 19790
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 11532 19310 11560 19790
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 11348 18698 11376 19246
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11624 18426 11652 19790
rect 11808 19378 11836 19994
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 12084 19310 12112 19654
rect 12268 19514 12296 19722
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12084 18850 12112 19246
rect 12268 18970 12296 19314
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 11808 18822 12112 18850
rect 12544 18834 12572 19246
rect 12532 18828 12584 18834
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9416 17202 9444 17478
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9416 16590 9444 16934
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 8864 16250 8892 16458
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 9140 15638 9168 16526
rect 9416 15910 9444 16526
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9036 15632 9088 15638
rect 9036 15574 9088 15580
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8496 15026 8524 15302
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 7576 14482 7604 14894
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8312 13938 8340 14418
rect 9048 14414 9076 15574
rect 9588 15496 9640 15502
rect 9692 15484 9720 16458
rect 9640 15456 9720 15484
rect 9588 15438 9640 15444
rect 9876 14464 9904 17478
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9968 16658 9996 17138
rect 10520 16998 10548 17614
rect 10612 17338 10640 18226
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9968 16182 9996 16594
rect 10336 16522 10364 16934
rect 10888 16794 10916 17818
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11072 16726 11100 17070
rect 11440 16794 11468 17138
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9968 15570 9996 16118
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15042 9996 15506
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10060 15162 10088 15438
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9968 15014 10088 15042
rect 10060 14822 10088 15014
rect 10336 14958 10364 16458
rect 11072 16046 11100 16662
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11704 15972 11756 15978
rect 11808 15960 11836 18822
rect 12532 18770 12584 18776
rect 12072 18760 12124 18766
rect 12716 18760 12768 18766
rect 12072 18702 12124 18708
rect 12544 18708 12716 18714
rect 12544 18702 12768 18708
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 16046 11928 16390
rect 11992 16182 12020 16458
rect 12084 16250 12112 18702
rect 12544 18698 12756 18702
rect 12532 18692 12756 18698
rect 12584 18686 12756 18692
rect 12532 18634 12584 18640
rect 12544 18358 12572 18634
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12820 18222 12848 18702
rect 13096 18698 13124 20556
rect 13176 20538 13228 20544
rect 14476 20398 14504 20810
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14476 19854 14504 20334
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13188 19242 13216 19654
rect 13832 19378 13860 19790
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13176 19236 13228 19242
rect 13176 19178 13228 19184
rect 13188 18698 13216 19178
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13188 18290 13216 18634
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12544 17746 12572 18158
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 17746 12848 18022
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12360 17270 12388 17546
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12360 16794 12388 17206
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12452 16522 12480 17274
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 12544 16130 12572 17070
rect 12636 16522 12664 17138
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12728 16436 12756 17478
rect 12820 17338 12848 17682
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12820 16794 12848 17070
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16794 12940 16934
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13004 16522 13032 17002
rect 13280 16794 13308 17138
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 12808 16448 12860 16454
rect 12728 16408 12808 16436
rect 12624 16176 12676 16182
rect 12544 16124 12624 16130
rect 12544 16118 12676 16124
rect 11992 16046 12020 16118
rect 12544 16102 12664 16118
rect 12728 16114 12756 16408
rect 12808 16390 12860 16396
rect 12912 16250 12940 16458
rect 12900 16244 12952 16250
rect 13464 16232 13492 19246
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13556 16590 13584 17478
rect 13648 16658 13676 18702
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14200 18358 14228 18566
rect 14188 18352 14240 18358
rect 14188 18294 14240 18300
rect 14384 18290 14412 19314
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13924 16794 13952 17546
rect 14384 17134 14412 18226
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13636 16244 13688 16250
rect 13464 16204 13636 16232
rect 12900 16186 12952 16192
rect 13636 16186 13688 16192
rect 12716 16108 12768 16114
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11980 16040 12032 16046
rect 12544 15994 12572 16102
rect 12716 16050 12768 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 11980 15982 12032 15988
rect 11756 15932 11836 15960
rect 11704 15914 11756 15920
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 10704 15638 10732 15846
rect 11624 15706 11652 15846
rect 11808 15706 11836 15932
rect 11992 15706 12020 15982
rect 12452 15978 12572 15994
rect 12440 15972 12572 15978
rect 12492 15966 12572 15972
rect 12440 15914 12492 15920
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10336 14618 10364 14894
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 9876 14436 9996 14464
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9876 14006 9904 14282
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 8312 13394 8340 13874
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8772 13326 8800 13738
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8036 12986 8064 13194
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6840 12714 6868 12786
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 8576 12708 8628 12714
rect 8576 12650 8628 12656
rect 6736 12300 6788 12306
rect 6788 12260 6868 12288
rect 6736 12242 6788 12248
rect 6642 12200 6698 12209
rect 6642 12135 6644 12144
rect 6696 12135 6698 12144
rect 6644 12106 6696 12112
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11914 6776 12038
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6656 11886 6776 11914
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5460 11014 5488 11766
rect 5920 11762 5948 11834
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 6552 11756 6604 11762
rect 6656 11744 6684 11886
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6604 11716 6684 11744
rect 6552 11698 6604 11704
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 5460 10606 5488 10950
rect 5644 10674 5672 11494
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10062 4660 10406
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 3712 9710 3832 9738
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3436 9382 3464 9454
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 2964 9036 3016 9042
rect 2884 8996 2964 9024
rect 2964 8978 3016 8984
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 1964 8430 1992 8774
rect 2976 8498 3004 8978
rect 3436 8974 3464 9318
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3712 8906 3740 9710
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8566 3372 8774
rect 3712 8566 3740 8842
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3700 8560 3752 8566
rect 3700 8502 3752 8508
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 6458 1440 7822
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1780 7546 1808 7754
rect 1964 7750 1992 8366
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1964 7410 1992 7686
rect 2240 7478 2268 8230
rect 2884 8090 2912 8366
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3712 7886 3740 8502
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 2884 6798 2912 7482
rect 2976 7002 3004 7822
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7546 3280 7686
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1412 6322 1440 6394
rect 1688 6390 1716 6598
rect 2976 6390 3004 6938
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 3068 6798 3096 6870
rect 3252 6798 3280 7482
rect 3620 7410 3648 7754
rect 3804 7750 3832 9046
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3896 8090 3924 8842
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3896 7886 3924 8026
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3988 7750 4016 9114
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8090 4660 9454
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4724 8294 4752 8910
rect 4816 8430 4844 10542
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5276 9586 5304 10406
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5368 8974 5396 9862
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5460 8922 5488 9998
rect 5552 9042 5580 10474
rect 5828 10062 5856 10610
rect 5920 10062 5948 10950
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6012 10266 6040 10542
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5736 9722 5764 9930
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 5368 8294 5396 8910
rect 5460 8894 5580 8922
rect 5552 8838 5580 8894
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4724 7886 4752 8230
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3804 6934 3832 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3252 6390 3280 6734
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 5778 1440 6258
rect 2976 5794 3004 6326
rect 1400 5772 1452 5778
rect 2976 5766 3096 5794
rect 1400 5714 1452 5720
rect 3068 5710 3096 5766
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3252 5370 3280 5714
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3344 5234 3372 6598
rect 3804 6390 3832 6870
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3436 5778 3464 6054
rect 3528 5914 3556 6054
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3896 5846 3924 6258
rect 3988 6118 4016 6734
rect 4448 6390 4476 6938
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 6458 4660 6734
rect 5552 6662 5580 6938
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4080 6118 4108 6258
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3436 5302 3464 5714
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 4080 5166 4108 5850
rect 4632 5778 4660 6394
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4724 5914 4752 6326
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4356 5302 4384 5714
rect 4724 5302 4752 5850
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4816 4826 4844 5646
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5552 5370 5580 5510
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5644 4826 5672 9522
rect 5736 8566 5764 9522
rect 5920 9466 5948 9998
rect 5828 9438 5948 9466
rect 6012 9450 6040 10202
rect 6564 10198 6592 11698
rect 6748 11150 6776 11766
rect 6840 11762 6868 12260
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 7024 11694 7052 12174
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 7116 10742 7144 12038
rect 7484 11898 7512 12174
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7116 10606 7144 10678
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7300 10554 7328 11630
rect 7392 11286 7420 11766
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7392 10674 7420 11222
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7300 10526 7420 10554
rect 7392 10470 7420 10526
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 7300 10062 7328 10406
rect 7392 10266 7420 10406
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7484 10146 7512 11494
rect 8312 10810 8340 11834
rect 8404 10810 8432 11834
rect 8588 11830 8616 12650
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8772 11762 8800 13262
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 12102 8892 12786
rect 9416 12306 9444 13874
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12986 9628 13126
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9968 12850 9996 14436
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10336 13258 10364 13942
rect 10704 13530 10732 14350
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 14074 11744 14214
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11808 13938 11836 15642
rect 12820 15502 12848 15846
rect 13004 15502 13032 15846
rect 13280 15502 13308 16050
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13372 15502 13400 15914
rect 13648 15502 13676 16186
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13832 15706 13860 16050
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 15026 12664 15302
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 13004 14958 13032 15438
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13556 15162 13584 15370
rect 14384 15366 14412 17070
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15212 15978 15240 16526
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 15212 15502 15240 15914
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 15212 15026 15240 15438
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 14074 12020 14350
rect 12176 14074 12204 14418
rect 12360 14074 12388 14826
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10324 13252 10376 13258
rect 10324 13194 10376 13200
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12306 9720 12582
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8864 11762 8892 12038
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8208 10668 8260 10674
rect 7944 10628 8208 10656
rect 7944 10538 7972 10628
rect 8208 10610 8260 10616
rect 8496 10538 8524 11086
rect 8680 10810 8708 11086
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 7392 10118 7512 10146
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 6000 9444 6052 9450
rect 5828 8974 5856 9438
rect 6000 9386 6052 9392
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9042 5948 9318
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 6104 8906 6132 9998
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6196 9178 6224 9590
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 6104 8498 6132 8842
rect 6288 8634 6316 9386
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 9042 6408 9318
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6472 8498 6500 9862
rect 6564 9178 6592 9998
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 8838 6592 8910
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6564 8294 6592 8774
rect 6656 8634 6684 9862
rect 6748 8906 6776 9998
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6840 9382 6868 9658
rect 7392 9654 7420 10118
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6840 9042 6868 9318
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6932 8974 6960 9522
rect 7392 9466 7420 9590
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 7300 9450 7420 9466
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7288 9444 7420 9450
rect 7340 9438 7420 9444
rect 7288 9386 7340 9392
rect 7484 9178 7512 9454
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 7484 8498 7512 9114
rect 8036 9042 8064 9318
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6012 6934 6040 8230
rect 8312 8090 8340 9522
rect 8496 9518 8524 10474
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8404 8974 8432 9386
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8404 8430 8432 8910
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8404 7818 8432 8366
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5724 6792 5776 6798
rect 5776 6740 5856 6746
rect 5724 6734 5856 6740
rect 5736 6718 5856 6734
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 5710 5764 6598
rect 5828 6118 5856 6718
rect 5920 6254 5948 6802
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5828 4622 5856 6054
rect 5920 5166 5948 6190
rect 6012 5370 6040 6666
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6012 4758 6040 5306
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 6104 4554 6132 6938
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6380 6390 6408 6598
rect 6564 6390 6592 6802
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7116 6474 7144 6734
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7024 6446 7144 6474
rect 7024 6390 7052 6446
rect 7392 6390 7420 6598
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6196 5166 6224 5578
rect 6380 5166 6408 6326
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 5778 6868 6190
rect 7484 6118 7512 6734
rect 8404 6458 8432 6802
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8496 6390 8524 8502
rect 8588 7818 8616 9862
rect 8772 8634 8800 11698
rect 8956 11642 8984 12038
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9508 11694 9536 11766
rect 8864 11614 8984 11642
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 8864 11218 8892 11614
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8956 11354 8984 11494
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 9048 11014 9076 11494
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9324 11082 9352 11290
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10674 9076 10950
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9692 10588 9720 11630
rect 9772 10600 9824 10606
rect 9692 10560 9772 10588
rect 9772 10542 9824 10548
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 9048 8566 9076 8774
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 9324 8498 9352 8978
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8772 7002 8800 7890
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8588 6118 8616 6938
rect 9048 6866 9076 7686
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6840 5234 6868 5714
rect 8864 5710 8892 6394
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 5914 8984 6190
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9140 5710 9168 6734
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9324 6338 9352 6666
rect 9416 6662 9444 8910
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9508 8498 9536 8570
rect 9876 8498 9904 12650
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10060 10470 10088 11834
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10152 9586 10180 11494
rect 10336 11150 10364 13194
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10336 10742 10364 11086
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10060 8566 10088 8842
rect 10152 8634 10180 9318
rect 10244 9178 10272 9318
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10336 8906 10364 10678
rect 10428 9586 10456 12922
rect 10704 12850 10732 13466
rect 11348 13326 11376 13670
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 11164 12646 11192 13262
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 12238 11192 12582
rect 11256 12442 11284 12786
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11348 12306 11376 13262
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11440 12714 11468 13126
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11440 12442 11468 12650
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11286 10732 11630
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10336 8650 10364 8842
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10244 8622 10364 8650
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9692 8090 9720 8434
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9968 8022 9996 8366
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 10152 7886 10180 8434
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10244 6746 10272 8622
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10336 8090 10364 8434
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10244 6730 10364 6746
rect 10244 6724 10376 6730
rect 10244 6718 10324 6724
rect 10324 6666 10376 6672
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 10336 6458 10364 6666
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 9324 6322 9444 6338
rect 9324 6316 9456 6322
rect 9324 6310 9404 6316
rect 9324 5914 9352 6310
rect 9404 6258 9456 6264
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6656 4622 6684 5102
rect 7208 4826 7236 5646
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 7668 5166 7696 5510
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8128 4826 8156 5102
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8404 4622 8432 5510
rect 8864 4690 8892 5646
rect 9140 5370 9168 5646
rect 10336 5642 10364 6394
rect 10428 5778 10456 9522
rect 10796 6390 10824 12174
rect 11532 11218 11560 13262
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11532 10674 11560 11154
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11428 10532 11480 10538
rect 11428 10474 11480 10480
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7002 10916 7686
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11072 6866 11100 8978
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11256 8498 11284 8774
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 8090 11192 8298
rect 11256 8294 11284 8434
rect 11348 8362 11376 9590
rect 11440 8514 11468 10474
rect 11532 9586 11560 10610
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11532 9042 11560 9522
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11440 8486 11560 8514
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11256 8022 11284 8230
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11440 7886 11468 8366
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11256 7546 11284 7822
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9508 5302 9536 5510
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 10520 4554 10548 6326
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10796 5778 10824 6122
rect 11072 5778 11100 6802
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 11532 2774 11560 8486
rect 11624 7410 11652 13398
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 11150 11744 12038
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11808 10690 11836 13874
rect 11992 13802 12020 13874
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 11694 11928 12786
rect 11992 12646 12020 13738
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 12084 12442 12112 12718
rect 12176 12714 12204 13194
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12072 11892 12124 11898
rect 12176 11880 12204 12310
rect 12124 11852 12204 11880
rect 12072 11834 12124 11840
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 12176 11506 12204 11698
rect 12268 11626 12296 13942
rect 12820 13938 12848 14214
rect 12808 13932 12860 13938
rect 12860 13892 12940 13920
rect 12808 13874 12860 13880
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 12918 12572 13670
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12912 12782 12940 13892
rect 15304 13734 15332 22066
rect 15476 22034 15528 22040
rect 15672 22030 15700 23462
rect 15948 23050 15976 23462
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 16224 22642 16252 29446
rect 16500 29306 16528 30330
rect 16488 29300 16540 29306
rect 16488 29242 16540 29248
rect 16488 27872 16540 27878
rect 16488 27814 16540 27820
rect 16302 27160 16358 27169
rect 16302 27095 16304 27104
rect 16356 27095 16358 27104
rect 16304 27066 16356 27072
rect 16304 26988 16356 26994
rect 16304 26930 16356 26936
rect 16316 26586 16344 26930
rect 16304 26580 16356 26586
rect 16304 26522 16356 26528
rect 16394 26480 16450 26489
rect 16394 26415 16396 26424
rect 16448 26415 16450 26424
rect 16396 26386 16448 26392
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 16316 26042 16344 26318
rect 16500 26042 16528 27814
rect 16304 26036 16356 26042
rect 16304 25978 16356 25984
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16396 25968 16448 25974
rect 16396 25910 16448 25916
rect 16408 25702 16436 25910
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 16408 23730 16436 24006
rect 16592 23730 16620 31078
rect 16684 30938 16712 31690
rect 16856 31272 16908 31278
rect 16856 31214 16908 31220
rect 16868 31142 16896 31214
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 16672 30932 16724 30938
rect 16672 30874 16724 30880
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16684 28626 16712 30262
rect 16764 30048 16816 30054
rect 16764 29990 16816 29996
rect 16776 29714 16804 29990
rect 16868 29714 16896 31078
rect 17224 30728 17276 30734
rect 17224 30670 17276 30676
rect 17236 30394 17264 30670
rect 17224 30388 17276 30394
rect 17224 30330 17276 30336
rect 17328 30274 17356 33798
rect 17604 31686 17632 35634
rect 17684 35488 17736 35494
rect 17684 35430 17736 35436
rect 17696 35086 17724 35430
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17788 35018 17816 40054
rect 17880 39982 17908 40990
rect 18800 40526 18828 41074
rect 18880 40996 18932 41002
rect 18880 40938 18932 40944
rect 18892 40526 18920 40938
rect 18788 40520 18840 40526
rect 18788 40462 18840 40468
rect 18880 40520 18932 40526
rect 18880 40462 18932 40468
rect 18696 40452 18748 40458
rect 18696 40394 18748 40400
rect 18236 40384 18288 40390
rect 18236 40326 18288 40332
rect 18248 40186 18276 40326
rect 18236 40180 18288 40186
rect 18236 40122 18288 40128
rect 17868 39976 17920 39982
rect 17868 39918 17920 39924
rect 18144 38276 18196 38282
rect 18144 38218 18196 38224
rect 18156 37806 18184 38218
rect 18144 37800 18196 37806
rect 18144 37742 18196 37748
rect 18156 36650 18184 37742
rect 18144 36644 18196 36650
rect 18144 36586 18196 36592
rect 18052 36576 18104 36582
rect 18052 36518 18104 36524
rect 18064 36242 18092 36518
rect 18052 36236 18104 36242
rect 18052 36178 18104 36184
rect 18156 35290 18184 36586
rect 18248 35630 18276 40122
rect 18708 39438 18736 40394
rect 18800 40118 18828 40462
rect 18892 40390 18920 40462
rect 19444 40390 19472 41482
rect 19904 41414 19932 43250
rect 20168 42696 20220 42702
rect 20168 42638 20220 42644
rect 19984 41540 20036 41546
rect 19984 41482 20036 41488
rect 19812 41386 19932 41414
rect 19524 40452 19576 40458
rect 19524 40394 19576 40400
rect 18880 40384 18932 40390
rect 18880 40326 18932 40332
rect 19432 40384 19484 40390
rect 19432 40326 19484 40332
rect 18788 40112 18840 40118
rect 18788 40054 18840 40060
rect 18892 39982 18920 40326
rect 19444 40050 19472 40326
rect 19432 40044 19484 40050
rect 19432 39986 19484 39992
rect 18880 39976 18932 39982
rect 18880 39918 18932 39924
rect 18788 39840 18840 39846
rect 18788 39782 18840 39788
rect 18800 39506 18828 39782
rect 18788 39500 18840 39506
rect 18788 39442 18840 39448
rect 18696 39432 18748 39438
rect 18696 39374 18748 39380
rect 18708 39098 18736 39374
rect 18696 39092 18748 39098
rect 18696 39034 18748 39040
rect 19340 38820 19392 38826
rect 19340 38762 19392 38768
rect 18420 38752 18472 38758
rect 18420 38694 18472 38700
rect 18432 37942 18460 38694
rect 19352 38350 19380 38762
rect 19340 38344 19392 38350
rect 19340 38286 19392 38292
rect 18788 38276 18840 38282
rect 18788 38218 18840 38224
rect 18420 37936 18472 37942
rect 18420 37878 18472 37884
rect 18328 37868 18380 37874
rect 18328 37810 18380 37816
rect 18340 37466 18368 37810
rect 18800 37754 18828 38218
rect 19064 38208 19116 38214
rect 19064 38150 19116 38156
rect 19076 37942 19104 38150
rect 19064 37936 19116 37942
rect 19064 37878 19116 37884
rect 18708 37738 18828 37754
rect 18696 37732 18828 37738
rect 18748 37726 18828 37732
rect 18696 37674 18748 37680
rect 18328 37460 18380 37466
rect 18328 37402 18380 37408
rect 18800 37233 18828 37726
rect 18786 37224 18842 37233
rect 19352 37210 19380 38286
rect 19444 37670 19472 39986
rect 19432 37664 19484 37670
rect 19432 37606 19484 37612
rect 19444 37330 19472 37606
rect 19536 37398 19564 40394
rect 19708 39296 19760 39302
rect 19708 39238 19760 39244
rect 19720 38962 19748 39238
rect 19708 38956 19760 38962
rect 19708 38898 19760 38904
rect 19708 38208 19760 38214
rect 19708 38150 19760 38156
rect 19524 37392 19576 37398
rect 19524 37334 19576 37340
rect 19432 37324 19484 37330
rect 19720 37274 19748 38150
rect 19432 37266 19484 37272
rect 19524 37256 19576 37262
rect 19352 37182 19472 37210
rect 19524 37198 19576 37204
rect 19628 37246 19748 37274
rect 18786 37159 18842 37168
rect 19444 36802 19472 37182
rect 19536 37126 19564 37198
rect 19524 37120 19576 37126
rect 19524 37062 19576 37068
rect 19076 36786 19472 36802
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 19064 36780 19472 36786
rect 19116 36774 19472 36780
rect 19064 36722 19116 36728
rect 18800 36553 18828 36722
rect 19338 36680 19394 36689
rect 19628 36650 19656 37246
rect 19338 36615 19340 36624
rect 19392 36615 19394 36624
rect 19616 36644 19668 36650
rect 19340 36586 19392 36592
rect 19616 36586 19668 36592
rect 18786 36544 18842 36553
rect 18786 36479 18842 36488
rect 18512 36032 18564 36038
rect 18512 35974 18564 35980
rect 18236 35624 18288 35630
rect 18236 35566 18288 35572
rect 18248 35290 18276 35566
rect 18144 35284 18196 35290
rect 18144 35226 18196 35232
rect 18236 35284 18288 35290
rect 18236 35226 18288 35232
rect 17776 35012 17828 35018
rect 17776 34954 17828 34960
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 17868 32904 17920 32910
rect 17868 32846 17920 32852
rect 17776 32768 17828 32774
rect 17776 32710 17828 32716
rect 17788 32026 17816 32710
rect 17880 32434 17908 32846
rect 18156 32502 18184 33254
rect 18144 32496 18196 32502
rect 18144 32438 18196 32444
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 17776 32020 17828 32026
rect 17776 31962 17828 31968
rect 17592 31680 17644 31686
rect 17592 31622 17644 31628
rect 17604 31482 17632 31622
rect 17592 31476 17644 31482
rect 17592 31418 17644 31424
rect 17408 31136 17460 31142
rect 17406 31104 17408 31113
rect 17460 31104 17462 31113
rect 17406 31039 17462 31048
rect 17788 30818 17816 31962
rect 18144 31748 18196 31754
rect 18144 31690 18196 31696
rect 18156 31346 18184 31690
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 17500 30796 17552 30802
rect 17788 30790 17908 30818
rect 17500 30738 17552 30744
rect 17236 30246 17356 30274
rect 17040 30116 17092 30122
rect 17040 30058 17092 30064
rect 16764 29708 16816 29714
rect 16764 29650 16816 29656
rect 16856 29708 16908 29714
rect 16856 29650 16908 29656
rect 16868 29102 16896 29650
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16856 29096 16908 29102
rect 16856 29038 16908 29044
rect 16672 28620 16724 28626
rect 16672 28562 16724 28568
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 16868 28014 16896 28426
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 16868 27606 16896 27950
rect 16856 27600 16908 27606
rect 16856 27542 16908 27548
rect 16960 27130 16988 29582
rect 17052 29170 17080 30058
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17144 29238 17172 29990
rect 17236 29510 17264 30246
rect 17316 30184 17368 30190
rect 17316 30126 17368 30132
rect 17224 29504 17276 29510
rect 17224 29446 17276 29452
rect 17132 29232 17184 29238
rect 17132 29174 17184 29180
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 17132 29096 17184 29102
rect 17184 29044 17264 29050
rect 17132 29038 17264 29044
rect 17144 29022 17264 29038
rect 17328 29034 17356 30126
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17420 29306 17448 29582
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17144 28150 17172 28494
rect 17132 28144 17184 28150
rect 17132 28086 17184 28092
rect 17040 27396 17092 27402
rect 17040 27338 17092 27344
rect 16764 27124 16816 27130
rect 16764 27066 16816 27072
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 16672 26920 16724 26926
rect 16672 26862 16724 26868
rect 16684 24857 16712 26862
rect 16776 25158 16804 27066
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16868 26450 16896 26930
rect 16948 26920 17000 26926
rect 16946 26888 16948 26897
rect 17000 26888 17002 26897
rect 16946 26823 17002 26832
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 16856 26444 16908 26450
rect 16856 26386 16908 26392
rect 16960 25265 16988 26726
rect 17052 26382 17080 27338
rect 17144 27334 17172 28086
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 17052 25838 17080 26318
rect 17040 25832 17092 25838
rect 17040 25774 17092 25780
rect 16946 25256 17002 25265
rect 17144 25226 17172 27270
rect 17236 27033 17264 29022
rect 17316 29028 17368 29034
rect 17316 28970 17368 28976
rect 17512 28642 17540 30738
rect 17880 30734 17908 30790
rect 17868 30728 17920 30734
rect 17868 30670 17920 30676
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17604 30258 17632 30534
rect 17880 30258 17908 30670
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17684 30252 17736 30258
rect 17684 30194 17736 30200
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17604 29850 17632 30194
rect 17592 29844 17644 29850
rect 17592 29786 17644 29792
rect 17592 29504 17644 29510
rect 17592 29446 17644 29452
rect 17604 29306 17632 29446
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17696 29034 17724 30194
rect 17880 29646 17908 30194
rect 18064 29753 18092 30602
rect 18050 29744 18106 29753
rect 18050 29679 18106 29688
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 17960 29572 18012 29578
rect 17960 29514 18012 29520
rect 17776 29504 17828 29510
rect 17774 29472 17776 29481
rect 17828 29472 17830 29481
rect 17774 29407 17830 29416
rect 17776 29232 17828 29238
rect 17776 29174 17828 29180
rect 17684 29028 17736 29034
rect 17684 28970 17736 28976
rect 17788 28966 17816 29174
rect 17972 29170 18000 29514
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17868 29096 17920 29102
rect 17868 29038 17920 29044
rect 17776 28960 17828 28966
rect 17776 28902 17828 28908
rect 17880 28778 17908 29038
rect 17328 28614 17540 28642
rect 17696 28750 17908 28778
rect 17972 28762 18000 29106
rect 17960 28756 18012 28762
rect 17328 27169 17356 28614
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17420 27452 17448 28494
rect 17696 27713 17724 28750
rect 17960 28698 18012 28704
rect 18064 28642 18092 29679
rect 17788 28614 18092 28642
rect 17682 27704 17738 27713
rect 17682 27639 17738 27648
rect 17788 27588 17816 28614
rect 18156 28558 18184 31282
rect 18248 31142 18276 33458
rect 18236 31136 18288 31142
rect 18236 31078 18288 31084
rect 18420 30592 18472 30598
rect 18420 30534 18472 30540
rect 18432 30054 18460 30534
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 18420 30048 18472 30054
rect 18420 29990 18472 29996
rect 18248 29714 18276 29990
rect 18340 29782 18368 29990
rect 18328 29776 18380 29782
rect 18328 29718 18380 29724
rect 18236 29708 18288 29714
rect 18236 29650 18288 29656
rect 18420 29640 18472 29646
rect 18420 29582 18472 29588
rect 18236 29300 18288 29306
rect 18236 29242 18288 29248
rect 18248 28694 18276 29242
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 18236 28688 18288 28694
rect 18236 28630 18288 28636
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18052 28484 18104 28490
rect 18052 28426 18104 28432
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 17696 27560 17816 27588
rect 17868 27600 17920 27606
rect 17420 27424 17632 27452
rect 17408 27328 17460 27334
rect 17408 27270 17460 27276
rect 17314 27160 17370 27169
rect 17314 27095 17370 27104
rect 17222 27024 17278 27033
rect 17222 26959 17278 26968
rect 17328 26926 17356 27095
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 17420 26518 17448 27270
rect 17498 26888 17554 26897
rect 17498 26823 17500 26832
rect 17552 26823 17554 26832
rect 17500 26794 17552 26800
rect 17604 26602 17632 27424
rect 17696 26790 17724 27560
rect 17868 27542 17920 27548
rect 17776 27396 17828 27402
rect 17776 27338 17828 27344
rect 17788 26994 17816 27338
rect 17880 27169 17908 27542
rect 17972 27470 18000 28154
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 17866 27160 17922 27169
rect 17866 27095 17922 27104
rect 17880 27062 17908 27095
rect 17868 27056 17920 27062
rect 17868 26998 17920 27004
rect 17972 26994 18000 27270
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17604 26574 17724 26602
rect 17408 26512 17460 26518
rect 17408 26454 17460 26460
rect 17420 26382 17448 26454
rect 17224 26376 17276 26382
rect 17222 26344 17224 26353
rect 17408 26376 17460 26382
rect 17276 26344 17278 26353
rect 17408 26318 17460 26324
rect 17222 26279 17278 26288
rect 17592 26240 17644 26246
rect 17592 26182 17644 26188
rect 16946 25191 17002 25200
rect 17132 25220 17184 25226
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16670 24848 16726 24857
rect 16670 24783 16726 24792
rect 16684 24138 16712 24783
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16776 24070 16804 25094
rect 16960 24206 16988 25191
rect 17132 25162 17184 25168
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 17052 24274 17080 24550
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 17236 24206 17264 24890
rect 17604 24886 17632 26182
rect 17696 25378 17724 26574
rect 17788 26314 17816 26726
rect 17972 26586 18000 26930
rect 17960 26580 18012 26586
rect 17960 26522 18012 26528
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17788 25498 17816 26250
rect 17868 26240 17920 26246
rect 17868 26182 17920 26188
rect 17880 25770 17908 26182
rect 17972 25906 18000 26318
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17868 25764 17920 25770
rect 17868 25706 17920 25712
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17696 25350 17908 25378
rect 17880 25226 17908 25350
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 17960 25220 18012 25226
rect 17960 25162 18012 25168
rect 17592 24880 17644 24886
rect 17592 24822 17644 24828
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16396 23724 16448 23730
rect 16396 23666 16448 23672
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 16776 23474 16804 24006
rect 17130 23760 17186 23769
rect 17040 23724 17092 23730
rect 17604 23730 17632 24822
rect 17880 23905 17908 25162
rect 17972 24410 18000 25162
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 17866 23896 17922 23905
rect 17866 23831 17922 23840
rect 17972 23730 18000 24346
rect 18064 23866 18092 28426
rect 18248 28082 18276 28494
rect 18340 28218 18368 28902
rect 18328 28212 18380 28218
rect 18432 28200 18460 29582
rect 18524 28626 18552 35974
rect 18604 35760 18656 35766
rect 18604 35702 18656 35708
rect 18616 35086 18644 35702
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 18616 34610 18644 35022
rect 19156 34944 19208 34950
rect 19156 34886 19208 34892
rect 19168 34746 19196 34886
rect 19156 34740 19208 34746
rect 19156 34682 19208 34688
rect 19248 34740 19300 34746
rect 19248 34682 19300 34688
rect 18604 34604 18656 34610
rect 18604 34546 18656 34552
rect 18616 34066 18644 34546
rect 19260 34542 19288 34682
rect 19340 34604 19392 34610
rect 19340 34546 19392 34552
rect 19248 34536 19300 34542
rect 19248 34478 19300 34484
rect 19260 34202 19288 34478
rect 19248 34196 19300 34202
rect 19248 34138 19300 34144
rect 18604 34060 18656 34066
rect 18604 34002 18656 34008
rect 18616 33658 18644 34002
rect 18604 33652 18656 33658
rect 18604 33594 18656 33600
rect 18788 33516 18840 33522
rect 18788 33458 18840 33464
rect 18972 33516 19024 33522
rect 18972 33458 19024 33464
rect 18800 33114 18828 33458
rect 18788 33108 18840 33114
rect 18788 33050 18840 33056
rect 18604 32360 18656 32366
rect 18604 32302 18656 32308
rect 18616 31754 18644 32302
rect 18604 31748 18656 31754
rect 18604 31690 18656 31696
rect 18880 30864 18932 30870
rect 18880 30806 18932 30812
rect 18788 30728 18840 30734
rect 18892 30716 18920 30806
rect 18840 30688 18920 30716
rect 18788 30670 18840 30676
rect 18694 30152 18750 30161
rect 18694 30087 18696 30096
rect 18748 30087 18750 30096
rect 18696 30058 18748 30064
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18616 28762 18644 29582
rect 18696 29572 18748 29578
rect 18696 29514 18748 29520
rect 18708 29238 18736 29514
rect 18696 29232 18748 29238
rect 18696 29174 18748 29180
rect 18696 29028 18748 29034
rect 18696 28970 18748 28976
rect 18604 28756 18656 28762
rect 18604 28698 18656 28704
rect 18512 28620 18564 28626
rect 18512 28562 18564 28568
rect 18708 28393 18736 28970
rect 18788 28688 18840 28694
rect 18788 28630 18840 28636
rect 18694 28384 18750 28393
rect 18694 28319 18750 28328
rect 18432 28172 18736 28200
rect 18328 28154 18380 28160
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18420 28008 18472 28014
rect 18420 27950 18472 27956
rect 18236 27668 18288 27674
rect 18236 27610 18288 27616
rect 18248 27538 18276 27610
rect 18432 27606 18460 27950
rect 18420 27600 18472 27606
rect 18420 27542 18472 27548
rect 18236 27532 18288 27538
rect 18236 27474 18288 27480
rect 18144 27328 18196 27334
rect 18144 27270 18196 27276
rect 18156 26994 18184 27270
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 18156 26450 18184 26930
rect 18248 26908 18276 27474
rect 18328 27328 18380 27334
rect 18328 27270 18380 27276
rect 18340 27130 18368 27270
rect 18328 27124 18380 27130
rect 18328 27066 18380 27072
rect 18432 26994 18460 27542
rect 18524 27334 18552 28018
rect 18708 27946 18736 28172
rect 18696 27940 18748 27946
rect 18696 27882 18748 27888
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 18328 26920 18380 26926
rect 18248 26880 18328 26908
rect 18248 26450 18276 26880
rect 18328 26862 18380 26868
rect 18328 26512 18380 26518
rect 18328 26454 18380 26460
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 18236 26036 18288 26042
rect 18236 25978 18288 25984
rect 18144 25492 18196 25498
rect 18144 25434 18196 25440
rect 18156 24750 18184 25434
rect 18248 25294 18276 25978
rect 18340 25770 18368 26454
rect 18524 26382 18552 27270
rect 18616 26858 18644 27270
rect 18604 26852 18656 26858
rect 18604 26794 18656 26800
rect 18708 26790 18736 27882
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 18432 26217 18460 26318
rect 18418 26208 18474 26217
rect 18418 26143 18474 26152
rect 18328 25764 18380 25770
rect 18328 25706 18380 25712
rect 18340 25362 18368 25706
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18420 25152 18472 25158
rect 18420 25094 18472 25100
rect 18432 24818 18460 25094
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 18328 24676 18380 24682
rect 18328 24618 18380 24624
rect 18340 24342 18368 24618
rect 18432 24585 18460 24754
rect 18604 24608 18656 24614
rect 18418 24576 18474 24585
rect 18604 24550 18656 24556
rect 18418 24511 18474 24520
rect 18328 24336 18380 24342
rect 18328 24278 18380 24284
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 17130 23695 17186 23704
rect 17592 23724 17644 23730
rect 17040 23666 17092 23672
rect 16500 23446 16804 23474
rect 16500 22778 16528 23446
rect 17052 23254 17080 23666
rect 17144 23662 17172 23695
rect 17592 23666 17644 23672
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 18064 23594 18092 23802
rect 18052 23588 18104 23594
rect 18052 23530 18104 23536
rect 17960 23520 18012 23526
rect 17590 23488 17646 23497
rect 17960 23462 18012 23468
rect 17590 23423 17646 23432
rect 17040 23248 17092 23254
rect 16868 23196 17040 23202
rect 16868 23190 17092 23196
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16868 23174 17080 23190
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16212 22636 16264 22642
rect 16212 22578 16264 22584
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16408 22234 16436 22374
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16304 22092 16356 22098
rect 16304 22034 16356 22040
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15396 21554 15424 21898
rect 15580 21690 15608 21966
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15580 20534 15608 20742
rect 15568 20528 15620 20534
rect 15568 20470 15620 20476
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15488 16590 15516 17614
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15396 16114 15424 16458
rect 15672 16250 15700 21966
rect 16316 21894 16344 22034
rect 16408 22030 16436 22170
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16316 21554 16344 21830
rect 16592 21622 16620 22918
rect 16684 22574 16712 23122
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16684 22098 16712 22510
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16580 21616 16632 21622
rect 16580 21558 16632 21564
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16132 21146 16160 21422
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16026 21040 16082 21049
rect 16026 20975 16028 20984
rect 16080 20975 16082 20984
rect 16028 20946 16080 20952
rect 16132 20466 16160 21082
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16592 20398 16620 20878
rect 16684 20466 16712 22034
rect 16868 21962 16896 23174
rect 17604 22710 17632 23423
rect 17592 22704 17644 22710
rect 17592 22646 17644 22652
rect 17972 22642 18000 23462
rect 18156 23118 18184 24210
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 18064 22778 18092 22986
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17512 22234 17540 22374
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 16948 22160 17000 22166
rect 16948 22102 17000 22108
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 16960 21622 16988 22102
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 17236 20942 17264 21626
rect 18064 21554 18092 22714
rect 18156 22642 18184 23054
rect 18248 22642 18276 24074
rect 18340 23730 18368 24278
rect 18616 24274 18644 24550
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18512 24200 18564 24206
rect 18510 24168 18512 24177
rect 18564 24168 18566 24177
rect 18510 24103 18566 24112
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18432 23866 18460 24006
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 18616 23662 18644 24210
rect 18800 24206 18828 28630
rect 18892 27674 18920 30688
rect 18984 29306 19012 33458
rect 19352 31754 19380 34546
rect 19812 34082 19840 41386
rect 19996 37788 20024 41482
rect 20076 38752 20128 38758
rect 20076 38694 20128 38700
rect 20088 38418 20116 38694
rect 20076 38412 20128 38418
rect 20076 38354 20128 38360
rect 20180 38026 20208 42638
rect 20444 42560 20496 42566
rect 20444 42502 20496 42508
rect 20260 42288 20312 42294
rect 20260 42230 20312 42236
rect 20272 41478 20300 42230
rect 20260 41472 20312 41478
rect 20260 41414 20312 41420
rect 20352 40996 20404 41002
rect 20352 40938 20404 40944
rect 20364 40730 20392 40938
rect 20352 40724 20404 40730
rect 20352 40666 20404 40672
rect 20364 40458 20392 40666
rect 20352 40452 20404 40458
rect 20352 40394 20404 40400
rect 20260 39024 20312 39030
rect 20260 38966 20312 38972
rect 20352 39024 20404 39030
rect 20352 38966 20404 38972
rect 20272 38282 20300 38966
rect 20364 38282 20392 38966
rect 20260 38276 20312 38282
rect 20260 38218 20312 38224
rect 20352 38276 20404 38282
rect 20352 38218 20404 38224
rect 20180 37998 20300 38026
rect 20076 37800 20128 37806
rect 19996 37760 20076 37788
rect 20076 37742 20128 37748
rect 19984 37392 20036 37398
rect 19984 37334 20036 37340
rect 19892 37120 19944 37126
rect 19892 37062 19944 37068
rect 19904 36786 19932 37062
rect 19892 36780 19944 36786
rect 19892 36722 19944 36728
rect 19904 36689 19932 36722
rect 19890 36680 19946 36689
rect 19890 36615 19946 36624
rect 19892 36576 19944 36582
rect 19892 36518 19944 36524
rect 19904 36378 19932 36518
rect 19892 36372 19944 36378
rect 19892 36314 19944 36320
rect 19996 35698 20024 37334
rect 20088 37194 20116 37742
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20076 37188 20128 37194
rect 20076 37130 20128 37136
rect 20180 36666 20208 37198
rect 20272 36922 20300 37998
rect 20260 36916 20312 36922
rect 20260 36858 20312 36864
rect 20180 36638 20300 36666
rect 20168 36576 20220 36582
rect 20166 36544 20168 36553
rect 20220 36544 20222 36553
rect 20166 36479 20222 36488
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 19720 34054 19840 34082
rect 19720 33096 19748 34054
rect 19800 33924 19852 33930
rect 19800 33866 19852 33872
rect 19812 33658 19840 33866
rect 19800 33652 19852 33658
rect 19800 33594 19852 33600
rect 19800 33516 19852 33522
rect 19800 33458 19852 33464
rect 19536 33068 19748 33096
rect 19536 32842 19564 33068
rect 19616 32972 19668 32978
rect 19616 32914 19668 32920
rect 19524 32836 19576 32842
rect 19524 32778 19576 32784
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19156 31408 19208 31414
rect 19156 31350 19208 31356
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 19076 30190 19104 30670
rect 19168 30598 19196 31350
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 19156 30252 19208 30258
rect 19156 30194 19208 30200
rect 19064 30184 19116 30190
rect 19064 30126 19116 30132
rect 19076 29730 19104 30126
rect 19168 29850 19196 30194
rect 19156 29844 19208 29850
rect 19156 29786 19208 29792
rect 19076 29702 19196 29730
rect 18972 29300 19024 29306
rect 18972 29242 19024 29248
rect 19064 29096 19116 29102
rect 19064 29038 19116 29044
rect 19076 28558 19104 29038
rect 19168 28642 19196 29702
rect 19249 29300 19301 29306
rect 19249 29242 19301 29248
rect 19260 29050 19288 29242
rect 19260 29022 19289 29050
rect 19261 28994 19289 29022
rect 19260 28966 19289 28994
rect 19260 28762 19288 28966
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19168 28614 19288 28642
rect 18972 28552 19024 28558
rect 18972 28494 19024 28500
rect 19064 28552 19116 28558
rect 19064 28494 19116 28500
rect 18984 27860 19012 28494
rect 19076 28014 19104 28494
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 19168 27860 19196 28018
rect 18984 27832 19196 27860
rect 18880 27668 18932 27674
rect 18880 27610 18932 27616
rect 18892 27062 18920 27610
rect 19168 27538 19196 27832
rect 19156 27532 19208 27538
rect 19156 27474 19208 27480
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 18880 27056 18932 27062
rect 18880 26998 18932 27004
rect 18972 26988 19024 26994
rect 18972 26930 19024 26936
rect 18984 26518 19012 26930
rect 19076 26897 19104 27270
rect 19168 26994 19196 27474
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 19062 26888 19118 26897
rect 19062 26823 19118 26832
rect 18972 26512 19024 26518
rect 18972 26454 19024 26460
rect 19168 26217 19196 26930
rect 19154 26208 19210 26217
rect 19154 26143 19210 26152
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 18788 24200 18840 24206
rect 19064 24200 19116 24206
rect 18840 24148 19064 24154
rect 18788 24142 19116 24148
rect 18800 24126 19104 24142
rect 19168 24070 19196 24346
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 18800 23730 18828 24006
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 19260 23662 19288 28614
rect 19352 24954 19380 31690
rect 19524 31680 19576 31686
rect 19524 31622 19576 31628
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19444 30394 19472 30738
rect 19536 30598 19564 31622
rect 19628 31346 19656 32914
rect 19720 32366 19748 33068
rect 19708 32360 19760 32366
rect 19708 32302 19760 32308
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19616 31340 19668 31346
rect 19616 31282 19668 31288
rect 19720 31278 19748 31826
rect 19708 31272 19760 31278
rect 19708 31214 19760 31220
rect 19708 30864 19760 30870
rect 19706 30832 19708 30841
rect 19760 30832 19762 30841
rect 19706 30767 19762 30776
rect 19616 30728 19668 30734
rect 19616 30670 19668 30676
rect 19708 30728 19760 30734
rect 19708 30670 19760 30676
rect 19524 30592 19576 30598
rect 19524 30534 19576 30540
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19536 30274 19564 30534
rect 19628 30394 19656 30670
rect 19616 30388 19668 30394
rect 19616 30330 19668 30336
rect 19444 30246 19564 30274
rect 19444 29170 19472 30246
rect 19720 29850 19748 30670
rect 19812 30122 19840 33458
rect 20076 32836 20128 32842
rect 20076 32778 20128 32784
rect 20088 32502 20116 32778
rect 20076 32496 20128 32502
rect 20076 32438 20128 32444
rect 19892 30932 19944 30938
rect 19892 30874 19944 30880
rect 19904 30802 19932 30874
rect 20272 30870 20300 36638
rect 20456 36378 20484 42502
rect 20536 40996 20588 41002
rect 20536 40938 20588 40944
rect 20812 40996 20864 41002
rect 20812 40938 20864 40944
rect 20548 40662 20576 40938
rect 20536 40656 20588 40662
rect 20536 40598 20588 40604
rect 20720 40384 20772 40390
rect 20720 40326 20772 40332
rect 20732 40050 20760 40326
rect 20720 40044 20772 40050
rect 20720 39986 20772 39992
rect 20824 39982 20852 40938
rect 20812 39976 20864 39982
rect 20812 39918 20864 39924
rect 20812 38956 20864 38962
rect 20812 38898 20864 38904
rect 20628 38820 20680 38826
rect 20628 38762 20680 38768
rect 20536 38752 20588 38758
rect 20536 38694 20588 38700
rect 20548 38350 20576 38694
rect 20536 38344 20588 38350
rect 20536 38286 20588 38292
rect 20640 37942 20668 38762
rect 20720 38276 20772 38282
rect 20720 38218 20772 38224
rect 20628 37936 20680 37942
rect 20628 37878 20680 37884
rect 20536 37868 20588 37874
rect 20536 37810 20588 37816
rect 20548 37670 20576 37810
rect 20536 37664 20588 37670
rect 20536 37606 20588 37612
rect 20444 36372 20496 36378
rect 20444 36314 20496 36320
rect 20548 35850 20576 37606
rect 20732 37126 20760 38218
rect 20824 37738 20852 38898
rect 20916 37754 20944 43250
rect 21100 42294 21128 43250
rect 21180 43240 21232 43246
rect 21180 43182 21232 43188
rect 21088 42288 21140 42294
rect 21088 42230 21140 42236
rect 21100 41682 21128 42230
rect 21088 41676 21140 41682
rect 21088 41618 21140 41624
rect 21088 41472 21140 41478
rect 21088 41414 21140 41420
rect 21192 41414 21220 43182
rect 21548 43104 21600 43110
rect 21548 43046 21600 43052
rect 21456 42696 21508 42702
rect 21456 42638 21508 42644
rect 21468 42362 21496 42638
rect 21456 42356 21508 42362
rect 21456 42298 21508 42304
rect 21468 41682 21496 42298
rect 21456 41676 21508 41682
rect 21456 41618 21508 41624
rect 21100 41138 21128 41414
rect 21192 41386 21404 41414
rect 21088 41132 21140 41138
rect 21088 41074 21140 41080
rect 21100 41018 21128 41074
rect 21008 40990 21128 41018
rect 21272 40996 21324 41002
rect 21008 40526 21036 40990
rect 21272 40938 21324 40944
rect 21180 40928 21232 40934
rect 21180 40870 21232 40876
rect 20996 40520 21048 40526
rect 20996 40462 21048 40468
rect 21192 40118 21220 40870
rect 21284 40526 21312 40938
rect 21272 40520 21324 40526
rect 21272 40462 21324 40468
rect 21180 40112 21232 40118
rect 21180 40054 21232 40060
rect 21088 39908 21140 39914
rect 21088 39850 21140 39856
rect 21100 39030 21128 39850
rect 21088 39024 21140 39030
rect 21088 38966 21140 38972
rect 20996 38548 21048 38554
rect 20996 38490 21048 38496
rect 21008 38298 21036 38490
rect 21100 38418 21128 38966
rect 21272 38480 21324 38486
rect 21272 38422 21324 38428
rect 21088 38412 21140 38418
rect 21088 38354 21140 38360
rect 21008 38270 21128 38298
rect 20996 38208 21048 38214
rect 20996 38150 21048 38156
rect 21008 37874 21036 38150
rect 20996 37868 21048 37874
rect 20996 37810 21048 37816
rect 21100 37754 21128 38270
rect 21180 38208 21232 38214
rect 21180 38150 21232 38156
rect 21192 37874 21220 38150
rect 21284 37874 21312 38422
rect 21180 37868 21232 37874
rect 21180 37810 21232 37816
rect 21272 37868 21324 37874
rect 21272 37810 21324 37816
rect 20812 37732 20864 37738
rect 20916 37726 21036 37754
rect 21100 37726 21220 37754
rect 20812 37674 20864 37680
rect 20824 37194 20852 37674
rect 20904 37664 20956 37670
rect 20904 37606 20956 37612
rect 20916 37330 20944 37606
rect 20904 37324 20956 37330
rect 20904 37266 20956 37272
rect 20812 37188 20864 37194
rect 20812 37130 20864 37136
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 20812 36712 20864 36718
rect 20812 36654 20864 36660
rect 20824 36122 20852 36654
rect 20824 36094 20944 36122
rect 20916 36038 20944 36094
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 20456 35822 20576 35850
rect 20352 32020 20404 32026
rect 20352 31962 20404 31968
rect 20260 30864 20312 30870
rect 19982 30832 20038 30841
rect 19892 30796 19944 30802
rect 20260 30806 20312 30812
rect 19982 30767 19984 30776
rect 19892 30738 19944 30744
rect 20036 30767 20038 30776
rect 19984 30738 20036 30744
rect 19892 30660 19944 30666
rect 19892 30602 19944 30608
rect 19904 30258 19932 30602
rect 19984 30388 20036 30394
rect 20036 30348 20208 30376
rect 19984 30330 20036 30336
rect 19892 30252 19944 30258
rect 19892 30194 19944 30200
rect 19800 30116 19852 30122
rect 19800 30058 19852 30064
rect 19708 29844 19760 29850
rect 19708 29786 19760 29792
rect 19800 29708 19852 29714
rect 19800 29650 19852 29656
rect 19524 29640 19576 29646
rect 19524 29582 19576 29588
rect 19536 29481 19564 29582
rect 19616 29504 19668 29510
rect 19522 29472 19578 29481
rect 19616 29446 19668 29452
rect 19522 29407 19578 29416
rect 19628 29170 19656 29446
rect 19812 29170 19840 29650
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19616 29164 19668 29170
rect 19616 29106 19668 29112
rect 19800 29164 19852 29170
rect 19800 29106 19852 29112
rect 19444 28558 19472 29106
rect 19524 29096 19576 29102
rect 19524 29038 19576 29044
rect 19432 28552 19484 28558
rect 19432 28494 19484 28500
rect 19430 28384 19486 28393
rect 19430 28319 19486 28328
rect 19444 27674 19472 28319
rect 19536 28218 19564 29038
rect 19616 29028 19668 29034
rect 19616 28970 19668 28976
rect 19628 28490 19656 28970
rect 19616 28484 19668 28490
rect 19616 28426 19668 28432
rect 19524 28212 19576 28218
rect 19524 28154 19576 28160
rect 19524 27872 19576 27878
rect 19524 27814 19576 27820
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19536 27130 19564 27814
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19444 25906 19472 27066
rect 19536 26246 19564 27066
rect 19524 26240 19576 26246
rect 19524 26182 19576 26188
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19536 25838 19564 26182
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19628 24954 19656 28426
rect 19340 24948 19392 24954
rect 19616 24948 19668 24954
rect 19392 24908 19564 24936
rect 19340 24890 19392 24896
rect 19536 24834 19564 24908
rect 19616 24890 19668 24896
rect 19536 24806 19656 24834
rect 19524 24744 19576 24750
rect 19352 24704 19524 24732
rect 19352 24070 19380 24704
rect 19524 24686 19576 24692
rect 19522 24440 19578 24449
rect 19522 24375 19578 24384
rect 19536 24274 19564 24375
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 19432 24200 19484 24206
rect 19430 24168 19432 24177
rect 19484 24168 19486 24177
rect 19430 24103 19486 24112
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19352 23662 19380 24006
rect 19444 23798 19472 24103
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18248 22234 18276 22578
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 17972 21350 18000 21422
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 15764 19514 15792 19722
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 16224 16522 16252 19722
rect 17144 19514 17172 20198
rect 17328 20058 17356 20334
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17236 18834 17264 19654
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16684 17678 16712 18022
rect 17052 17746 17080 18226
rect 17420 18222 17448 20946
rect 17972 20942 18000 21286
rect 18156 20942 18184 21830
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18248 20874 18276 22170
rect 18512 21956 18564 21962
rect 18512 21898 18564 21904
rect 18524 21554 18552 21898
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18524 20924 18552 21490
rect 18432 20896 18552 20924
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17788 19514 17816 19654
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17408 18216 17460 18222
rect 17328 18176 17408 18204
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 17052 16726 17080 17478
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 16212 16516 16264 16522
rect 16212 16458 16264 16464
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 17130 16144 17186 16153
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 15844 16108 15896 16114
rect 17130 16079 17132 16088
rect 15844 16050 15896 16056
rect 17184 16079 17186 16088
rect 17132 16050 17184 16056
rect 15856 15910 15884 16050
rect 17328 16046 17356 18176
rect 17408 18158 17460 18164
rect 17696 17746 17724 19110
rect 17788 18970 17816 19450
rect 17972 19446 18000 20334
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17972 18290 18000 19382
rect 18064 18834 18092 19858
rect 18432 19854 18460 20896
rect 18616 20602 18644 23462
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18800 22710 18828 22918
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18892 21554 18920 21966
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19168 21146 19196 21490
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18616 19922 18644 20538
rect 19076 20534 19104 20742
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18432 19446 18460 19790
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18420 19440 18472 19446
rect 18420 19382 18472 19388
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18340 18970 18368 19246
rect 18432 18970 18460 19382
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18432 18358 18460 18906
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18432 17882 18460 18158
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 17338 17448 17478
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18156 16590 18184 17070
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15396 15026 15424 15846
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13530 15332 13670
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12440 12368 12492 12374
rect 12360 12316 12440 12322
rect 12360 12310 12492 12316
rect 12360 12294 12480 12310
rect 12360 11762 12388 12294
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12452 11898 12480 12174
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12820 11898 12848 12106
rect 12912 12102 12940 12718
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 11900 11014 11928 11494
rect 12176 11478 12480 11506
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11716 10662 11836 10690
rect 11716 10130 11744 10662
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11808 10266 11836 10542
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 12084 10130 12112 10950
rect 12452 10606 12480 11478
rect 12544 11354 12572 11766
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12544 10962 12572 11086
rect 12636 10962 12664 11698
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12820 11082 12848 11562
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12820 10962 12848 11018
rect 12544 10934 12848 10962
rect 12820 10810 12848 10934
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12912 10538 12940 12038
rect 13004 11218 13032 13126
rect 13464 12918 13492 13126
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13372 12306 13400 12854
rect 13464 12442 13492 12854
rect 13740 12850 13768 13126
rect 14568 12918 14596 13262
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14936 12918 14964 13194
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13372 11898 13400 12242
rect 13556 12238 13584 12582
rect 13648 12238 13676 12650
rect 15028 12442 15056 12718
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13176 11824 13228 11830
rect 13096 11784 13176 11812
rect 13096 11354 13124 11784
rect 13176 11766 13228 11772
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13188 11558 13216 11630
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 13004 10826 13032 11154
rect 13188 11014 13216 11494
rect 13372 11370 13400 11630
rect 13280 11342 13400 11370
rect 13464 11354 13492 11698
rect 13452 11348 13504 11354
rect 13280 11014 13308 11342
rect 13452 11290 13504 11296
rect 13648 11218 13676 12174
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11354 13768 11494
rect 13924 11354 13952 11630
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14016 11218 14044 11766
rect 14568 11762 14596 12038
rect 15120 11898 15148 12854
rect 15856 12238 15884 15846
rect 16500 15162 16528 15982
rect 17328 15910 17356 15982
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 16684 15434 16712 15846
rect 17420 15434 17448 15982
rect 17512 15706 17540 16526
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18156 15910 18184 16390
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14346 16252 14758
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16408 13394 16436 13670
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16500 12850 16528 13738
rect 16592 12986 16620 14962
rect 17052 14958 17080 15370
rect 18050 15192 18106 15201
rect 18156 15162 18184 15846
rect 18248 15502 18276 16186
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18050 15127 18106 15136
rect 18144 15156 18196 15162
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16948 14476 17000 14482
rect 17052 14464 17080 14894
rect 17972 14618 18000 14962
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17000 14436 17080 14464
rect 16948 14418 17000 14424
rect 17052 13870 17080 14436
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17052 13326 17080 13806
rect 17972 13734 18000 14214
rect 18064 13938 18092 15127
rect 18144 15098 18196 15104
rect 18340 14958 18368 17682
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 15706 18460 16390
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18340 14550 18368 14894
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18432 14074 18460 14894
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18524 14006 18552 14282
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 11354 14504 11630
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13004 10798 13124 10826
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11716 9042 11744 10066
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12176 9178 12204 9454
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11716 7886 11744 8774
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11808 7886 11836 8026
rect 11900 7954 11928 8570
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11900 7342 11928 7890
rect 12084 7750 12112 8502
rect 12176 8090 12204 8502
rect 12268 8430 12296 9386
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8566 12388 8910
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12820 8498 12848 8978
rect 13004 8838 13032 10798
rect 13096 10742 13124 10798
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 13188 10452 13216 10950
rect 13280 10606 13308 10950
rect 14016 10810 14044 11154
rect 15120 11082 15148 11834
rect 15856 11762 15884 12174
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13268 10464 13320 10470
rect 13188 10424 13268 10452
rect 13268 10406 13320 10412
rect 13280 10130 13308 10406
rect 13372 10266 13400 10610
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13648 10130 13676 10542
rect 13740 10266 13768 10746
rect 14464 10736 14516 10742
rect 14568 10690 14596 11018
rect 15488 10742 15516 11494
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 14516 10684 14596 10690
rect 14464 10678 14596 10684
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 14476 10662 14596 10678
rect 15764 10674 15792 11154
rect 16132 11150 16160 12038
rect 16500 11694 16528 12786
rect 17880 12714 17908 13126
rect 17868 12708 17920 12714
rect 17868 12650 17920 12656
rect 17880 12238 17908 12650
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16592 11762 16620 12106
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16500 11218 16528 11630
rect 17604 11354 17632 12174
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13740 10062 13768 10202
rect 13924 10130 13952 10406
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 14568 9994 14596 10662
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13004 8566 13032 8774
rect 13096 8634 13124 8910
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 13096 8498 13124 8570
rect 13188 8498 13216 8842
rect 14568 8566 14596 9930
rect 15856 9042 15884 9998
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7478 12112 7686
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 12176 7410 12204 8026
rect 12452 7546 12480 8298
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 7750 12848 8230
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12820 7410 12848 7686
rect 13188 7478 13216 8434
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13556 7546 13584 7754
rect 14568 7750 14596 8502
rect 15304 8430 15332 8978
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15304 7954 15332 8366
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 18064 7750 18092 13874
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18524 13394 18552 13806
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18432 12986 18460 13330
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18156 8566 18184 12922
rect 18616 12434 18644 19722
rect 19260 19310 19288 23598
rect 19536 23186 19564 24006
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19628 23050 19656 24806
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19720 23866 19748 24142
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19812 23798 19840 29106
rect 19904 28778 19932 30194
rect 20180 30190 20208 30348
rect 20168 30184 20220 30190
rect 20168 30126 20220 30132
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 19904 28750 20024 28778
rect 19892 26988 19944 26994
rect 19892 26930 19944 26936
rect 19904 26314 19932 26930
rect 19892 26308 19944 26314
rect 19892 26250 19944 26256
rect 19892 24404 19944 24410
rect 19892 24346 19944 24352
rect 19904 24138 19932 24346
rect 19996 24274 20024 28750
rect 20088 28082 20116 29582
rect 20180 28694 20208 30126
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 20272 29102 20300 29582
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20168 28688 20220 28694
rect 20168 28630 20220 28636
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 20258 27568 20314 27577
rect 20088 27402 20116 27542
rect 20258 27503 20314 27512
rect 20076 27396 20128 27402
rect 20076 27338 20128 27344
rect 20088 25888 20116 27338
rect 20272 26897 20300 27503
rect 20258 26888 20314 26897
rect 20258 26823 20260 26832
rect 20312 26823 20314 26832
rect 20260 26794 20312 26800
rect 20260 26444 20312 26450
rect 20260 26386 20312 26392
rect 20168 25900 20220 25906
rect 20088 25860 20168 25888
rect 20168 25842 20220 25848
rect 20272 25838 20300 26386
rect 20260 25832 20312 25838
rect 20260 25774 20312 25780
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19800 23792 19852 23798
rect 19800 23734 19852 23740
rect 19892 23588 19944 23594
rect 19892 23530 19944 23536
rect 19904 23186 19932 23530
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19616 23044 19668 23050
rect 19616 22986 19668 22992
rect 19628 22778 19656 22986
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19352 20058 19380 20878
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19812 19854 19840 22714
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19260 18766 19288 19246
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19800 18692 19852 18698
rect 19800 18634 19852 18640
rect 19340 18624 19392 18630
rect 19720 18601 19748 18634
rect 19340 18566 19392 18572
rect 19706 18592 19762 18601
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 18708 15570 18736 16526
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18800 15502 18828 16390
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18800 14890 18828 15438
rect 18892 15366 18920 15642
rect 18984 15434 19012 16526
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19168 15638 19196 16390
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 19076 15162 19104 15506
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18892 14822 18920 14962
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18788 14408 18840 14414
rect 18892 14396 18920 14758
rect 18840 14368 18920 14396
rect 18788 14350 18840 14356
rect 19076 14328 19104 15098
rect 19260 14822 19288 15574
rect 19352 15162 19380 18566
rect 19706 18527 19762 18536
rect 19720 18290 19748 18527
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19812 17762 19840 18634
rect 19996 18426 20024 24210
rect 20088 23730 20116 24618
rect 20180 23798 20208 24754
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20272 23866 20300 24006
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 20180 23526 20208 23734
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20088 20262 20116 20878
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19628 17740 19840 17762
rect 19628 17734 19708 17740
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19444 15706 19472 16050
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19156 14340 19208 14346
rect 19076 14300 19156 14328
rect 19156 14282 19208 14288
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18800 13462 18828 13806
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 19444 12850 19472 14486
rect 19536 13258 19564 16458
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19352 12646 19380 12718
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 18616 12406 19012 12434
rect 18984 11286 19012 12406
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19168 11898 19196 12174
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18340 10606 18368 11086
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18616 10742 18644 10950
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18340 10062 18368 10542
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18340 9568 18368 9998
rect 18420 9580 18472 9586
rect 18340 9540 18420 9568
rect 18420 9522 18472 9528
rect 18328 9036 18380 9042
rect 18432 9024 18460 9522
rect 19352 9042 19380 12582
rect 19444 11694 19472 12786
rect 19628 12714 19656 17734
rect 19760 17734 19840 17740
rect 19892 17740 19944 17746
rect 19708 17682 19760 17688
rect 19892 17682 19944 17688
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 16590 19748 17478
rect 19904 17202 19932 17682
rect 19996 17678 20024 18362
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19720 16182 19748 16526
rect 19708 16176 19760 16182
rect 19708 16118 19760 16124
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19720 14414 19748 15098
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19720 13326 19748 14350
rect 19812 14226 19840 16526
rect 19892 16516 19944 16522
rect 19892 16458 19944 16464
rect 19904 15706 19932 16458
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19904 15026 19932 15302
rect 19996 15162 20024 16050
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19984 14272 20036 14278
rect 19812 14198 19932 14226
rect 19984 14214 20036 14220
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19616 12708 19668 12714
rect 19616 12650 19668 12656
rect 19812 12170 19840 14010
rect 19904 13326 19932 14198
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19904 12986 19932 13262
rect 19996 13258 20024 14214
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 20088 13138 20116 20198
rect 20364 18358 20392 31962
rect 20456 30734 20484 35822
rect 20916 35562 20944 35974
rect 20904 35556 20956 35562
rect 20904 35498 20956 35504
rect 20536 35488 20588 35494
rect 20536 35430 20588 35436
rect 20548 34678 20576 35430
rect 20916 34746 20944 35498
rect 20904 34740 20956 34746
rect 20904 34682 20956 34688
rect 20536 34672 20588 34678
rect 20536 34614 20588 34620
rect 21008 34202 21036 37726
rect 21192 36718 21220 37726
rect 21376 37346 21404 41386
rect 21468 41002 21496 41618
rect 21560 41546 21588 43046
rect 21652 42226 21680 43318
rect 23112 43308 23164 43314
rect 23112 43250 23164 43256
rect 23756 43308 23808 43314
rect 23756 43250 23808 43256
rect 22008 42628 22060 42634
rect 22008 42570 22060 42576
rect 21640 42220 21692 42226
rect 21640 42162 21692 42168
rect 21548 41540 21600 41546
rect 21548 41482 21600 41488
rect 21560 41138 21588 41482
rect 21652 41138 21680 42162
rect 21916 42016 21968 42022
rect 21916 41958 21968 41964
rect 21928 41614 21956 41958
rect 21916 41608 21968 41614
rect 21916 41550 21968 41556
rect 21548 41132 21600 41138
rect 21548 41074 21600 41080
rect 21640 41132 21692 41138
rect 21640 41074 21692 41080
rect 21456 40996 21508 41002
rect 21456 40938 21508 40944
rect 21456 38956 21508 38962
rect 21456 38898 21508 38904
rect 21468 38554 21496 38898
rect 21456 38548 21508 38554
rect 21456 38490 21508 38496
rect 21468 38350 21496 38490
rect 21456 38344 21508 38350
rect 21456 38286 21508 38292
rect 21456 37800 21508 37806
rect 21456 37742 21508 37748
rect 21284 37318 21404 37346
rect 21180 36712 21232 36718
rect 21180 36654 21232 36660
rect 21192 36242 21220 36654
rect 21180 36236 21232 36242
rect 21180 36178 21232 36184
rect 21180 35760 21232 35766
rect 21180 35702 21232 35708
rect 20996 34196 21048 34202
rect 20996 34138 21048 34144
rect 21088 33856 21140 33862
rect 21088 33798 21140 33804
rect 21100 33658 21128 33798
rect 21088 33652 21140 33658
rect 21088 33594 21140 33600
rect 20720 33448 20772 33454
rect 20720 33390 20772 33396
rect 20628 33380 20680 33386
rect 20628 33322 20680 33328
rect 20640 32502 20668 33322
rect 20628 32496 20680 32502
rect 20628 32438 20680 32444
rect 20536 32428 20588 32434
rect 20536 32370 20588 32376
rect 20548 32026 20576 32370
rect 20536 32020 20588 32026
rect 20536 31962 20588 31968
rect 20640 31890 20668 32438
rect 20732 32434 20760 33390
rect 20904 33108 20956 33114
rect 20904 33050 20956 33056
rect 20812 32496 20864 32502
rect 20812 32438 20864 32444
rect 20720 32428 20772 32434
rect 20720 32370 20772 32376
rect 20732 32298 20760 32370
rect 20720 32292 20772 32298
rect 20720 32234 20772 32240
rect 20628 31884 20680 31890
rect 20628 31826 20680 31832
rect 20628 30796 20680 30802
rect 20628 30738 20680 30744
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 20536 30728 20588 30734
rect 20536 30670 20588 30676
rect 20456 30326 20484 30670
rect 20444 30320 20496 30326
rect 20444 30262 20496 30268
rect 20548 30258 20576 30670
rect 20640 30394 20668 30738
rect 20628 30388 20680 30394
rect 20628 30330 20680 30336
rect 20536 30252 20588 30258
rect 20536 30194 20588 30200
rect 20824 30122 20852 32438
rect 20916 32434 20944 33050
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 21192 31346 21220 35702
rect 21284 33114 21312 37318
rect 21468 37194 21496 37742
rect 21456 37188 21508 37194
rect 21456 37130 21508 37136
rect 21364 36780 21416 36786
rect 21364 36722 21416 36728
rect 21376 36038 21404 36722
rect 21468 36174 21496 37130
rect 21652 36650 21680 41074
rect 21928 41070 21956 41550
rect 22020 41274 22048 42570
rect 22468 42152 22520 42158
rect 22468 42094 22520 42100
rect 22480 41818 22508 42094
rect 22560 42016 22612 42022
rect 22560 41958 22612 41964
rect 22468 41812 22520 41818
rect 22468 41754 22520 41760
rect 22572 41614 22600 41958
rect 22560 41608 22612 41614
rect 22560 41550 22612 41556
rect 22376 41540 22428 41546
rect 22376 41482 22428 41488
rect 22928 41540 22980 41546
rect 22928 41482 22980 41488
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 21916 41064 21968 41070
rect 21916 41006 21968 41012
rect 22388 41002 22416 41482
rect 22560 41472 22612 41478
rect 22560 41414 22612 41420
rect 22376 40996 22428 41002
rect 22376 40938 22428 40944
rect 22572 40526 22600 41414
rect 22744 41064 22796 41070
rect 22744 41006 22796 41012
rect 22560 40520 22612 40526
rect 22560 40462 22612 40468
rect 22560 40384 22612 40390
rect 22560 40326 22612 40332
rect 22100 40044 22152 40050
rect 22100 39986 22152 39992
rect 22112 39846 22140 39986
rect 22572 39982 22600 40326
rect 22560 39976 22612 39982
rect 22560 39918 22612 39924
rect 22100 39840 22152 39846
rect 22100 39782 22152 39788
rect 22112 39438 22140 39782
rect 22192 39500 22244 39506
rect 22192 39442 22244 39448
rect 22100 39432 22152 39438
rect 22100 39374 22152 39380
rect 21824 39364 21876 39370
rect 21824 39306 21876 39312
rect 21836 38962 21864 39306
rect 22112 39030 22140 39374
rect 22100 39024 22152 39030
rect 22100 38966 22152 38972
rect 21824 38956 21876 38962
rect 21824 38898 21876 38904
rect 21916 38344 21968 38350
rect 22204 38332 22232 39442
rect 22652 39296 22704 39302
rect 22652 39238 22704 39244
rect 22468 38888 22520 38894
rect 22468 38830 22520 38836
rect 22480 38554 22508 38830
rect 22560 38752 22612 38758
rect 22560 38694 22612 38700
rect 22468 38548 22520 38554
rect 22468 38490 22520 38496
rect 22572 38350 22600 38694
rect 22664 38418 22692 39238
rect 22652 38412 22704 38418
rect 22652 38354 22704 38360
rect 21968 38321 22232 38332
rect 22560 38344 22612 38350
rect 21968 38312 22246 38321
rect 21968 38304 22190 38312
rect 21916 38286 21968 38292
rect 21928 37942 21956 38286
rect 22560 38286 22612 38292
rect 22190 38247 22246 38256
rect 21916 37936 21968 37942
rect 21916 37878 21968 37884
rect 22468 37460 22520 37466
rect 22468 37402 22520 37408
rect 21640 36644 21692 36650
rect 21640 36586 21692 36592
rect 21640 36236 21692 36242
rect 21640 36178 21692 36184
rect 21456 36168 21508 36174
rect 21456 36110 21508 36116
rect 21364 36032 21416 36038
rect 21364 35974 21416 35980
rect 21376 34950 21404 35974
rect 21364 34944 21416 34950
rect 21364 34886 21416 34892
rect 21376 33522 21404 34886
rect 21468 33930 21496 36110
rect 21548 35692 21600 35698
rect 21548 35634 21600 35640
rect 21456 33924 21508 33930
rect 21456 33866 21508 33872
rect 21364 33516 21416 33522
rect 21364 33458 21416 33464
rect 21272 33108 21324 33114
rect 21272 33050 21324 33056
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 21456 32836 21508 32842
rect 21456 32778 21508 32784
rect 21376 32502 21404 32778
rect 21364 32496 21416 32502
rect 21364 32438 21416 32444
rect 21468 32026 21496 32778
rect 21456 32020 21508 32026
rect 21456 31962 21508 31968
rect 21560 31958 21588 35634
rect 21652 35630 21680 36178
rect 21640 35624 21692 35630
rect 21640 35566 21692 35572
rect 22376 35624 22428 35630
rect 22376 35566 22428 35572
rect 22100 35488 22152 35494
rect 22100 35430 22152 35436
rect 22112 35154 22140 35430
rect 22100 35148 22152 35154
rect 22100 35090 22152 35096
rect 22192 35012 22244 35018
rect 22192 34954 22244 34960
rect 21916 34944 21968 34950
rect 21916 34886 21968 34892
rect 21928 33658 21956 34886
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 22020 34218 22048 34478
rect 22098 34232 22154 34241
rect 22020 34190 22098 34218
rect 22098 34167 22154 34176
rect 22112 33998 22140 34167
rect 22100 33992 22152 33998
rect 22100 33934 22152 33940
rect 21916 33652 21968 33658
rect 21916 33594 21968 33600
rect 21732 32768 21784 32774
rect 21732 32710 21784 32716
rect 21548 31952 21600 31958
rect 21548 31894 21600 31900
rect 21560 31482 21588 31894
rect 21548 31476 21600 31482
rect 21548 31418 21600 31424
rect 21640 31476 21692 31482
rect 21640 31418 21692 31424
rect 21180 31340 21232 31346
rect 21180 31282 21232 31288
rect 21548 30932 21600 30938
rect 21548 30874 21600 30880
rect 21088 30728 21140 30734
rect 21088 30670 21140 30676
rect 21100 30394 21128 30670
rect 21088 30388 21140 30394
rect 21088 30330 21140 30336
rect 20812 30116 20864 30122
rect 20812 30058 20864 30064
rect 20720 29640 20772 29646
rect 20718 29608 20720 29617
rect 20772 29608 20774 29617
rect 20718 29543 20774 29552
rect 20536 27464 20588 27470
rect 20536 27406 20588 27412
rect 20444 27396 20496 27402
rect 20444 27338 20496 27344
rect 20456 26858 20484 27338
rect 20548 27062 20576 27406
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 20536 27056 20588 27062
rect 20536 26998 20588 27004
rect 20444 26852 20496 26858
rect 20444 26794 20496 26800
rect 20456 26586 20484 26794
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20456 25974 20484 26522
rect 20640 26450 20668 27066
rect 20732 26926 20760 29543
rect 20994 29200 21050 29209
rect 20994 29135 20996 29144
rect 21048 29135 21050 29144
rect 20996 29106 21048 29112
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 20824 27441 20852 28494
rect 20810 27432 20866 27441
rect 20810 27367 20866 27376
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20812 26852 20864 26858
rect 20812 26794 20864 26800
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20536 26308 20588 26314
rect 20536 26250 20588 26256
rect 20444 25968 20496 25974
rect 20444 25910 20496 25916
rect 20548 25906 20576 26250
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20824 25430 20852 26794
rect 20812 25424 20864 25430
rect 20812 25366 20864 25372
rect 21100 25294 21128 30330
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 21180 30048 21232 30054
rect 21180 29990 21232 29996
rect 21192 29850 21220 29990
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 21284 28762 21312 30194
rect 21560 30190 21588 30874
rect 21652 30258 21680 31418
rect 21640 30252 21692 30258
rect 21640 30194 21692 30200
rect 21548 30184 21600 30190
rect 21548 30126 21600 30132
rect 21652 29889 21680 30194
rect 21638 29880 21694 29889
rect 21638 29815 21694 29824
rect 21364 29504 21416 29510
rect 21364 29446 21416 29452
rect 21376 29306 21404 29446
rect 21364 29300 21416 29306
rect 21364 29242 21416 29248
rect 21376 28762 21404 29242
rect 21456 28960 21508 28966
rect 21456 28902 21508 28908
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 21364 28756 21416 28762
rect 21364 28698 21416 28704
rect 21468 28490 21496 28902
rect 21456 28484 21508 28490
rect 21456 28426 21508 28432
rect 21548 28484 21600 28490
rect 21548 28426 21600 28432
rect 21180 26920 21232 26926
rect 21178 26888 21180 26897
rect 21232 26888 21234 26897
rect 21178 26823 21234 26832
rect 21560 26382 21588 28426
rect 21640 28076 21692 28082
rect 21640 28018 21692 28024
rect 21652 27538 21680 28018
rect 21744 27878 21772 32710
rect 21916 32564 21968 32570
rect 21916 32506 21968 32512
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 21836 31142 21864 32370
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 21824 30660 21876 30666
rect 21824 30602 21876 30608
rect 21836 30326 21864 30602
rect 21824 30320 21876 30326
rect 21824 30262 21876 30268
rect 21824 29844 21876 29850
rect 21824 29786 21876 29792
rect 21836 29510 21864 29786
rect 21824 29504 21876 29510
rect 21824 29446 21876 29452
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 21836 28762 21864 29106
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 21732 27872 21784 27878
rect 21732 27814 21784 27820
rect 21928 27554 21956 32506
rect 22008 32224 22060 32230
rect 22008 32166 22060 32172
rect 22020 31822 22048 32166
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22100 31748 22152 31754
rect 22100 31690 22152 31696
rect 22112 30938 22140 31690
rect 22204 31482 22232 34954
rect 22388 33862 22416 35566
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 22376 32496 22428 32502
rect 22376 32438 22428 32444
rect 22388 31890 22416 32438
rect 22376 31884 22428 31890
rect 22376 31826 22428 31832
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 22192 30864 22244 30870
rect 22192 30806 22244 30812
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 22020 30598 22048 30670
rect 22008 30592 22060 30598
rect 22008 30534 22060 30540
rect 22020 30258 22048 30534
rect 22204 30258 22232 30806
rect 22008 30252 22060 30258
rect 22192 30252 22244 30258
rect 22008 30194 22060 30200
rect 22112 30212 22192 30240
rect 22112 29510 22140 30212
rect 22192 30194 22244 30200
rect 22190 29880 22246 29889
rect 22296 29866 22324 31282
rect 22480 30666 22508 37402
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22664 36242 22692 36654
rect 22652 36236 22704 36242
rect 22652 36178 22704 36184
rect 22756 35834 22784 41006
rect 22836 38344 22888 38350
rect 22836 38286 22888 38292
rect 22848 36854 22876 38286
rect 22836 36848 22888 36854
rect 22836 36790 22888 36796
rect 22940 35834 22968 41482
rect 23020 39976 23072 39982
rect 23020 39918 23072 39924
rect 23032 38486 23060 39918
rect 23020 38480 23072 38486
rect 23020 38422 23072 38428
rect 23018 38312 23074 38321
rect 23018 38247 23020 38256
rect 23072 38247 23074 38256
rect 23020 38218 23072 38224
rect 23020 37800 23072 37806
rect 23020 37742 23072 37748
rect 23032 37466 23060 37742
rect 23020 37460 23072 37466
rect 23020 37402 23072 37408
rect 23020 37324 23072 37330
rect 23020 37266 23072 37272
rect 23032 37126 23060 37266
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 23032 36718 23060 37062
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 23020 36236 23072 36242
rect 23020 36178 23072 36184
rect 22744 35828 22796 35834
rect 22744 35770 22796 35776
rect 22928 35828 22980 35834
rect 22928 35770 22980 35776
rect 22560 35760 22612 35766
rect 23032 35714 23060 36178
rect 22560 35702 22612 35708
rect 22572 34746 22600 35702
rect 22940 35686 23060 35714
rect 22836 34944 22888 34950
rect 22836 34886 22888 34892
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 22848 34678 22876 34886
rect 22836 34672 22888 34678
rect 22836 34614 22888 34620
rect 22744 33108 22796 33114
rect 22744 33050 22796 33056
rect 22756 32434 22784 33050
rect 22744 32428 22796 32434
rect 22744 32370 22796 32376
rect 22560 32224 22612 32230
rect 22560 32166 22612 32172
rect 22572 32026 22600 32166
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22744 31884 22796 31890
rect 22744 31826 22796 31832
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22468 30660 22520 30666
rect 22468 30602 22520 30608
rect 22376 30592 22428 30598
rect 22374 30560 22376 30569
rect 22428 30560 22430 30569
rect 22374 30495 22430 30504
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22480 30054 22508 30194
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 22466 29880 22522 29889
rect 22296 29838 22360 29866
rect 22190 29815 22246 29824
rect 22100 29504 22152 29510
rect 22100 29446 22152 29452
rect 22098 29200 22154 29209
rect 22008 29164 22060 29170
rect 22098 29135 22100 29144
rect 22008 29106 22060 29112
rect 22152 29135 22154 29144
rect 22100 29106 22152 29112
rect 22020 28694 22048 29106
rect 22008 28688 22060 28694
rect 22008 28630 22060 28636
rect 22204 28626 22232 29815
rect 22332 29764 22360 29838
rect 22466 29815 22468 29824
rect 22520 29815 22522 29824
rect 22468 29786 22520 29792
rect 22296 29736 22360 29764
rect 22192 28620 22244 28626
rect 22192 28562 22244 28568
rect 22204 28490 22232 28562
rect 22192 28484 22244 28490
rect 22192 28426 22244 28432
rect 22008 27872 22060 27878
rect 22008 27814 22060 27820
rect 22020 27606 22048 27814
rect 21640 27532 21692 27538
rect 21640 27474 21692 27480
rect 21744 27526 21956 27554
rect 22008 27600 22060 27606
rect 22008 27542 22060 27548
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 21456 26240 21508 26246
rect 21456 26182 21508 26188
rect 21180 25968 21232 25974
rect 21180 25910 21232 25916
rect 21192 25498 21220 25910
rect 21180 25492 21232 25498
rect 21180 25434 21232 25440
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 20444 25152 20496 25158
rect 20444 25094 20496 25100
rect 20456 24138 20484 25094
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20444 24132 20496 24138
rect 20444 24074 20496 24080
rect 20442 23896 20498 23905
rect 20442 23831 20444 23840
rect 20496 23831 20498 23840
rect 20444 23802 20496 23808
rect 20732 22710 20760 24346
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20536 22432 20588 22438
rect 20536 22374 20588 22380
rect 20456 21962 20484 22374
rect 20444 21956 20496 21962
rect 20444 21898 20496 21904
rect 20548 21622 20576 22374
rect 20640 22234 20668 22578
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20640 21894 20668 22170
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20536 21616 20588 21622
rect 20536 21558 20588 21564
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 19786 20484 21286
rect 20548 20058 20576 21558
rect 20628 21412 20680 21418
rect 20628 21354 20680 21360
rect 20640 21078 20668 21354
rect 20628 21072 20680 21078
rect 20628 21014 20680 21020
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20640 19922 20668 21014
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20732 19786 20760 20402
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20732 19446 20760 19722
rect 20720 19440 20772 19446
rect 20772 19388 20852 19394
rect 20720 19382 20852 19388
rect 20732 19366 20852 19382
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20732 18970 20760 19246
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20824 18426 20852 19366
rect 20916 19310 20944 25230
rect 21284 24886 21312 26182
rect 21468 25974 21496 26182
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 21364 25900 21416 25906
rect 21364 25842 21416 25848
rect 21376 24954 21404 25842
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21652 25294 21680 25638
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21364 24948 21416 24954
rect 21364 24890 21416 24896
rect 21272 24880 21324 24886
rect 21272 24822 21324 24828
rect 21744 23322 21772 27526
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 21836 27130 21864 27406
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 21836 26042 21864 27066
rect 22112 26858 22140 27406
rect 22100 26852 22152 26858
rect 22100 26794 22152 26800
rect 22296 26382 22324 29736
rect 22468 29232 22520 29238
rect 22468 29174 22520 29180
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22388 28558 22416 28902
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22374 27704 22430 27713
rect 22374 27639 22376 27648
rect 22428 27639 22430 27648
rect 22376 27610 22428 27616
rect 22480 26790 22508 29174
rect 22560 29096 22612 29102
rect 22560 29038 22612 29044
rect 22572 28762 22600 29038
rect 22560 28756 22612 28762
rect 22560 28698 22612 28704
rect 22560 27396 22612 27402
rect 22560 27338 22612 27344
rect 22572 26926 22600 27338
rect 22560 26920 22612 26926
rect 22560 26862 22612 26868
rect 22468 26784 22520 26790
rect 22468 26726 22520 26732
rect 22284 26376 22336 26382
rect 22336 26336 22416 26364
rect 22284 26318 22336 26324
rect 22100 26240 22152 26246
rect 22100 26182 22152 26188
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 22112 25974 22140 26182
rect 22100 25968 22152 25974
rect 22100 25910 22152 25916
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22020 25702 22048 25842
rect 22204 25786 22232 26182
rect 22112 25758 22232 25786
rect 22284 25764 22336 25770
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 22112 25498 22140 25758
rect 22284 25706 22336 25712
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 22112 25294 22140 25434
rect 22296 25294 22324 25706
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22100 25152 22152 25158
rect 22098 25120 22100 25129
rect 22284 25152 22336 25158
rect 22152 25120 22154 25129
rect 22284 25094 22336 25100
rect 22098 25055 22154 25064
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21836 24274 21864 24550
rect 22204 24410 22232 24890
rect 22296 24818 22324 25094
rect 22388 24954 22416 26336
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22480 24857 22508 26726
rect 22572 26586 22600 26862
rect 22560 26580 22612 26586
rect 22560 26522 22612 26528
rect 22560 26240 22612 26246
rect 22560 26182 22612 26188
rect 22572 25906 22600 26182
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22466 24848 22522 24857
rect 22284 24812 22336 24818
rect 22466 24783 22522 24792
rect 22284 24754 22336 24760
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 21824 24268 21876 24274
rect 21824 24210 21876 24216
rect 21916 24132 21968 24138
rect 21916 24074 21968 24080
rect 22468 24132 22520 24138
rect 22468 24074 22520 24080
rect 21928 23866 21956 24074
rect 22480 23866 22508 24074
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 22560 23792 22612 23798
rect 22560 23734 22612 23740
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21088 22500 21140 22506
rect 21088 22442 21140 22448
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21008 19530 21036 21830
rect 21100 21554 21128 22442
rect 21468 22094 21496 22578
rect 21824 22568 21876 22574
rect 21824 22510 21876 22516
rect 21732 22432 21784 22438
rect 21732 22374 21784 22380
rect 21376 22066 21496 22094
rect 21376 21690 21404 22066
rect 21744 22030 21772 22374
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21100 19718 21128 20334
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21008 19502 21128 19530
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20916 18766 20944 19246
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20824 17270 20852 18362
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20916 17610 20944 18090
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20812 17264 20864 17270
rect 20864 17224 20944 17252
rect 20812 17206 20864 17212
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20824 16794 20852 17070
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20180 14906 20208 15982
rect 20272 15910 20300 16526
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20364 15094 20392 15642
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20456 15094 20484 15302
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20444 14952 20496 14958
rect 20180 14878 20300 14906
rect 20548 14940 20576 15370
rect 20640 15094 20668 16390
rect 20732 15910 20760 16526
rect 20916 16250 20944 17224
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20812 16176 20864 16182
rect 20812 16118 20864 16124
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20496 14912 20576 14940
rect 20444 14894 20496 14900
rect 20272 14550 20300 14878
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 20272 14346 20300 14486
rect 20548 14482 20576 14912
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 19996 13110 20116 13138
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19800 12164 19852 12170
rect 19800 12106 19852 12112
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19536 11218 19564 12038
rect 19996 11898 20024 13110
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20088 12102 20116 12786
rect 20180 12374 20208 12854
rect 20168 12368 20220 12374
rect 20168 12310 20220 12316
rect 20272 12238 20300 14282
rect 20548 14074 20576 14418
rect 20732 14414 20760 15846
rect 20824 15706 20852 16118
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20916 15706 20944 15914
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20916 15162 20944 15642
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 21008 15026 21036 15302
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21100 14906 21128 19502
rect 21192 17082 21220 21422
rect 21468 20942 21496 21966
rect 21836 21894 21864 22510
rect 21824 21888 21876 21894
rect 21824 21830 21876 21836
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21836 20874 21864 21286
rect 21824 20868 21876 20874
rect 21824 20810 21876 20816
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21192 17054 21312 17082
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21192 16250 21220 16458
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21284 15450 21312 17054
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21376 15978 21404 16934
rect 21468 16590 21496 18566
rect 21836 17202 21864 19654
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21376 15570 21404 15914
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21284 15422 21404 15450
rect 21008 14878 21128 14906
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 21008 12434 21036 14878
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 21100 13394 21128 14214
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20732 12406 21036 12434
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19628 11354 19656 11630
rect 19996 11558 20024 11834
rect 20088 11626 20116 12038
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19524 11212 19576 11218
rect 19892 11212 19944 11218
rect 19524 11154 19576 11160
rect 19812 11172 19892 11200
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19444 10810 19472 11018
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19812 9586 19840 11172
rect 19892 11154 19944 11160
rect 20180 11082 20208 12106
rect 20732 11830 20760 12406
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 20548 11218 20576 11630
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20180 10674 20208 11018
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20088 9654 20116 10406
rect 20180 9994 20208 10610
rect 21100 10130 21128 10950
rect 21284 10538 21312 14350
rect 21376 11762 21404 15422
rect 21640 14884 21692 14890
rect 21640 14826 21692 14832
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14346 21496 14758
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21652 13870 21680 14826
rect 21744 14822 21772 16526
rect 21836 16114 21864 17138
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21822 15600 21878 15609
rect 21822 15535 21878 15544
rect 21836 15502 21864 15535
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21744 14550 21772 14758
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21652 13462 21680 13806
rect 21928 13530 21956 23258
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22480 22710 22508 22918
rect 22572 22778 22600 23734
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22468 22704 22520 22710
rect 22468 22646 22520 22652
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22296 20602 22324 21490
rect 22388 21434 22416 22510
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 22572 21570 22600 22374
rect 22664 21690 22692 31078
rect 22756 29238 22784 31826
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 22742 28520 22798 28529
rect 22742 28455 22798 28464
rect 22756 24682 22784 28455
rect 22836 27396 22888 27402
rect 22836 27338 22888 27344
rect 22848 27305 22876 27338
rect 22834 27296 22890 27305
rect 22834 27231 22890 27240
rect 22940 26790 22968 35686
rect 23020 35148 23072 35154
rect 23020 35090 23072 35096
rect 23032 34406 23060 35090
rect 23020 34400 23072 34406
rect 23020 34342 23072 34348
rect 23124 33114 23152 43250
rect 23572 42832 23624 42838
rect 23572 42774 23624 42780
rect 23296 42628 23348 42634
rect 23296 42570 23348 42576
rect 23308 41614 23336 42570
rect 23480 42560 23532 42566
rect 23480 42502 23532 42508
rect 23492 41682 23520 42502
rect 23584 41750 23612 42774
rect 23572 41744 23624 41750
rect 23624 41692 23704 41698
rect 23572 41686 23704 41692
rect 23480 41676 23532 41682
rect 23584 41670 23704 41686
rect 23480 41618 23532 41624
rect 23296 41608 23348 41614
rect 23296 41550 23348 41556
rect 23572 41540 23624 41546
rect 23572 41482 23624 41488
rect 23480 41472 23532 41478
rect 23480 41414 23532 41420
rect 23492 41138 23520 41414
rect 23584 41274 23612 41482
rect 23572 41268 23624 41274
rect 23572 41210 23624 41216
rect 23480 41132 23532 41138
rect 23480 41074 23532 41080
rect 23572 41064 23624 41070
rect 23386 41032 23442 41041
rect 23676 41052 23704 41670
rect 23624 41024 23704 41052
rect 23572 41006 23624 41012
rect 23386 40967 23442 40976
rect 23400 40118 23428 40967
rect 23388 40112 23440 40118
rect 23388 40054 23440 40060
rect 23480 39092 23532 39098
rect 23480 39034 23532 39040
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 23388 37120 23440 37126
rect 23388 37062 23440 37068
rect 23216 36922 23244 37062
rect 23204 36916 23256 36922
rect 23204 36858 23256 36864
rect 23400 36242 23428 37062
rect 23492 36854 23520 39034
rect 23676 37670 23704 41024
rect 23664 37664 23716 37670
rect 23664 37606 23716 37612
rect 23664 37120 23716 37126
rect 23664 37062 23716 37068
rect 23676 36854 23704 37062
rect 23480 36848 23532 36854
rect 23480 36790 23532 36796
rect 23664 36848 23716 36854
rect 23664 36790 23716 36796
rect 23388 36236 23440 36242
rect 23388 36178 23440 36184
rect 23492 36106 23520 36790
rect 23480 36100 23532 36106
rect 23480 36042 23532 36048
rect 23492 35766 23520 36042
rect 23480 35760 23532 35766
rect 23480 35702 23532 35708
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23204 34944 23256 34950
rect 23256 34904 23336 34932
rect 23204 34886 23256 34892
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 23216 33522 23244 33798
rect 23204 33516 23256 33522
rect 23204 33458 23256 33464
rect 23112 33108 23164 33114
rect 23112 33050 23164 33056
rect 23020 33040 23072 33046
rect 23020 32982 23072 32988
rect 23032 32502 23060 32982
rect 23020 32496 23072 32502
rect 23020 32438 23072 32444
rect 23032 30394 23060 32438
rect 23308 31482 23336 34904
rect 23400 34762 23428 35090
rect 23400 34746 23520 34762
rect 23400 34740 23532 34746
rect 23400 34734 23480 34740
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 23020 30388 23072 30394
rect 23020 30330 23072 30336
rect 23032 29646 23060 30330
rect 23308 30190 23336 31418
rect 23400 31414 23428 34734
rect 23480 34682 23532 34688
rect 23768 34626 23796 43250
rect 26240 43240 26292 43246
rect 26240 43182 26292 43188
rect 33876 43240 33928 43246
rect 33876 43182 33928 43188
rect 25872 43104 25924 43110
rect 25872 43046 25924 43052
rect 25884 42702 25912 43046
rect 23940 42696 23992 42702
rect 23940 42638 23992 42644
rect 24676 42696 24728 42702
rect 24676 42638 24728 42644
rect 25872 42696 25924 42702
rect 25872 42638 25924 42644
rect 23952 42294 23980 42638
rect 24584 42560 24636 42566
rect 24584 42502 24636 42508
rect 24596 42294 24624 42502
rect 23940 42288 23992 42294
rect 23940 42230 23992 42236
rect 24584 42288 24636 42294
rect 24584 42230 24636 42236
rect 23952 41818 23980 42230
rect 24308 42220 24360 42226
rect 24308 42162 24360 42168
rect 23940 41812 23992 41818
rect 23940 41754 23992 41760
rect 23848 41676 23900 41682
rect 23848 41618 23900 41624
rect 23860 41206 23888 41618
rect 23848 41200 23900 41206
rect 23848 41142 23900 41148
rect 23952 39030 23980 41754
rect 24320 41682 24348 42162
rect 24688 42022 24716 42638
rect 25872 42560 25924 42566
rect 25872 42502 25924 42508
rect 26056 42560 26108 42566
rect 26056 42502 26108 42508
rect 25688 42220 25740 42226
rect 25688 42162 25740 42168
rect 24676 42016 24728 42022
rect 24676 41958 24728 41964
rect 24584 41744 24636 41750
rect 24584 41686 24636 41692
rect 24308 41676 24360 41682
rect 24308 41618 24360 41624
rect 24320 40050 24348 41618
rect 24400 41608 24452 41614
rect 24400 41550 24452 41556
rect 24412 41002 24440 41550
rect 24400 40996 24452 41002
rect 24400 40938 24452 40944
rect 24596 40526 24624 41686
rect 24688 41614 24716 41958
rect 25700 41818 25728 42162
rect 25688 41812 25740 41818
rect 25688 41754 25740 41760
rect 24676 41608 24728 41614
rect 24676 41550 24728 41556
rect 25700 41546 25728 41754
rect 25688 41540 25740 41546
rect 25688 41482 25740 41488
rect 24768 41472 24820 41478
rect 24768 41414 24820 41420
rect 24780 41138 24808 41414
rect 24768 41132 24820 41138
rect 24768 41074 24820 41080
rect 24860 40588 24912 40594
rect 24860 40530 24912 40536
rect 24584 40520 24636 40526
rect 24584 40462 24636 40468
rect 24400 40180 24452 40186
rect 24400 40122 24452 40128
rect 24308 40044 24360 40050
rect 24308 39986 24360 39992
rect 24320 39438 24348 39986
rect 24308 39432 24360 39438
rect 24308 39374 24360 39380
rect 24320 39098 24348 39374
rect 24308 39092 24360 39098
rect 24308 39034 24360 39040
rect 23940 39024 23992 39030
rect 23940 38966 23992 38972
rect 23952 36922 23980 38966
rect 24124 38820 24176 38826
rect 24124 38762 24176 38768
rect 24032 38752 24084 38758
rect 24032 38694 24084 38700
rect 24044 38418 24072 38694
rect 24032 38412 24084 38418
rect 24032 38354 24084 38360
rect 24136 38298 24164 38762
rect 24412 38758 24440 40122
rect 24596 40050 24624 40462
rect 24872 40050 24900 40530
rect 25136 40520 25188 40526
rect 25136 40462 25188 40468
rect 25412 40520 25464 40526
rect 25412 40462 25464 40468
rect 24584 40044 24636 40050
rect 24584 39986 24636 39992
rect 24860 40044 24912 40050
rect 25148 40032 25176 40462
rect 25228 40044 25280 40050
rect 25148 40004 25228 40032
rect 24860 39986 24912 39992
rect 25228 39986 25280 39992
rect 24768 39840 24820 39846
rect 24768 39782 24820 39788
rect 24584 39568 24636 39574
rect 24584 39510 24636 39516
rect 24400 38752 24452 38758
rect 24400 38694 24452 38700
rect 24412 38350 24440 38694
rect 24596 38350 24624 39510
rect 24780 39438 24808 39782
rect 25240 39438 25268 39986
rect 25424 39930 25452 40462
rect 25332 39914 25452 39930
rect 25320 39908 25452 39914
rect 25372 39902 25452 39908
rect 25320 39850 25372 39856
rect 25332 39438 25360 39850
rect 24768 39432 24820 39438
rect 24768 39374 24820 39380
rect 25228 39432 25280 39438
rect 25228 39374 25280 39380
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 24860 38956 24912 38962
rect 24860 38898 24912 38904
rect 25044 38956 25096 38962
rect 25044 38898 25096 38904
rect 24872 38554 24900 38898
rect 24860 38548 24912 38554
rect 24860 38490 24912 38496
rect 25056 38434 25084 38898
rect 25240 38826 25268 39374
rect 25332 39098 25360 39374
rect 25596 39296 25648 39302
rect 25596 39238 25648 39244
rect 25320 39092 25372 39098
rect 25320 39034 25372 39040
rect 25608 39030 25636 39238
rect 25596 39024 25648 39030
rect 25596 38966 25648 38972
rect 25320 38956 25372 38962
rect 25320 38898 25372 38904
rect 25412 38956 25464 38962
rect 25412 38898 25464 38904
rect 25228 38820 25280 38826
rect 25228 38762 25280 38768
rect 25332 38554 25360 38898
rect 25320 38548 25372 38554
rect 25320 38490 25372 38496
rect 25424 38434 25452 38898
rect 25056 38406 25452 38434
rect 25608 38418 25636 38966
rect 24044 38270 24164 38298
rect 24400 38344 24452 38350
rect 24400 38286 24452 38292
rect 24584 38344 24636 38350
rect 24584 38286 24636 38292
rect 25044 38344 25096 38350
rect 25044 38286 25096 38292
rect 23940 36916 23992 36922
rect 23940 36858 23992 36864
rect 23952 36038 23980 36858
rect 23940 36032 23992 36038
rect 23940 35974 23992 35980
rect 23492 34598 23796 34626
rect 23492 32026 23520 34598
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 23676 33998 23704 34478
rect 23756 34400 23808 34406
rect 23756 34342 23808 34348
rect 23664 33992 23716 33998
rect 23664 33934 23716 33940
rect 23768 33522 23796 34342
rect 23860 33658 23888 34478
rect 23940 33924 23992 33930
rect 23940 33866 23992 33872
rect 23952 33658 23980 33866
rect 23848 33652 23900 33658
rect 23848 33594 23900 33600
rect 23940 33652 23992 33658
rect 23940 33594 23992 33600
rect 23756 33516 23808 33522
rect 23756 33458 23808 33464
rect 24044 33402 24072 38270
rect 24596 38214 24624 38286
rect 24584 38208 24636 38214
rect 24584 38150 24636 38156
rect 24768 37664 24820 37670
rect 24768 37606 24820 37612
rect 24780 37330 24808 37606
rect 24768 37324 24820 37330
rect 24768 37266 24820 37272
rect 24860 37324 24912 37330
rect 24860 37266 24912 37272
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 24124 34604 24176 34610
rect 24124 34546 24176 34552
rect 23584 33374 24072 33402
rect 23480 32020 23532 32026
rect 23480 31962 23532 31968
rect 23492 31822 23520 31962
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23388 31408 23440 31414
rect 23388 31350 23440 31356
rect 23584 30734 23612 33374
rect 23664 32768 23716 32774
rect 23664 32710 23716 32716
rect 23676 32366 23704 32710
rect 24032 32496 24084 32502
rect 24032 32438 24084 32444
rect 23664 32360 23716 32366
rect 23664 32302 23716 32308
rect 23676 31822 23704 32302
rect 24044 32026 24072 32438
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 23676 30870 23704 31758
rect 24032 31748 24084 31754
rect 24032 31690 24084 31696
rect 24044 31142 24072 31690
rect 24136 31346 24164 34546
rect 24412 33998 24440 36110
rect 24676 35624 24728 35630
rect 24676 35566 24728 35572
rect 24688 35290 24716 35566
rect 24676 35284 24728 35290
rect 24676 35226 24728 35232
rect 24780 35154 24808 37266
rect 24768 35148 24820 35154
rect 24768 35090 24820 35096
rect 24872 34746 24900 37266
rect 25056 37262 25084 38286
rect 25044 37256 25096 37262
rect 25044 37198 25096 37204
rect 25056 36922 25084 37198
rect 25044 36916 25096 36922
rect 25044 36858 25096 36864
rect 25320 36576 25372 36582
rect 25320 36518 25372 36524
rect 25332 36106 25360 36518
rect 25320 36100 25372 36106
rect 25320 36042 25372 36048
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 25148 35766 25176 35974
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 25424 35630 25452 38406
rect 25596 38412 25648 38418
rect 25596 38354 25648 38360
rect 25688 38276 25740 38282
rect 25688 38218 25740 38224
rect 25596 38208 25648 38214
rect 25596 38150 25648 38156
rect 25504 37868 25556 37874
rect 25504 37810 25556 37816
rect 25516 36378 25544 37810
rect 25608 36922 25636 38150
rect 25700 37262 25728 38218
rect 25688 37256 25740 37262
rect 25688 37198 25740 37204
rect 25596 36916 25648 36922
rect 25596 36858 25648 36864
rect 25780 36644 25832 36650
rect 25780 36586 25832 36592
rect 25504 36372 25556 36378
rect 25504 36314 25556 36320
rect 25792 36106 25820 36586
rect 25780 36100 25832 36106
rect 25780 36042 25832 36048
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 25412 35488 25464 35494
rect 25412 35430 25464 35436
rect 25320 34944 25372 34950
rect 25320 34886 25372 34892
rect 25332 34746 25360 34886
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 25320 34740 25372 34746
rect 25320 34682 25372 34688
rect 25424 34542 25452 35430
rect 25596 34672 25648 34678
rect 25596 34614 25648 34620
rect 25136 34536 25188 34542
rect 25136 34478 25188 34484
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24412 32978 24440 33934
rect 24768 33924 24820 33930
rect 24768 33866 24820 33872
rect 24780 33658 24808 33866
rect 25148 33862 25176 34478
rect 25320 34400 25372 34406
rect 25320 34342 25372 34348
rect 25136 33856 25188 33862
rect 25136 33798 25188 33804
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24400 32972 24452 32978
rect 24400 32914 24452 32920
rect 24308 32428 24360 32434
rect 24412 32416 24440 32914
rect 25148 32910 25176 33798
rect 25332 33454 25360 34342
rect 25412 33516 25464 33522
rect 25412 33458 25464 33464
rect 25228 33448 25280 33454
rect 25228 33390 25280 33396
rect 25320 33448 25372 33454
rect 25320 33390 25372 33396
rect 25240 33114 25268 33390
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 25136 32904 25188 32910
rect 25136 32846 25188 32852
rect 24360 32388 24440 32416
rect 24584 32428 24636 32434
rect 24308 32370 24360 32376
rect 24584 32370 24636 32376
rect 24124 31340 24176 31346
rect 24124 31282 24176 31288
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 23664 30864 23716 30870
rect 23664 30806 23716 30812
rect 23388 30728 23440 30734
rect 23572 30728 23624 30734
rect 23440 30688 23520 30716
rect 23388 30670 23440 30676
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 23204 30048 23256 30054
rect 23204 29990 23256 29996
rect 23216 29646 23244 29990
rect 23020 29640 23072 29646
rect 23020 29582 23072 29588
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23216 29345 23244 29582
rect 23202 29336 23258 29345
rect 23202 29271 23258 29280
rect 23308 29170 23336 30126
rect 23492 29646 23520 30688
rect 23624 30676 23704 30682
rect 23572 30670 23704 30676
rect 23584 30654 23704 30670
rect 23676 29646 23704 30654
rect 23848 29776 23900 29782
rect 23848 29718 23900 29724
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23492 29481 23520 29582
rect 23478 29472 23534 29481
rect 23478 29407 23534 29416
rect 23388 29232 23440 29238
rect 23388 29174 23440 29180
rect 23572 29232 23624 29238
rect 23572 29174 23624 29180
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 23020 29096 23072 29102
rect 23020 29038 23072 29044
rect 23032 28558 23060 29038
rect 23124 28762 23152 29106
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23112 28756 23164 28762
rect 23112 28698 23164 28704
rect 23124 28558 23152 28698
rect 23308 28558 23336 28902
rect 23400 28558 23428 29174
rect 23480 28688 23532 28694
rect 23480 28630 23532 28636
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23112 27668 23164 27674
rect 23112 27610 23164 27616
rect 23018 27568 23074 27577
rect 23018 27503 23020 27512
rect 23072 27503 23074 27512
rect 23020 27474 23072 27480
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23032 27130 23060 27270
rect 23020 27124 23072 27130
rect 23020 27066 23072 27072
rect 23124 26926 23152 27610
rect 23492 27112 23520 28630
rect 23584 28082 23612 29174
rect 23664 29028 23716 29034
rect 23664 28970 23716 28976
rect 23676 28762 23704 28970
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23664 28212 23716 28218
rect 23664 28154 23716 28160
rect 23572 28076 23624 28082
rect 23572 28018 23624 28024
rect 23676 27946 23704 28154
rect 23768 28082 23796 29582
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23664 27940 23716 27946
rect 23664 27882 23716 27888
rect 23400 27084 23520 27112
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 22928 26784 22980 26790
rect 22928 26726 22980 26732
rect 23112 26784 23164 26790
rect 23112 26726 23164 26732
rect 23124 26450 23152 26726
rect 23400 26518 23428 27084
rect 23768 27033 23796 28018
rect 23860 27538 23888 29718
rect 23938 29472 23994 29481
rect 23938 29407 23994 29416
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 23754 27024 23810 27033
rect 23480 26988 23532 26994
rect 23754 26959 23810 26968
rect 23480 26930 23532 26936
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 23112 26444 23164 26450
rect 23112 26386 23164 26392
rect 23400 26382 23428 26454
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 23020 25696 23072 25702
rect 23020 25638 23072 25644
rect 23032 25362 23060 25638
rect 23020 25356 23072 25362
rect 23020 25298 23072 25304
rect 23308 25294 23336 25706
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23400 25226 23428 25434
rect 23388 25220 23440 25226
rect 23388 25162 23440 25168
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 22744 24676 22796 24682
rect 22744 24618 22796 24624
rect 22756 23730 22784 24618
rect 23032 23866 23060 25094
rect 23400 24886 23428 25162
rect 23388 24880 23440 24886
rect 23388 24822 23440 24828
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 23020 23860 23072 23866
rect 23020 23802 23072 23808
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 23124 23474 23152 24754
rect 23492 24274 23520 26930
rect 23848 26512 23900 26518
rect 23848 26454 23900 26460
rect 23572 26444 23624 26450
rect 23572 26386 23624 26392
rect 23584 26330 23612 26386
rect 23756 26376 23808 26382
rect 23584 26302 23704 26330
rect 23756 26318 23808 26324
rect 23572 26240 23624 26246
rect 23572 26182 23624 26188
rect 23584 25362 23612 26182
rect 23676 25838 23704 26302
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23768 25702 23796 26318
rect 23860 25906 23888 26454
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23756 25696 23808 25702
rect 23756 25638 23808 25644
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 23952 25294 23980 29407
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23940 25288 23992 25294
rect 23940 25230 23992 25236
rect 23572 25220 23624 25226
rect 23572 25162 23624 25168
rect 23584 25129 23612 25162
rect 23570 25120 23626 25129
rect 23570 25055 23626 25064
rect 23480 24268 23532 24274
rect 23480 24210 23532 24216
rect 23032 23446 23152 23474
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22848 21894 22876 23054
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22572 21542 22692 21570
rect 22388 21418 22508 21434
rect 22388 21412 22520 21418
rect 22388 21406 22468 21412
rect 22468 21354 22520 21360
rect 22480 20942 22508 21354
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22480 20398 22508 20878
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 22020 19922 22048 20198
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22388 19174 22416 20334
rect 22480 19786 22508 20334
rect 22468 19780 22520 19786
rect 22468 19722 22520 19728
rect 22480 19514 22508 19722
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22192 18216 22244 18222
rect 22192 18158 22244 18164
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 22020 17202 22048 17750
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 22020 16114 22048 17138
rect 22100 17060 22152 17066
rect 22100 17002 22152 17008
rect 22112 16658 22140 17002
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22204 16454 22232 18158
rect 22480 17678 22508 19450
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22480 17338 22508 17614
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 16590 22600 16934
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22112 15910 22140 16390
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22112 15026 22140 15846
rect 22204 15638 22232 15982
rect 22192 15632 22244 15638
rect 22468 15632 22520 15638
rect 22192 15574 22244 15580
rect 22466 15600 22468 15609
rect 22520 15600 22522 15609
rect 22466 15535 22522 15544
rect 22284 15496 22336 15502
rect 22468 15496 22520 15502
rect 22284 15438 22336 15444
rect 22388 15456 22468 15484
rect 22296 15366 22324 15438
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22204 14958 22232 15302
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 22112 13938 22140 14282
rect 22296 14074 22324 14962
rect 22388 14618 22416 15456
rect 22468 15438 22520 15444
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22388 13870 22416 14554
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19536 9110 19564 9522
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 18380 8996 18460 9024
rect 18328 8978 18380 8984
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18432 8430 18460 8996
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11900 7002 11928 7278
rect 14568 7274 14596 7686
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 18064 6914 18092 7686
rect 17972 6886 18092 6914
rect 17972 6322 18000 6886
rect 18432 6866 18460 8366
rect 19076 7954 19104 8774
rect 19352 8294 19380 8978
rect 19536 8974 19564 9046
rect 19720 9042 19748 9522
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7546 18736 7754
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 19352 7410 19380 8230
rect 19628 8090 19656 8366
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19720 7954 19748 8978
rect 20180 8974 20208 9930
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20364 8974 20392 9522
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19812 8090 19840 8842
rect 19996 8430 20024 8842
rect 20180 8566 20208 8910
rect 20364 8634 20392 8910
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20168 8560 20220 8566
rect 20168 8502 20220 8508
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19720 7562 19748 7890
rect 19812 7886 19840 8026
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19628 7534 19748 7562
rect 19628 7478 19656 7534
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18432 6322 18460 6802
rect 18708 6390 18736 7142
rect 19628 7002 19656 7414
rect 19996 7342 20024 8366
rect 20364 8022 20392 8570
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20180 7546 20208 7754
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20364 7478 20392 7822
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 20180 6458 20208 7278
rect 20548 7002 20576 7686
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 20824 6390 20852 7210
rect 21192 6730 21220 9930
rect 21376 9518 21404 10066
rect 21468 9586 21496 12242
rect 22204 12170 22232 12378
rect 22388 12238 22416 13330
rect 22468 13252 22520 13258
rect 22468 13194 22520 13200
rect 22480 12986 22508 13194
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22664 12306 22692 21542
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22756 18970 22784 19246
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22756 17066 22784 17546
rect 22744 17060 22796 17066
rect 22744 17002 22796 17008
rect 22848 16946 22876 21830
rect 22756 16918 22876 16946
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 22296 11694 22324 12106
rect 22388 11898 22416 12174
rect 22756 12170 22784 16918
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22848 15094 22876 16458
rect 22940 15910 22968 16526
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22836 15088 22888 15094
rect 22836 15030 22888 15036
rect 22836 14340 22888 14346
rect 22836 14282 22888 14288
rect 22848 13870 22876 14282
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22848 13258 22876 13806
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 22940 12986 22968 13874
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 23032 12434 23060 23446
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23112 22636 23164 22642
rect 23112 22578 23164 22584
rect 23124 22234 23152 22578
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23216 21622 23244 21966
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 23216 21146 23244 21422
rect 23204 21140 23256 21146
rect 23204 21082 23256 21088
rect 23308 21026 23336 21830
rect 23216 20998 23336 21026
rect 23216 18834 23244 20998
rect 23400 19496 23428 22918
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23492 20534 23520 20742
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23308 19468 23428 19496
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 23124 13938 23152 14758
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23204 12436 23256 12442
rect 23032 12406 23152 12434
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22388 11762 22416 11834
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22480 11286 22508 12038
rect 22940 11830 22968 12242
rect 22928 11824 22980 11830
rect 22928 11766 22980 11772
rect 22652 11688 22704 11694
rect 22652 11630 22704 11636
rect 22664 11354 22692 11630
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22468 11280 22520 11286
rect 22468 11222 22520 11228
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22388 10810 22416 11086
rect 22836 11076 22888 11082
rect 22888 11036 22968 11064
rect 22836 11018 22888 11024
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22204 10266 22232 10542
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22008 9648 22060 9654
rect 22008 9590 22060 9596
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21652 9042 21680 9318
rect 21744 9178 21772 9454
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 22020 8974 22048 9590
rect 22296 9450 22324 9998
rect 22284 9444 22336 9450
rect 22284 9386 22336 9392
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22112 8838 22140 9318
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22296 8430 22324 8910
rect 22388 8634 22416 9114
rect 22664 9110 22692 9998
rect 22848 9926 22876 9998
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22756 9042 22784 9114
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22480 8634 22508 8842
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22756 8430 22784 8978
rect 22848 8634 22876 9862
rect 22940 9110 22968 11036
rect 23020 10600 23072 10606
rect 23020 10542 23072 10548
rect 22928 9104 22980 9110
rect 22928 9046 22980 9052
rect 23032 8906 23060 10542
rect 23020 8900 23072 8906
rect 23020 8842 23072 8848
rect 23124 8786 23152 12406
rect 23204 12378 23256 12384
rect 23216 11218 23244 12378
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 23308 11150 23336 19468
rect 23388 18760 23440 18766
rect 23492 18748 23520 19654
rect 23584 19446 23612 19654
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23440 18720 23520 18748
rect 23388 18702 23440 18708
rect 23676 18170 23704 25230
rect 23756 22568 23808 22574
rect 23756 22510 23808 22516
rect 23768 22098 23796 22510
rect 24044 22166 24072 31078
rect 24136 29730 24164 31282
rect 24216 31272 24268 31278
rect 24214 31240 24216 31249
rect 24268 31240 24270 31249
rect 24214 31175 24270 31184
rect 24596 30938 24624 32370
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 24860 31748 24912 31754
rect 24860 31690 24912 31696
rect 24872 31482 24900 31690
rect 25056 31482 25084 32166
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 24584 30184 24636 30190
rect 24584 30126 24636 30132
rect 24492 30048 24544 30054
rect 24492 29990 24544 29996
rect 24136 29702 24256 29730
rect 24504 29714 24532 29990
rect 24596 29850 24624 30126
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24124 29640 24176 29646
rect 24124 29582 24176 29588
rect 24136 29170 24164 29582
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 24136 28626 24164 29106
rect 24124 28620 24176 28626
rect 24124 28562 24176 28568
rect 24228 26790 24256 29702
rect 24492 29708 24544 29714
rect 24492 29650 24544 29656
rect 24584 29708 24636 29714
rect 24584 29650 24636 29656
rect 24504 29481 24532 29650
rect 24490 29472 24546 29481
rect 24490 29407 24546 29416
rect 24400 29232 24452 29238
rect 24400 29174 24452 29180
rect 24308 29164 24360 29170
rect 24308 29106 24360 29112
rect 24320 28694 24348 29106
rect 24412 28694 24440 29174
rect 24596 29034 24624 29650
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24308 28688 24360 28694
rect 24308 28630 24360 28636
rect 24400 28688 24452 28694
rect 24400 28630 24452 28636
rect 24320 28490 24348 28630
rect 24308 28484 24360 28490
rect 24308 28426 24360 28432
rect 24492 27872 24544 27878
rect 24492 27814 24544 27820
rect 24504 27674 24532 27814
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24688 27538 24716 29990
rect 25240 29782 25268 31282
rect 25320 30728 25372 30734
rect 25320 30670 25372 30676
rect 25228 29776 25280 29782
rect 25228 29718 25280 29724
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24780 29306 24808 29582
rect 24950 29472 25006 29481
rect 24950 29407 25006 29416
rect 24768 29300 24820 29306
rect 24768 29242 24820 29248
rect 24964 27878 24992 29407
rect 25240 29306 25268 29718
rect 25332 29578 25360 30670
rect 25320 29572 25372 29578
rect 25320 29514 25372 29520
rect 25228 29300 25280 29306
rect 25228 29242 25280 29248
rect 25240 29170 25268 29242
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25044 28960 25096 28966
rect 25044 28902 25096 28908
rect 25056 28150 25084 28902
rect 25044 28144 25096 28150
rect 25044 28086 25096 28092
rect 25240 28082 25268 29106
rect 25332 28082 25360 29514
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25320 28076 25372 28082
rect 25320 28018 25372 28024
rect 24952 27872 25004 27878
rect 24952 27814 25004 27820
rect 25240 27674 25268 28018
rect 25318 27704 25374 27713
rect 25228 27668 25280 27674
rect 25318 27639 25374 27648
rect 25228 27610 25280 27616
rect 24400 27532 24452 27538
rect 24400 27474 24452 27480
rect 24676 27532 24728 27538
rect 24676 27474 24728 27480
rect 24412 26994 24440 27474
rect 25240 27130 25268 27610
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24228 26382 24256 26726
rect 24412 26450 24440 26930
rect 25332 26926 25360 27639
rect 25424 27010 25452 33458
rect 25608 32434 25636 34614
rect 25884 34202 25912 42502
rect 26068 41682 26096 42502
rect 26252 42362 26280 43182
rect 33784 43104 33836 43110
rect 33784 43046 33836 43052
rect 33140 42900 33192 42906
rect 33140 42842 33192 42848
rect 29552 42764 29604 42770
rect 29552 42706 29604 42712
rect 31760 42764 31812 42770
rect 31760 42706 31812 42712
rect 27620 42628 27672 42634
rect 27620 42570 27672 42576
rect 28724 42628 28776 42634
rect 28724 42570 28776 42576
rect 26424 42560 26476 42566
rect 26424 42502 26476 42508
rect 26792 42560 26844 42566
rect 26792 42502 26844 42508
rect 26436 42362 26464 42502
rect 26240 42356 26292 42362
rect 26240 42298 26292 42304
rect 26424 42356 26476 42362
rect 26424 42298 26476 42304
rect 26700 42220 26752 42226
rect 26700 42162 26752 42168
rect 26240 42152 26292 42158
rect 26240 42094 26292 42100
rect 26252 41818 26280 42094
rect 26240 41812 26292 41818
rect 26240 41754 26292 41760
rect 26056 41676 26108 41682
rect 26056 41618 26108 41624
rect 26252 41274 26280 41754
rect 26712 41546 26740 42162
rect 26700 41540 26752 41546
rect 26700 41482 26752 41488
rect 26608 41472 26660 41478
rect 26608 41414 26660 41420
rect 26148 41268 26200 41274
rect 26148 41210 26200 41216
rect 26240 41268 26292 41274
rect 26240 41210 26292 41216
rect 26160 41154 26188 41210
rect 26160 41138 26280 41154
rect 26620 41138 26648 41414
rect 26160 41132 26292 41138
rect 26160 41126 26240 41132
rect 26240 41074 26292 41080
rect 26608 41132 26660 41138
rect 26608 41074 26660 41080
rect 26056 40928 26108 40934
rect 26056 40870 26108 40876
rect 26424 40928 26476 40934
rect 26424 40870 26476 40876
rect 26068 40662 26096 40870
rect 26056 40656 26108 40662
rect 26056 40598 26108 40604
rect 26436 40526 26464 40870
rect 26424 40520 26476 40526
rect 26424 40462 26476 40468
rect 26056 40384 26108 40390
rect 26056 40326 26108 40332
rect 26068 39982 26096 40326
rect 26056 39976 26108 39982
rect 26056 39918 26108 39924
rect 26700 38752 26752 38758
rect 26700 38694 26752 38700
rect 26712 38350 26740 38694
rect 26700 38344 26752 38350
rect 26700 38286 26752 38292
rect 26424 37936 26476 37942
rect 26424 37878 26476 37884
rect 26240 35828 26292 35834
rect 26240 35770 26292 35776
rect 26252 35086 26280 35770
rect 26332 35488 26384 35494
rect 26332 35430 26384 35436
rect 26344 35154 26372 35430
rect 26332 35148 26384 35154
rect 26332 35090 26384 35096
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 25872 34196 25924 34202
rect 25872 34138 25924 34144
rect 26436 34066 26464 37878
rect 26516 37664 26568 37670
rect 26516 37606 26568 37612
rect 26528 37330 26556 37606
rect 26516 37324 26568 37330
rect 26516 37266 26568 37272
rect 26424 34060 26476 34066
rect 26424 34002 26476 34008
rect 26240 33856 26292 33862
rect 26240 33798 26292 33804
rect 26332 33856 26384 33862
rect 26332 33798 26384 33804
rect 26252 33590 26280 33798
rect 26240 33584 26292 33590
rect 26240 33526 26292 33532
rect 26344 33522 26372 33798
rect 26332 33516 26384 33522
rect 26332 33458 26384 33464
rect 25964 33448 26016 33454
rect 25964 33390 26016 33396
rect 25780 32836 25832 32842
rect 25780 32778 25832 32784
rect 25596 32428 25648 32434
rect 25596 32370 25648 32376
rect 25608 32026 25636 32370
rect 25792 32298 25820 32778
rect 25976 32314 26004 33390
rect 26056 33312 26108 33318
rect 26056 33254 26108 33260
rect 26068 32502 26096 33254
rect 26344 33114 26372 33458
rect 26436 33454 26464 34002
rect 26700 33924 26752 33930
rect 26700 33866 26752 33872
rect 26424 33448 26476 33454
rect 26424 33390 26476 33396
rect 26332 33108 26384 33114
rect 26332 33050 26384 33056
rect 26056 32496 26108 32502
rect 26056 32438 26108 32444
rect 26332 32496 26384 32502
rect 26332 32438 26384 32444
rect 26056 32360 26108 32366
rect 25976 32308 26056 32314
rect 25976 32302 26108 32308
rect 25780 32292 25832 32298
rect 25976 32286 26096 32302
rect 25780 32234 25832 32240
rect 25596 32020 25648 32026
rect 25596 31962 25648 31968
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 25792 30802 25820 31758
rect 26068 31278 26096 32286
rect 26148 31748 26200 31754
rect 26148 31690 26200 31696
rect 26160 31482 26188 31690
rect 26148 31476 26200 31482
rect 26148 31418 26200 31424
rect 26056 31272 26108 31278
rect 26056 31214 26108 31220
rect 25688 30796 25740 30802
rect 25688 30738 25740 30744
rect 25780 30796 25832 30802
rect 25780 30738 25832 30744
rect 25700 30394 25728 30738
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 25688 30388 25740 30394
rect 25688 30330 25740 30336
rect 26252 30326 26280 30534
rect 26148 30320 26200 30326
rect 26148 30262 26200 30268
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 26160 30172 26188 30262
rect 26160 30144 26280 30172
rect 26056 30116 26108 30122
rect 26056 30058 26108 30064
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25504 29504 25556 29510
rect 25504 29446 25556 29452
rect 25516 28014 25544 29446
rect 25608 29102 25636 29582
rect 25686 29336 25742 29345
rect 25686 29271 25742 29280
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 25700 28558 25728 29271
rect 25792 29170 25820 29582
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25884 29238 25912 29446
rect 25872 29232 25924 29238
rect 25872 29174 25924 29180
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 25792 28762 25820 29106
rect 25780 28756 25832 28762
rect 25780 28698 25832 28704
rect 25688 28552 25740 28558
rect 25884 28540 25912 29174
rect 26068 28694 26096 30058
rect 26148 30048 26200 30054
rect 26148 29990 26200 29996
rect 26160 29481 26188 29990
rect 26146 29472 26202 29481
rect 26146 29407 26202 29416
rect 26160 28762 26188 29407
rect 26252 29209 26280 30144
rect 26238 29200 26294 29209
rect 26238 29135 26294 29144
rect 26148 28756 26200 28762
rect 26148 28698 26200 28704
rect 26056 28688 26108 28694
rect 26056 28630 26108 28636
rect 25964 28552 26016 28558
rect 25884 28512 25964 28540
rect 25688 28494 25740 28500
rect 25964 28494 26016 28500
rect 25700 28014 25728 28494
rect 26068 28422 26096 28630
rect 26056 28416 26108 28422
rect 26056 28358 26108 28364
rect 25780 28076 25832 28082
rect 25780 28018 25832 28024
rect 25504 28008 25556 28014
rect 25504 27950 25556 27956
rect 25688 28008 25740 28014
rect 25688 27950 25740 27956
rect 25424 26994 25544 27010
rect 25424 26988 25556 26994
rect 25424 26982 25504 26988
rect 25504 26930 25556 26936
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25412 26920 25464 26926
rect 25412 26862 25464 26868
rect 24400 26444 24452 26450
rect 24400 26386 24452 26392
rect 24216 26376 24268 26382
rect 24216 26318 24268 26324
rect 24228 24342 24256 26318
rect 24860 26308 24912 26314
rect 24860 26250 24912 26256
rect 24872 26042 24900 26250
rect 24860 26036 24912 26042
rect 24860 25978 24912 25984
rect 25228 25968 25280 25974
rect 25228 25910 25280 25916
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24964 25498 24992 25842
rect 25044 25696 25096 25702
rect 25044 25638 25096 25644
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24216 24336 24268 24342
rect 24216 24278 24268 24284
rect 24228 23730 24256 24278
rect 24596 24206 24624 25230
rect 24676 24812 24728 24818
rect 24676 24754 24728 24760
rect 24688 24274 24716 24754
rect 25056 24750 25084 25638
rect 25240 24818 25268 25910
rect 25424 25294 25452 26862
rect 25516 26246 25544 26930
rect 25792 26926 25820 28018
rect 26252 27402 26280 29135
rect 26344 28490 26372 32438
rect 26516 30252 26568 30258
rect 26516 30194 26568 30200
rect 26528 29850 26556 30194
rect 26608 30184 26660 30190
rect 26608 30126 26660 30132
rect 26620 29850 26648 30126
rect 26516 29844 26568 29850
rect 26516 29786 26568 29792
rect 26608 29844 26660 29850
rect 26608 29786 26660 29792
rect 26608 29708 26660 29714
rect 26608 29650 26660 29656
rect 26516 29640 26568 29646
rect 26516 29582 26568 29588
rect 26528 29510 26556 29582
rect 26516 29504 26568 29510
rect 26516 29446 26568 29452
rect 26620 29238 26648 29650
rect 26608 29232 26660 29238
rect 26608 29174 26660 29180
rect 26608 29096 26660 29102
rect 26608 29038 26660 29044
rect 26424 28960 26476 28966
rect 26424 28902 26476 28908
rect 26436 28694 26464 28902
rect 26424 28688 26476 28694
rect 26424 28630 26476 28636
rect 26516 28552 26568 28558
rect 26620 28540 26648 29038
rect 26568 28512 26648 28540
rect 26516 28494 26568 28500
rect 26332 28484 26384 28490
rect 26332 28426 26384 28432
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 25780 26920 25832 26926
rect 25780 26862 25832 26868
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25516 25906 25544 26182
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 25516 25430 25544 25842
rect 25504 25424 25556 25430
rect 25504 25366 25556 25372
rect 25412 25288 25464 25294
rect 25412 25230 25464 25236
rect 25320 25220 25372 25226
rect 25320 25162 25372 25168
rect 25332 24954 25360 25162
rect 25320 24948 25372 24954
rect 25320 24890 25372 24896
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 24860 24676 24912 24682
rect 24860 24618 24912 24624
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24872 24206 24900 24618
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24584 24064 24636 24070
rect 24636 24012 24900 24018
rect 24584 24006 24900 24012
rect 24596 23990 24900 24006
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24320 23526 24348 23666
rect 24308 23520 24360 23526
rect 24308 23462 24360 23468
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24216 22772 24268 22778
rect 24216 22714 24268 22720
rect 24124 22500 24176 22506
rect 24124 22442 24176 22448
rect 24032 22160 24084 22166
rect 24032 22102 24084 22108
rect 24136 22098 24164 22442
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 23768 21350 23796 22034
rect 24228 21622 24256 22714
rect 24688 22710 24716 23054
rect 24872 22710 24900 23990
rect 24964 23866 24992 24142
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25056 23662 25084 24686
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 25226 24440 25282 24449
rect 25226 24375 25282 24384
rect 25136 24336 25188 24342
rect 25136 24278 25188 24284
rect 25148 24206 25176 24278
rect 25240 24206 25268 24375
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 24676 22704 24728 22710
rect 24676 22646 24728 22652
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24216 21616 24268 21622
rect 24216 21558 24268 21564
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 24780 21010 24808 22646
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24872 21690 24900 22510
rect 25148 22030 25176 23462
rect 25228 23044 25280 23050
rect 25228 22986 25280 22992
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 24952 21888 25004 21894
rect 25240 21876 25268 22986
rect 25004 21848 25268 21876
rect 24952 21830 25004 21836
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 25240 21554 25268 21848
rect 25332 21622 25360 24550
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23768 19242 23796 19790
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 23756 19236 23808 19242
rect 23756 19178 23808 19184
rect 23584 18142 23704 18170
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23492 12782 23520 13670
rect 23584 13462 23612 18142
rect 23768 18034 23796 19178
rect 24136 18970 24164 19246
rect 24964 18970 24992 20946
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 24400 18692 24452 18698
rect 24400 18634 24452 18640
rect 24308 18216 24360 18222
rect 24308 18158 24360 18164
rect 23676 18006 23796 18034
rect 23676 15502 23704 18006
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23768 17270 23796 17818
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23860 16794 23888 17138
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24136 16250 24164 16594
rect 24216 16584 24268 16590
rect 24216 16526 24268 16532
rect 24228 16250 24256 16526
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 23756 16176 23808 16182
rect 23756 16118 23808 16124
rect 23768 15570 23796 16118
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23952 15502 23980 16050
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23952 15366 23980 15438
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 23756 14340 23808 14346
rect 23756 14282 23808 14288
rect 23768 14074 23796 14282
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 24136 14006 24164 14758
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 23572 13456 23624 13462
rect 23572 13398 23624 13404
rect 23584 12850 23612 13398
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23676 12374 23704 12718
rect 23768 12434 23796 13126
rect 23768 12406 24164 12434
rect 23664 12368 23716 12374
rect 23664 12310 23716 12316
rect 24136 12238 24164 12406
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24136 11830 24164 12174
rect 24124 11824 24176 11830
rect 24124 11766 24176 11772
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24136 11218 24164 11494
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23308 10266 23336 10950
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 22940 8758 23152 8786
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21284 7478 21312 7686
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21192 6390 21220 6666
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 21180 6384 21232 6390
rect 21180 6326 21232 6332
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 21744 5914 21772 6666
rect 21836 6322 21864 7142
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 22112 5234 22140 5578
rect 22204 5302 22232 7890
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22296 5302 22324 7482
rect 22468 6656 22520 6662
rect 22468 6598 22520 6604
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22388 5098 22416 5646
rect 22480 5234 22508 6598
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22664 5642 22692 6054
rect 22848 5710 22876 8570
rect 22940 7886 22968 8758
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22652 5636 22704 5642
rect 22652 5578 22704 5584
rect 22940 5574 22968 7822
rect 23032 6662 23060 8434
rect 23216 7478 23244 9590
rect 23308 9518 23336 9998
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 23400 9178 23428 9998
rect 23676 9722 23704 9998
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23768 9654 23796 10406
rect 24136 10130 24164 11154
rect 24228 10674 24256 13262
rect 24320 12442 24348 18158
rect 24412 17882 24440 18634
rect 24964 18222 24992 18906
rect 25056 18358 25084 19654
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 24952 18216 25004 18222
rect 24952 18158 25004 18164
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 24400 17264 24452 17270
rect 24400 17206 24452 17212
rect 24412 16794 24440 17206
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24504 14958 24532 17070
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24780 16046 24808 16730
rect 24964 16590 24992 17682
rect 25056 17610 25084 18294
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 25056 17270 25084 17546
rect 25044 17264 25096 17270
rect 25044 17206 25096 17212
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24780 15638 24808 15982
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24872 14362 24900 16186
rect 25056 16114 25084 16390
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25056 15978 25084 16050
rect 25044 15972 25096 15978
rect 25044 15914 25096 15920
rect 25056 15502 25084 15914
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25148 15314 25176 21490
rect 25240 20788 25268 21490
rect 25320 20800 25372 20806
rect 25240 20760 25320 20788
rect 25320 20742 25372 20748
rect 25424 19514 25452 25230
rect 25516 24750 25544 25366
rect 25504 24744 25556 24750
rect 25608 24721 25636 26726
rect 26252 26382 26280 27338
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26240 25492 26292 25498
rect 26240 25434 26292 25440
rect 25872 25220 25924 25226
rect 25872 25162 25924 25168
rect 25884 24886 25912 25162
rect 25688 24880 25740 24886
rect 25688 24822 25740 24828
rect 25872 24880 25924 24886
rect 26056 24880 26108 24886
rect 25924 24840 26056 24868
rect 25872 24822 25924 24828
rect 26056 24822 26108 24828
rect 25700 24750 25728 24822
rect 25688 24744 25740 24750
rect 25504 24686 25556 24692
rect 25594 24712 25650 24721
rect 25688 24686 25740 24692
rect 25594 24647 25650 24656
rect 25608 24596 25636 24647
rect 25516 24568 25636 24596
rect 25516 23118 25544 24568
rect 25700 24206 25728 24686
rect 26252 24682 26280 25434
rect 26344 24818 26372 28426
rect 26516 28416 26568 28422
rect 26514 28384 26516 28393
rect 26568 28384 26570 28393
rect 26514 28319 26570 28328
rect 26424 28144 26476 28150
rect 26424 28086 26476 28092
rect 26436 26994 26464 28086
rect 26608 28076 26660 28082
rect 26608 28018 26660 28024
rect 26516 27872 26568 27878
rect 26516 27814 26568 27820
rect 26528 27470 26556 27814
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26514 27024 26570 27033
rect 26424 26988 26476 26994
rect 26620 27010 26648 28018
rect 26712 27062 26740 33866
rect 26804 33658 26832 42502
rect 27632 42362 27660 42570
rect 27620 42356 27672 42362
rect 27620 42298 27672 42304
rect 26884 42288 26936 42294
rect 26884 42230 26936 42236
rect 26896 41614 26924 42230
rect 27712 42152 27764 42158
rect 27712 42094 27764 42100
rect 27068 42016 27120 42022
rect 27068 41958 27120 41964
rect 26884 41608 26936 41614
rect 26884 41550 26936 41556
rect 27080 41002 27108 41958
rect 27068 40996 27120 41002
rect 27068 40938 27120 40944
rect 27620 40384 27672 40390
rect 27620 40326 27672 40332
rect 27632 40118 27660 40326
rect 27620 40112 27672 40118
rect 27620 40054 27672 40060
rect 26976 39976 27028 39982
rect 26976 39918 27028 39924
rect 26988 38758 27016 39918
rect 26976 38752 27028 38758
rect 26976 38694 27028 38700
rect 26988 38350 27016 38694
rect 27252 38480 27304 38486
rect 27252 38422 27304 38428
rect 26976 38344 27028 38350
rect 26976 38286 27028 38292
rect 27160 38208 27212 38214
rect 27160 38150 27212 38156
rect 27172 37874 27200 38150
rect 27264 37874 27292 38422
rect 27528 38412 27580 38418
rect 27528 38354 27580 38360
rect 27540 38321 27568 38354
rect 27526 38312 27582 38321
rect 27526 38247 27582 38256
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 27252 37868 27304 37874
rect 27252 37810 27304 37816
rect 27620 37664 27672 37670
rect 27620 37606 27672 37612
rect 27068 37460 27120 37466
rect 27068 37402 27120 37408
rect 27080 36174 27108 37402
rect 27632 37262 27660 37606
rect 27620 37256 27672 37262
rect 27620 37198 27672 37204
rect 27344 36712 27396 36718
rect 27344 36654 27396 36660
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 27080 35018 27108 36110
rect 27356 36038 27384 36654
rect 27632 36650 27660 37198
rect 27620 36644 27672 36650
rect 27620 36586 27672 36592
rect 27344 36032 27396 36038
rect 27344 35974 27396 35980
rect 27068 35012 27120 35018
rect 27068 34954 27120 34960
rect 27160 35012 27212 35018
rect 27160 34954 27212 34960
rect 27080 33930 27108 34954
rect 27172 34746 27200 34954
rect 27160 34740 27212 34746
rect 27160 34682 27212 34688
rect 27068 33924 27120 33930
rect 27068 33866 27120 33872
rect 26792 33652 26844 33658
rect 26792 33594 26844 33600
rect 27080 32910 27108 33866
rect 27252 33584 27304 33590
rect 27252 33526 27304 33532
rect 27068 32904 27120 32910
rect 27068 32846 27120 32852
rect 27080 31822 27108 32846
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 27068 31816 27120 31822
rect 27068 31758 27120 31764
rect 26792 31408 26844 31414
rect 26792 31350 26844 31356
rect 26804 30598 26832 31350
rect 26792 30592 26844 30598
rect 26792 30534 26844 30540
rect 26804 30258 26832 30534
rect 26792 30252 26844 30258
rect 26792 30194 26844 30200
rect 26804 29646 26832 30194
rect 26792 29640 26844 29646
rect 26792 29582 26844 29588
rect 26804 29306 26832 29582
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26804 29102 26832 29242
rect 27172 29238 27200 32370
rect 27264 32026 27292 33526
rect 27252 32020 27304 32026
rect 27252 31962 27304 31968
rect 27264 31346 27292 31962
rect 27356 31906 27384 35974
rect 27724 34202 27752 42094
rect 27896 42084 27948 42090
rect 27896 42026 27948 42032
rect 27804 41132 27856 41138
rect 27804 41074 27856 41080
rect 27816 40905 27844 41074
rect 27802 40896 27858 40905
rect 27802 40831 27858 40840
rect 27908 40730 27936 42026
rect 28736 41818 28764 42570
rect 29000 42560 29052 42566
rect 29000 42502 29052 42508
rect 29012 42226 29040 42502
rect 29000 42220 29052 42226
rect 29000 42162 29052 42168
rect 28724 41812 28776 41818
rect 28724 41754 28776 41760
rect 28080 41744 28132 41750
rect 28080 41686 28132 41692
rect 28092 41138 28120 41686
rect 28172 41608 28224 41614
rect 28172 41550 28224 41556
rect 28184 41274 28212 41550
rect 28632 41472 28684 41478
rect 28632 41414 28684 41420
rect 28552 41386 28672 41414
rect 28172 41268 28224 41274
rect 28172 41210 28224 41216
rect 28264 41268 28316 41274
rect 28264 41210 28316 41216
rect 28080 41132 28132 41138
rect 28080 41074 28132 41080
rect 27896 40724 27948 40730
rect 27896 40666 27948 40672
rect 28092 40526 28120 41074
rect 28276 41002 28304 41210
rect 28552 41138 28580 41386
rect 28736 41290 28764 41754
rect 29012 41750 29040 42162
rect 29000 41744 29052 41750
rect 29000 41686 29052 41692
rect 29564 41682 29592 42706
rect 29828 42628 29880 42634
rect 29828 42570 29880 42576
rect 30472 42628 30524 42634
rect 30472 42570 30524 42576
rect 29840 42362 29868 42570
rect 29828 42356 29880 42362
rect 29828 42298 29880 42304
rect 30104 42152 30156 42158
rect 30104 42094 30156 42100
rect 29552 41676 29604 41682
rect 29552 41618 29604 41624
rect 29736 41676 29788 41682
rect 29736 41618 29788 41624
rect 29276 41608 29328 41614
rect 29276 41550 29328 41556
rect 29184 41540 29236 41546
rect 29184 41482 29236 41488
rect 28644 41262 28764 41290
rect 28908 41268 28960 41274
rect 28540 41132 28592 41138
rect 28540 41074 28592 41080
rect 28356 41064 28408 41070
rect 28356 41006 28408 41012
rect 28264 40996 28316 41002
rect 28264 40938 28316 40944
rect 28172 40724 28224 40730
rect 28172 40666 28224 40672
rect 27804 40520 27856 40526
rect 27804 40462 27856 40468
rect 27988 40520 28040 40526
rect 28080 40520 28132 40526
rect 27988 40462 28040 40468
rect 28078 40488 28080 40497
rect 28132 40488 28134 40497
rect 27816 40361 27844 40462
rect 27896 40384 27948 40390
rect 27802 40352 27858 40361
rect 27896 40326 27948 40332
rect 27802 40287 27858 40296
rect 27908 39982 27936 40326
rect 28000 40186 28028 40462
rect 28078 40423 28134 40432
rect 27988 40180 28040 40186
rect 27988 40122 28040 40128
rect 27896 39976 27948 39982
rect 27896 39918 27948 39924
rect 27896 37800 27948 37806
rect 27896 37742 27948 37748
rect 27908 37126 27936 37742
rect 27896 37120 27948 37126
rect 27896 37062 27948 37068
rect 27804 36100 27856 36106
rect 27804 36042 27856 36048
rect 27816 35834 27844 36042
rect 27804 35828 27856 35834
rect 27804 35770 27856 35776
rect 27712 34196 27764 34202
rect 27712 34138 27764 34144
rect 27436 32836 27488 32842
rect 27436 32778 27488 32784
rect 27448 32298 27476 32778
rect 27436 32292 27488 32298
rect 27436 32234 27488 32240
rect 27356 31878 27568 31906
rect 27252 31340 27304 31346
rect 27252 31282 27304 31288
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27436 29640 27488 29646
rect 27436 29582 27488 29588
rect 27252 29572 27304 29578
rect 27252 29514 27304 29520
rect 27160 29232 27212 29238
rect 27160 29174 27212 29180
rect 26792 29096 26844 29102
rect 26792 29038 26844 29044
rect 27068 28960 27120 28966
rect 27068 28902 27120 28908
rect 26884 28620 26936 28626
rect 26884 28562 26936 28568
rect 26790 28520 26846 28529
rect 26790 28455 26846 28464
rect 26804 28422 26832 28455
rect 26792 28416 26844 28422
rect 26792 28358 26844 28364
rect 26570 26982 26648 27010
rect 26700 27056 26752 27062
rect 26700 26998 26752 27004
rect 26514 26959 26516 26968
rect 26424 26930 26476 26936
rect 26568 26959 26570 26968
rect 26516 26930 26568 26936
rect 26804 26874 26832 28358
rect 26896 27713 26924 28562
rect 27080 28558 27108 28902
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 26882 27704 26938 27713
rect 26882 27639 26938 27648
rect 27172 27606 27200 29174
rect 27264 27946 27292 29514
rect 27356 29170 27384 29582
rect 27448 29306 27476 29582
rect 27436 29300 27488 29306
rect 27436 29242 27488 29248
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27252 27940 27304 27946
rect 27252 27882 27304 27888
rect 27264 27674 27292 27882
rect 27252 27668 27304 27674
rect 27252 27610 27304 27616
rect 27160 27600 27212 27606
rect 27160 27542 27212 27548
rect 27172 27130 27200 27542
rect 27160 27124 27212 27130
rect 27160 27066 27212 27072
rect 26620 26846 26832 26874
rect 26332 24812 26384 24818
rect 26332 24754 26384 24760
rect 26516 24744 26568 24750
rect 26516 24686 26568 24692
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 25596 24132 25648 24138
rect 25596 24074 25648 24080
rect 25608 23202 25636 24074
rect 25700 23594 25728 24142
rect 25688 23588 25740 23594
rect 25688 23530 25740 23536
rect 25792 23526 25820 24210
rect 26068 24206 26096 24550
rect 26252 24206 26280 24618
rect 26528 24449 26556 24686
rect 26514 24440 26570 24449
rect 26514 24375 26570 24384
rect 26528 24206 26556 24375
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26148 24132 26200 24138
rect 26148 24074 26200 24080
rect 26160 24018 26188 24074
rect 26160 23990 26280 24018
rect 26252 23798 26280 23990
rect 26148 23792 26200 23798
rect 26148 23734 26200 23740
rect 26240 23792 26292 23798
rect 26240 23734 26292 23740
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 25872 23588 25924 23594
rect 25872 23530 25924 23536
rect 25780 23520 25832 23526
rect 25780 23462 25832 23468
rect 25608 23174 25728 23202
rect 25504 23112 25556 23118
rect 25504 23054 25556 23060
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25608 22778 25636 23054
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25516 20534 25544 22578
rect 25700 22094 25728 23174
rect 25884 23118 25912 23530
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25964 23112 26016 23118
rect 25964 23054 26016 23060
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25792 22234 25820 22578
rect 25976 22438 26004 23054
rect 25964 22432 26016 22438
rect 25964 22374 26016 22380
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 25700 22066 25912 22094
rect 25596 21956 25648 21962
rect 25596 21898 25648 21904
rect 25608 21690 25636 21898
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25700 21690 25728 21830
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25884 21026 25912 22066
rect 25976 21554 26004 22374
rect 25964 21548 26016 21554
rect 25964 21490 26016 21496
rect 25976 21350 26004 21490
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25700 20998 25912 21026
rect 25504 20528 25556 20534
rect 25504 20470 25556 20476
rect 25516 19718 25544 20470
rect 25504 19712 25556 19718
rect 25504 19654 25556 19660
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25240 18766 25268 19110
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25240 17746 25268 18702
rect 25424 18630 25452 19450
rect 25516 19446 25544 19654
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25516 17746 25544 18022
rect 25228 17740 25280 17746
rect 25228 17682 25280 17688
rect 25504 17740 25556 17746
rect 25504 17682 25556 17688
rect 25240 17338 25268 17682
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 25504 17060 25556 17066
rect 25504 17002 25556 17008
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 24688 14334 24900 14362
rect 24964 15286 25176 15314
rect 24688 13326 24716 14334
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24780 14006 24808 14214
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24308 12436 24360 12442
rect 24308 12378 24360 12384
rect 24780 12238 24808 13942
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24872 12646 24900 13330
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24964 12306 24992 15286
rect 25424 15042 25452 16934
rect 25516 16590 25544 17002
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25608 16250 25636 16526
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 25608 15201 25636 15302
rect 25594 15192 25650 15201
rect 25594 15127 25650 15136
rect 25332 15014 25452 15042
rect 25332 14958 25360 15014
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25320 14340 25372 14346
rect 25320 14282 25372 14288
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25148 13326 25176 14010
rect 25228 13456 25280 13462
rect 25332 13444 25360 14282
rect 25280 13416 25360 13444
rect 25228 13398 25280 13404
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25148 12918 25176 13262
rect 25136 12912 25188 12918
rect 25136 12854 25188 12860
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24504 11830 24532 12038
rect 24492 11824 24544 11830
rect 24492 11766 24544 11772
rect 24860 11552 24912 11558
rect 24860 11494 24912 11500
rect 24872 11286 24900 11494
rect 24860 11280 24912 11286
rect 24860 11222 24912 11228
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24228 10554 24256 10610
rect 25148 10606 25176 12582
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25240 11558 25268 12378
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 25240 10810 25268 11018
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25136 10600 25188 10606
rect 24228 10526 24348 10554
rect 25136 10542 25188 10548
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23572 9512 23624 9518
rect 23572 9454 23624 9460
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23204 7472 23256 7478
rect 23204 7414 23256 7420
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23308 5914 23336 7278
rect 23400 6730 23428 7414
rect 23584 7342 23612 9454
rect 24216 9104 24268 9110
rect 24216 9046 24268 9052
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23768 7546 23796 8230
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 23584 6866 23612 7278
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23400 6458 23428 6666
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23492 6254 23520 6598
rect 23584 6390 23612 6802
rect 23768 6798 23796 7482
rect 24136 7410 24164 7958
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24136 7002 24164 7346
rect 24124 6996 24176 7002
rect 24124 6938 24176 6944
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23768 5778 23796 6734
rect 24228 6730 24256 9046
rect 24320 8294 24348 10526
rect 25044 10124 25096 10130
rect 24964 10084 25044 10112
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24596 9178 24624 9454
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24320 7478 24348 8230
rect 24412 7954 24440 8366
rect 24492 8356 24544 8362
rect 24492 8298 24544 8304
rect 24504 7954 24532 8298
rect 24400 7948 24452 7954
rect 24400 7890 24452 7896
rect 24492 7948 24544 7954
rect 24492 7890 24544 7896
rect 24412 7478 24440 7890
rect 24780 7478 24808 8910
rect 24964 7750 24992 10084
rect 25044 10066 25096 10072
rect 25044 9988 25096 9994
rect 25044 9930 25096 9936
rect 25056 8974 25084 9930
rect 25148 9466 25176 10542
rect 25148 9438 25268 9466
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 25148 9042 25176 9318
rect 25136 9036 25188 9042
rect 25136 8978 25188 8984
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25056 8480 25084 8774
rect 25148 8634 25176 8978
rect 25240 8634 25268 9438
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25136 8492 25188 8498
rect 25056 8452 25136 8480
rect 25136 8434 25188 8440
rect 25148 7954 25176 8434
rect 25240 8430 25268 8570
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25332 7886 25360 12786
rect 25424 9450 25452 15014
rect 25596 14952 25648 14958
rect 25596 14894 25648 14900
rect 25608 14074 25636 14894
rect 25700 14090 25728 20998
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25792 20602 25820 20878
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25792 16810 25820 20538
rect 25884 20398 25912 20742
rect 25976 20466 26004 21286
rect 26068 20534 26096 23666
rect 26160 22930 26188 23734
rect 26424 22976 26476 22982
rect 26160 22902 26280 22930
rect 26424 22918 26476 22924
rect 26252 22778 26280 22902
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 26056 20528 26108 20534
rect 26056 20470 26108 20476
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 25872 20392 25924 20398
rect 25872 20334 25924 20340
rect 25964 19168 26016 19174
rect 25964 19110 26016 19116
rect 25976 18766 26004 19110
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 26160 17252 26188 22714
rect 26252 22574 26280 22714
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26436 21962 26464 22918
rect 26516 22500 26568 22506
rect 26516 22442 26568 22448
rect 26424 21956 26476 21962
rect 26424 21898 26476 21904
rect 26332 20868 26384 20874
rect 26332 20810 26384 20816
rect 26344 20602 26372 20810
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26344 18426 26372 19314
rect 26528 19310 26556 22442
rect 26620 22094 26648 26846
rect 26700 26784 26752 26790
rect 26700 26726 26752 26732
rect 26712 25430 26740 26726
rect 26700 25424 26752 25430
rect 26700 25366 26752 25372
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 27160 25288 27212 25294
rect 27160 25230 27212 25236
rect 26700 24608 26752 24614
rect 26700 24550 26752 24556
rect 26712 24188 26740 24550
rect 26988 24410 27016 25230
rect 27172 24682 27200 25230
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27252 24676 27304 24682
rect 27252 24618 27304 24624
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26792 24200 26844 24206
rect 26712 24160 26792 24188
rect 26792 24142 26844 24148
rect 26804 23662 26832 24142
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 27172 23866 27200 24074
rect 27160 23860 27212 23866
rect 27160 23802 27212 23808
rect 26792 23656 26844 23662
rect 26792 23598 26844 23604
rect 27264 23594 27292 24618
rect 27356 23798 27384 29106
rect 27540 28642 27568 31878
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 27724 30938 27752 31690
rect 27712 30932 27764 30938
rect 27712 30874 27764 30880
rect 27804 30388 27856 30394
rect 27804 30330 27856 30336
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27448 28614 27568 28642
rect 27448 28150 27476 28614
rect 27632 28558 27660 29582
rect 27816 29238 27844 30330
rect 27908 29714 27936 37062
rect 28184 34542 28212 40666
rect 28368 40390 28396 41006
rect 28448 40928 28500 40934
rect 28448 40870 28500 40876
rect 28356 40384 28408 40390
rect 28460 40361 28488 40870
rect 28552 40594 28580 41074
rect 28644 41018 28672 41262
rect 28908 41210 28960 41216
rect 28920 41138 28948 41210
rect 29196 41206 29224 41482
rect 29184 41200 29236 41206
rect 29184 41142 29236 41148
rect 28908 41132 28960 41138
rect 28908 41074 28960 41080
rect 29092 41132 29144 41138
rect 29092 41074 29144 41080
rect 28644 40990 28764 41018
rect 28632 40928 28684 40934
rect 28630 40896 28632 40905
rect 28736 40916 28764 40990
rect 28684 40896 28686 40905
rect 28736 40888 28856 40916
rect 28630 40831 28686 40840
rect 28724 40656 28776 40662
rect 28724 40598 28776 40604
rect 28540 40588 28592 40594
rect 28540 40530 28592 40536
rect 28356 40326 28408 40332
rect 28446 40352 28502 40361
rect 28446 40287 28502 40296
rect 28552 40186 28580 40530
rect 28540 40180 28592 40186
rect 28540 40122 28592 40128
rect 28356 39908 28408 39914
rect 28356 39850 28408 39856
rect 28368 38962 28396 39850
rect 28540 39092 28592 39098
rect 28540 39034 28592 39040
rect 28356 38956 28408 38962
rect 28356 38898 28408 38904
rect 28368 38418 28396 38898
rect 28448 38752 28500 38758
rect 28448 38694 28500 38700
rect 28356 38412 28408 38418
rect 28356 38354 28408 38360
rect 28460 38350 28488 38694
rect 28264 38344 28316 38350
rect 28264 38286 28316 38292
rect 28448 38344 28500 38350
rect 28448 38286 28500 38292
rect 28276 38010 28304 38286
rect 28448 38208 28500 38214
rect 28448 38150 28500 38156
rect 28264 38004 28316 38010
rect 28264 37946 28316 37952
rect 28460 35834 28488 38150
rect 28552 37874 28580 39034
rect 28736 39030 28764 40598
rect 28828 40202 28856 40888
rect 28908 40520 28960 40526
rect 28906 40488 28908 40497
rect 28960 40488 28962 40497
rect 28906 40423 28962 40432
rect 28908 40384 28960 40390
rect 28906 40352 28908 40361
rect 28960 40352 28962 40361
rect 28906 40287 28962 40296
rect 28828 40174 28948 40202
rect 28724 39024 28776 39030
rect 28644 38984 28724 39012
rect 28644 38418 28672 38984
rect 28724 38966 28776 38972
rect 28816 38888 28868 38894
rect 28816 38830 28868 38836
rect 28724 38752 28776 38758
rect 28724 38694 28776 38700
rect 28632 38412 28684 38418
rect 28632 38354 28684 38360
rect 28540 37868 28592 37874
rect 28540 37810 28592 37816
rect 28736 37754 28764 38694
rect 28828 38282 28856 38830
rect 28816 38276 28868 38282
rect 28816 38218 28868 38224
rect 28828 37806 28856 38218
rect 28644 37738 28764 37754
rect 28816 37800 28868 37806
rect 28816 37742 28868 37748
rect 28632 37732 28764 37738
rect 28684 37726 28764 37732
rect 28632 37674 28684 37680
rect 28816 37664 28868 37670
rect 28816 37606 28868 37612
rect 28828 36718 28856 37606
rect 28920 36718 28948 40174
rect 29000 37800 29052 37806
rect 29000 37742 29052 37748
rect 29012 36922 29040 37742
rect 29000 36916 29052 36922
rect 29000 36858 29052 36864
rect 28816 36712 28868 36718
rect 28816 36654 28868 36660
rect 28908 36712 28960 36718
rect 28908 36654 28960 36660
rect 28920 36122 28948 36654
rect 28828 36106 28948 36122
rect 28828 36100 28960 36106
rect 28828 36094 28908 36100
rect 28448 35828 28500 35834
rect 28448 35770 28500 35776
rect 28828 35018 28856 36094
rect 28908 36042 28960 36048
rect 29012 35986 29040 36858
rect 29104 36854 29132 41074
rect 29288 40934 29316 41550
rect 29748 41138 29776 41618
rect 30012 41540 30064 41546
rect 30012 41482 30064 41488
rect 29736 41132 29788 41138
rect 29736 41074 29788 41080
rect 29276 40928 29328 40934
rect 29276 40870 29328 40876
rect 29092 36848 29144 36854
rect 29092 36790 29144 36796
rect 29090 36272 29146 36281
rect 29090 36207 29146 36216
rect 29104 36174 29132 36207
rect 29092 36168 29144 36174
rect 29092 36110 29144 36116
rect 28920 35958 29040 35986
rect 28920 35630 28948 35958
rect 28908 35624 28960 35630
rect 28908 35566 28960 35572
rect 28816 35012 28868 35018
rect 28816 34954 28868 34960
rect 28724 34944 28776 34950
rect 28724 34886 28776 34892
rect 28736 34746 28764 34886
rect 28724 34740 28776 34746
rect 28724 34682 28776 34688
rect 29104 34678 29132 36110
rect 29288 35290 29316 40870
rect 30024 40730 30052 41482
rect 30012 40724 30064 40730
rect 30012 40666 30064 40672
rect 30116 39642 30144 42094
rect 30484 41818 30512 42570
rect 31392 42560 31444 42566
rect 31392 42502 31444 42508
rect 31404 42362 31432 42502
rect 31392 42356 31444 42362
rect 31392 42298 31444 42304
rect 31484 42356 31536 42362
rect 31484 42298 31536 42304
rect 31496 42242 31524 42298
rect 30840 42220 30892 42226
rect 30840 42162 30892 42168
rect 31208 42220 31260 42226
rect 31208 42162 31260 42168
rect 31404 42214 31524 42242
rect 31772 42226 31800 42706
rect 32128 42696 32180 42702
rect 32128 42638 32180 42644
rect 30656 42084 30708 42090
rect 30656 42026 30708 42032
rect 30472 41812 30524 41818
rect 30472 41754 30524 41760
rect 30484 41546 30512 41754
rect 30472 41540 30524 41546
rect 30472 41482 30524 41488
rect 30472 40928 30524 40934
rect 30472 40870 30524 40876
rect 30484 40526 30512 40870
rect 30668 40594 30696 42026
rect 30852 41478 30880 42162
rect 31220 41818 31248 42162
rect 31300 42152 31352 42158
rect 31300 42094 31352 42100
rect 31208 41812 31260 41818
rect 31208 41754 31260 41760
rect 31116 41744 31168 41750
rect 31116 41686 31168 41692
rect 30840 41472 30892 41478
rect 30840 41414 30892 41420
rect 30852 41274 30880 41414
rect 30840 41268 30892 41274
rect 30840 41210 30892 41216
rect 30932 41132 30984 41138
rect 30932 41074 30984 41080
rect 30944 41041 30972 41074
rect 30930 41032 30986 41041
rect 31128 41002 31156 41686
rect 31312 41682 31340 42094
rect 31300 41676 31352 41682
rect 31300 41618 31352 41624
rect 31404 41426 31432 42214
rect 31496 42208 31524 42214
rect 31576 42220 31628 42226
rect 31496 42180 31576 42208
rect 31576 42162 31628 42168
rect 31760 42220 31812 42226
rect 31760 42162 31812 42168
rect 31852 42152 31904 42158
rect 31588 42078 31754 42106
rect 31852 42094 31904 42100
rect 31588 42022 31616 42078
rect 31576 42016 31628 42022
rect 31576 41958 31628 41964
rect 31726 41970 31754 42078
rect 31864 42022 31892 42094
rect 31852 42016 31904 42022
rect 31726 41942 31800 41970
rect 31852 41958 31904 41964
rect 31484 41812 31536 41818
rect 31484 41754 31536 41760
rect 31496 41614 31524 41754
rect 31668 41744 31720 41750
rect 31668 41686 31720 41692
rect 31484 41608 31536 41614
rect 31536 41568 31616 41596
rect 31484 41550 31536 41556
rect 31484 41472 31536 41478
rect 31404 41420 31484 41426
rect 31404 41414 31536 41420
rect 31404 41398 31524 41414
rect 31496 41274 31524 41398
rect 31484 41268 31536 41274
rect 31484 41210 31536 41216
rect 30930 40967 30986 40976
rect 31116 40996 31168 41002
rect 30656 40588 30708 40594
rect 30656 40530 30708 40536
rect 30472 40520 30524 40526
rect 30472 40462 30524 40468
rect 30564 40384 30616 40390
rect 30564 40326 30616 40332
rect 30576 39642 30604 40326
rect 30944 40089 30972 40967
rect 31116 40938 31168 40944
rect 31128 40662 31156 40938
rect 31496 40882 31524 41210
rect 31588 41138 31616 41568
rect 31680 41478 31708 41686
rect 31772 41682 31800 41942
rect 31760 41676 31812 41682
rect 31760 41618 31812 41624
rect 31668 41472 31720 41478
rect 31668 41414 31720 41420
rect 31772 41138 31800 41618
rect 31864 41614 31892 41958
rect 31852 41608 31904 41614
rect 31852 41550 31904 41556
rect 31576 41132 31628 41138
rect 31576 41074 31628 41080
rect 31760 41132 31812 41138
rect 31760 41074 31812 41080
rect 31496 40854 31708 40882
rect 31484 40724 31536 40730
rect 31484 40666 31536 40672
rect 31116 40656 31168 40662
rect 31116 40598 31168 40604
rect 30930 40080 30986 40089
rect 30930 40015 30986 40024
rect 31116 40044 31168 40050
rect 31116 39986 31168 39992
rect 30104 39636 30156 39642
rect 30104 39578 30156 39584
rect 30564 39636 30616 39642
rect 30564 39578 30616 39584
rect 31128 39574 31156 39986
rect 31116 39568 31168 39574
rect 31116 39510 31168 39516
rect 30840 39500 30892 39506
rect 30840 39442 30892 39448
rect 30564 39296 30616 39302
rect 30564 39238 30616 39244
rect 30380 38752 30432 38758
rect 30380 38694 30432 38700
rect 29552 38208 29604 38214
rect 29552 38150 29604 38156
rect 29564 38010 29592 38150
rect 29552 38004 29604 38010
rect 29552 37946 29604 37952
rect 30392 37194 30420 38694
rect 30472 37800 30524 37806
rect 30472 37742 30524 37748
rect 30380 37188 30432 37194
rect 30380 37130 30432 37136
rect 30484 36582 30512 37742
rect 29920 36576 29972 36582
rect 29920 36518 29972 36524
rect 30472 36576 30524 36582
rect 30472 36518 30524 36524
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 29564 35766 29592 35974
rect 29552 35760 29604 35766
rect 29552 35702 29604 35708
rect 29828 35488 29880 35494
rect 29828 35430 29880 35436
rect 29276 35284 29328 35290
rect 29276 35226 29328 35232
rect 29840 35154 29868 35430
rect 29828 35148 29880 35154
rect 29828 35090 29880 35096
rect 29736 35012 29788 35018
rect 29736 34954 29788 34960
rect 29092 34672 29144 34678
rect 29092 34614 29144 34620
rect 29748 34542 29776 34954
rect 27988 34536 28040 34542
rect 27988 34478 28040 34484
rect 28172 34536 28224 34542
rect 28172 34478 28224 34484
rect 28908 34536 28960 34542
rect 28908 34478 28960 34484
rect 29736 34536 29788 34542
rect 29736 34478 29788 34484
rect 28000 33658 28028 34478
rect 28724 33924 28776 33930
rect 28724 33866 28776 33872
rect 28356 33856 28408 33862
rect 28356 33798 28408 33804
rect 27988 33652 28040 33658
rect 27988 33594 28040 33600
rect 28368 33538 28396 33798
rect 28276 33522 28396 33538
rect 28736 33522 28764 33866
rect 28264 33516 28396 33522
rect 28316 33510 28396 33516
rect 28724 33516 28776 33522
rect 28264 33458 28316 33464
rect 28724 33458 28776 33464
rect 28276 33046 28304 33458
rect 28264 33040 28316 33046
rect 28264 32982 28316 32988
rect 28080 32836 28132 32842
rect 28080 32778 28132 32784
rect 28092 32434 28120 32778
rect 28080 32428 28132 32434
rect 28080 32370 28132 32376
rect 28736 31958 28764 33458
rect 28920 33454 28948 34478
rect 28908 33448 28960 33454
rect 28908 33390 28960 33396
rect 29748 32978 29776 34478
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29748 32502 29776 32914
rect 28816 32496 28868 32502
rect 28816 32438 28868 32444
rect 29736 32496 29788 32502
rect 29736 32438 29788 32444
rect 28724 31952 28776 31958
rect 28724 31894 28776 31900
rect 28356 31408 28408 31414
rect 28356 31350 28408 31356
rect 28172 31272 28224 31278
rect 28172 31214 28224 31220
rect 28184 30938 28212 31214
rect 28264 31136 28316 31142
rect 28264 31078 28316 31084
rect 28172 30932 28224 30938
rect 28172 30874 28224 30880
rect 28276 30802 28304 31078
rect 28264 30796 28316 30802
rect 28264 30738 28316 30744
rect 27896 29708 27948 29714
rect 27896 29650 27948 29656
rect 27908 29238 27936 29650
rect 27804 29232 27856 29238
rect 27804 29174 27856 29180
rect 27896 29232 27948 29238
rect 27896 29174 27948 29180
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27528 28484 27580 28490
rect 27528 28426 27580 28432
rect 27436 28144 27488 28150
rect 27436 28086 27488 28092
rect 27540 27538 27568 28426
rect 27632 27674 27660 28494
rect 27724 28082 27752 28494
rect 27816 28234 27844 29174
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 27816 28206 27936 28234
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27804 28076 27856 28082
rect 27804 28018 27856 28024
rect 27620 27668 27672 27674
rect 27620 27610 27672 27616
rect 27528 27532 27580 27538
rect 27528 27474 27580 27480
rect 27816 26858 27844 28018
rect 27908 26926 27936 28206
rect 28092 28064 28120 29106
rect 28172 29028 28224 29034
rect 28172 28970 28224 28976
rect 28184 28665 28212 28970
rect 28170 28656 28226 28665
rect 28170 28591 28226 28600
rect 28172 28076 28224 28082
rect 28092 28036 28172 28064
rect 28172 28018 28224 28024
rect 28368 26994 28396 31350
rect 28736 30802 28764 31894
rect 28828 31822 28856 32438
rect 29184 32224 29236 32230
rect 29184 32166 29236 32172
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 29000 31816 29052 31822
rect 29000 31758 29052 31764
rect 28828 31686 28856 31758
rect 29012 31686 29040 31758
rect 29196 31754 29224 32166
rect 29184 31748 29236 31754
rect 29184 31690 29236 31696
rect 28816 31680 28868 31686
rect 28816 31622 28868 31628
rect 29000 31680 29052 31686
rect 29000 31622 29052 31628
rect 29012 31464 29040 31622
rect 28828 31436 29040 31464
rect 28828 31346 28856 31436
rect 29196 31414 29224 31690
rect 29184 31408 29236 31414
rect 29184 31350 29236 31356
rect 29460 31408 29512 31414
rect 29460 31350 29512 31356
rect 28816 31340 28868 31346
rect 28816 31282 28868 31288
rect 28724 30796 28776 30802
rect 28724 30738 28776 30744
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28540 29640 28592 29646
rect 28540 29582 28592 29588
rect 28552 29238 28580 29582
rect 28644 29238 28672 30602
rect 29000 29572 29052 29578
rect 29000 29514 29052 29520
rect 28540 29232 28592 29238
rect 28632 29232 28684 29238
rect 28540 29174 28592 29180
rect 28630 29200 28632 29209
rect 28684 29200 28686 29209
rect 28630 29135 28686 29144
rect 28724 28620 28776 28626
rect 28724 28562 28776 28568
rect 28736 28218 28764 28562
rect 28816 28416 28868 28422
rect 28816 28358 28868 28364
rect 28448 28212 28500 28218
rect 28448 28154 28500 28160
rect 28724 28212 28776 28218
rect 28724 28154 28776 28160
rect 28460 28082 28488 28154
rect 28736 28098 28764 28154
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28552 28070 28764 28098
rect 28552 28014 28580 28070
rect 28540 28008 28592 28014
rect 28540 27950 28592 27956
rect 28632 27940 28684 27946
rect 28632 27882 28684 27888
rect 28644 27538 28672 27882
rect 28632 27532 28684 27538
rect 28632 27474 28684 27480
rect 28736 27010 28764 28070
rect 28828 27470 28856 28358
rect 28906 27976 28962 27985
rect 28906 27911 28962 27920
rect 28816 27464 28868 27470
rect 28816 27406 28868 27412
rect 28356 26988 28408 26994
rect 28736 26982 28856 27010
rect 28920 26994 28948 27911
rect 29012 27169 29040 29514
rect 29184 29300 29236 29306
rect 29184 29242 29236 29248
rect 29092 27940 29144 27946
rect 29092 27882 29144 27888
rect 28998 27160 29054 27169
rect 28998 27095 29054 27104
rect 29104 27010 29132 27882
rect 29196 27606 29224 29242
rect 29276 28756 29328 28762
rect 29276 28698 29328 28704
rect 29184 27600 29236 27606
rect 29184 27542 29236 27548
rect 29288 27538 29316 28698
rect 29472 28082 29500 31350
rect 29552 31340 29604 31346
rect 29552 31282 29604 31288
rect 29564 30938 29592 31282
rect 29552 30932 29604 30938
rect 29552 30874 29604 30880
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29748 29034 29776 29582
rect 29736 29028 29788 29034
rect 29736 28970 29788 28976
rect 29840 28762 29868 29582
rect 29828 28756 29880 28762
rect 29828 28698 29880 28704
rect 29932 28558 29960 36518
rect 30472 36372 30524 36378
rect 30472 36314 30524 36320
rect 30104 36304 30156 36310
rect 30104 36246 30156 36252
rect 30116 36174 30144 36246
rect 30104 36168 30156 36174
rect 30104 36110 30156 36116
rect 30012 34536 30064 34542
rect 30012 34478 30064 34484
rect 30024 33658 30052 34478
rect 30012 33652 30064 33658
rect 30012 33594 30064 33600
rect 30116 33538 30144 36110
rect 30484 36106 30512 36314
rect 30576 36122 30604 39238
rect 30748 37732 30800 37738
rect 30748 37674 30800 37680
rect 30656 37256 30708 37262
rect 30656 37198 30708 37204
rect 30668 36786 30696 37198
rect 30656 36780 30708 36786
rect 30656 36722 30708 36728
rect 30668 36378 30696 36722
rect 30656 36372 30708 36378
rect 30656 36314 30708 36320
rect 30472 36100 30524 36106
rect 30576 36094 30696 36122
rect 30472 36042 30524 36048
rect 30484 35834 30512 36042
rect 30472 35828 30524 35834
rect 30472 35770 30524 35776
rect 30196 35556 30248 35562
rect 30196 35498 30248 35504
rect 30208 34202 30236 35498
rect 30288 35012 30340 35018
rect 30288 34954 30340 34960
rect 30300 34678 30328 34954
rect 30288 34672 30340 34678
rect 30288 34614 30340 34620
rect 30196 34196 30248 34202
rect 30196 34138 30248 34144
rect 30024 33510 30144 33538
rect 30024 30784 30052 33510
rect 30668 32910 30696 36094
rect 30760 34542 30788 37674
rect 30748 34536 30800 34542
rect 30748 34478 30800 34484
rect 30852 34066 30880 39442
rect 30932 39364 30984 39370
rect 30932 39306 30984 39312
rect 30840 34060 30892 34066
rect 30840 34002 30892 34008
rect 30656 32904 30708 32910
rect 30656 32846 30708 32852
rect 30104 32768 30156 32774
rect 30104 32710 30156 32716
rect 30116 32502 30144 32710
rect 30104 32496 30156 32502
rect 30104 32438 30156 32444
rect 30196 32428 30248 32434
rect 30196 32370 30248 32376
rect 30208 31414 30236 32370
rect 30288 32292 30340 32298
rect 30288 32234 30340 32240
rect 30300 31754 30328 32234
rect 30668 32230 30696 32846
rect 30656 32224 30708 32230
rect 30656 32166 30708 32172
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30288 31748 30340 31754
rect 30288 31690 30340 31696
rect 30196 31408 30248 31414
rect 30196 31350 30248 31356
rect 30300 31210 30328 31690
rect 30392 31482 30420 31758
rect 30380 31476 30432 31482
rect 30380 31418 30432 31424
rect 30288 31204 30340 31210
rect 30288 31146 30340 31152
rect 30300 30802 30328 31146
rect 30944 31142 30972 39306
rect 31128 38758 31156 39510
rect 31496 39506 31524 40666
rect 31484 39500 31536 39506
rect 31484 39442 31536 39448
rect 31392 38956 31444 38962
rect 31392 38898 31444 38904
rect 31116 38752 31168 38758
rect 31116 38694 31168 38700
rect 31116 37256 31168 37262
rect 31116 37198 31168 37204
rect 31208 37256 31260 37262
rect 31208 37198 31260 37204
rect 31128 36786 31156 37198
rect 31116 36780 31168 36786
rect 31116 36722 31168 36728
rect 31128 36378 31156 36722
rect 31220 36650 31248 37198
rect 31300 37120 31352 37126
rect 31300 37062 31352 37068
rect 31312 36718 31340 37062
rect 31404 36922 31432 38898
rect 31484 37256 31536 37262
rect 31484 37198 31536 37204
rect 31392 36916 31444 36922
rect 31392 36858 31444 36864
rect 31496 36854 31524 37198
rect 31576 37120 31628 37126
rect 31576 37062 31628 37068
rect 31484 36848 31536 36854
rect 31482 36816 31484 36825
rect 31536 36816 31538 36825
rect 31588 36786 31616 37062
rect 31482 36751 31538 36760
rect 31576 36780 31628 36786
rect 31576 36722 31628 36728
rect 31300 36712 31352 36718
rect 31300 36654 31352 36660
rect 31208 36644 31260 36650
rect 31208 36586 31260 36592
rect 31116 36372 31168 36378
rect 31116 36314 31168 36320
rect 31024 36168 31076 36174
rect 31024 36110 31076 36116
rect 31208 36168 31260 36174
rect 31208 36110 31260 36116
rect 31036 35630 31064 36110
rect 31220 36038 31248 36110
rect 31680 36106 31708 40854
rect 31772 40594 31800 41074
rect 31760 40588 31812 40594
rect 31760 40530 31812 40536
rect 31758 40080 31814 40089
rect 31758 40015 31814 40024
rect 32036 40044 32088 40050
rect 31772 37194 31800 40015
rect 32036 39986 32088 39992
rect 32048 39642 32076 39986
rect 32036 39636 32088 39642
rect 32036 39578 32088 39584
rect 32048 39506 32076 39578
rect 32036 39500 32088 39506
rect 32036 39442 32088 39448
rect 31852 39432 31904 39438
rect 31852 39374 31904 39380
rect 31864 38894 31892 39374
rect 31944 39364 31996 39370
rect 31944 39306 31996 39312
rect 31956 39098 31984 39306
rect 32140 39098 32168 42638
rect 33152 42362 33180 42842
rect 33508 42696 33560 42702
rect 33508 42638 33560 42644
rect 33232 42560 33284 42566
rect 33232 42502 33284 42508
rect 33140 42356 33192 42362
rect 33140 42298 33192 42304
rect 32864 41676 32916 41682
rect 32864 41618 32916 41624
rect 32772 41472 32824 41478
rect 32772 41414 32824 41420
rect 32588 40928 32640 40934
rect 32588 40870 32640 40876
rect 32404 40384 32456 40390
rect 32404 40326 32456 40332
rect 32416 40118 32444 40326
rect 32404 40112 32456 40118
rect 32404 40054 32456 40060
rect 32416 39930 32444 40054
rect 32324 39902 32444 39930
rect 32496 39908 32548 39914
rect 32220 39636 32272 39642
rect 32220 39578 32272 39584
rect 32232 39438 32260 39578
rect 32324 39438 32352 39902
rect 32496 39850 32548 39856
rect 32404 39840 32456 39846
rect 32404 39782 32456 39788
rect 32220 39432 32272 39438
rect 32220 39374 32272 39380
rect 32312 39432 32364 39438
rect 32312 39374 32364 39380
rect 32220 39296 32272 39302
rect 32220 39238 32272 39244
rect 31944 39092 31996 39098
rect 31944 39034 31996 39040
rect 32128 39092 32180 39098
rect 32128 39034 32180 39040
rect 32140 38962 32168 39034
rect 32128 38956 32180 38962
rect 32128 38898 32180 38904
rect 31852 38888 31904 38894
rect 31852 38830 31904 38836
rect 32128 38820 32180 38826
rect 32128 38762 32180 38768
rect 31944 38752 31996 38758
rect 31944 38694 31996 38700
rect 31852 38548 31904 38554
rect 31852 38490 31904 38496
rect 31760 37188 31812 37194
rect 31760 37130 31812 37136
rect 31758 36136 31814 36145
rect 31484 36100 31536 36106
rect 31484 36042 31536 36048
rect 31668 36100 31720 36106
rect 31864 36122 31892 38490
rect 31956 38214 31984 38694
rect 32140 38554 32168 38762
rect 32128 38548 32180 38554
rect 32128 38490 32180 38496
rect 32232 38418 32260 39238
rect 32220 38412 32272 38418
rect 32220 38354 32272 38360
rect 32416 38350 32444 39782
rect 32508 39522 32536 39850
rect 32600 39642 32628 40870
rect 32784 40526 32812 41414
rect 32876 41206 32904 41618
rect 33244 41614 33272 42502
rect 33324 41676 33376 41682
rect 33324 41618 33376 41624
rect 33232 41608 33284 41614
rect 33232 41550 33284 41556
rect 32864 41200 32916 41206
rect 32864 41142 32916 41148
rect 33244 41138 33272 41550
rect 33140 41132 33192 41138
rect 33140 41074 33192 41080
rect 33232 41132 33284 41138
rect 33232 41074 33284 41080
rect 33048 41064 33100 41070
rect 33048 41006 33100 41012
rect 33060 40662 33088 41006
rect 33048 40656 33100 40662
rect 33048 40598 33100 40604
rect 32864 40588 32916 40594
rect 32864 40530 32916 40536
rect 32772 40520 32824 40526
rect 32772 40462 32824 40468
rect 32876 40186 32904 40530
rect 32864 40180 32916 40186
rect 32864 40122 32916 40128
rect 33152 40118 33180 41074
rect 33244 40526 33272 41074
rect 33336 41002 33364 41618
rect 33416 41540 33468 41546
rect 33416 41482 33468 41488
rect 33428 41138 33456 41482
rect 33416 41132 33468 41138
rect 33416 41074 33468 41080
rect 33324 40996 33376 41002
rect 33324 40938 33376 40944
rect 33428 40526 33456 41074
rect 33232 40520 33284 40526
rect 33232 40462 33284 40468
rect 33416 40520 33468 40526
rect 33416 40462 33468 40468
rect 33140 40112 33192 40118
rect 33140 40054 33192 40060
rect 32680 39840 32732 39846
rect 32680 39782 32732 39788
rect 32588 39636 32640 39642
rect 32588 39578 32640 39584
rect 32508 39494 32628 39522
rect 32692 39506 32720 39782
rect 33520 39642 33548 42638
rect 33796 42362 33824 43046
rect 33888 42906 33916 43182
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 33876 42900 33928 42906
rect 33876 42842 33928 42848
rect 33784 42356 33836 42362
rect 33784 42298 33836 42304
rect 33888 42226 33916 42842
rect 34336 42764 34388 42770
rect 34336 42706 34388 42712
rect 33968 42696 34020 42702
rect 33968 42638 34020 42644
rect 33980 42362 34008 42638
rect 34060 42628 34112 42634
rect 34060 42570 34112 42576
rect 34152 42628 34204 42634
rect 34152 42570 34204 42576
rect 33968 42356 34020 42362
rect 33968 42298 34020 42304
rect 33876 42220 33928 42226
rect 33876 42162 33928 42168
rect 33600 42152 33652 42158
rect 33600 42094 33652 42100
rect 33612 41274 33640 42094
rect 33888 41682 33916 42162
rect 33876 41676 33928 41682
rect 33876 41618 33928 41624
rect 33980 41546 34008 42298
rect 34072 41818 34100 42570
rect 34164 42294 34192 42570
rect 34152 42288 34204 42294
rect 34152 42230 34204 42236
rect 34060 41812 34112 41818
rect 34060 41754 34112 41760
rect 34164 41614 34192 42230
rect 34348 42226 34376 42706
rect 35348 42560 35400 42566
rect 35348 42502 35400 42508
rect 34336 42220 34388 42226
rect 34336 42162 34388 42168
rect 34704 42152 34756 42158
rect 34704 42094 34756 42100
rect 34716 41818 34744 42094
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34704 41812 34756 41818
rect 34704 41754 34756 41760
rect 34428 41744 34480 41750
rect 34428 41686 34480 41692
rect 34152 41608 34204 41614
rect 34152 41550 34204 41556
rect 33968 41540 34020 41546
rect 33968 41482 34020 41488
rect 33600 41268 33652 41274
rect 33600 41210 33652 41216
rect 34440 41070 34468 41686
rect 35360 41546 35388 42502
rect 35594 42460 35902 42469
rect 35594 42458 35600 42460
rect 35656 42458 35680 42460
rect 35736 42458 35760 42460
rect 35816 42458 35840 42460
rect 35896 42458 35902 42460
rect 35656 42406 35658 42458
rect 35838 42406 35840 42458
rect 35594 42404 35600 42406
rect 35656 42404 35680 42406
rect 35736 42404 35760 42406
rect 35816 42404 35840 42406
rect 35896 42404 35902 42406
rect 35594 42395 35902 42404
rect 37464 42152 37516 42158
rect 37464 42094 37516 42100
rect 38568 42152 38620 42158
rect 38568 42094 38620 42100
rect 35992 42084 36044 42090
rect 35992 42026 36044 42032
rect 35348 41540 35400 41546
rect 35348 41482 35400 41488
rect 35164 41472 35216 41478
rect 35164 41414 35216 41420
rect 35176 41274 35204 41414
rect 35594 41372 35902 41381
rect 35594 41370 35600 41372
rect 35656 41370 35680 41372
rect 35736 41370 35760 41372
rect 35816 41370 35840 41372
rect 35896 41370 35902 41372
rect 35656 41318 35658 41370
rect 35838 41318 35840 41370
rect 35594 41316 35600 41318
rect 35656 41316 35680 41318
rect 35736 41316 35760 41318
rect 35816 41316 35840 41318
rect 35896 41316 35902 41318
rect 35594 41307 35902 41316
rect 35164 41268 35216 41274
rect 35164 41210 35216 41216
rect 34796 41200 34848 41206
rect 34796 41142 34848 41148
rect 34428 41064 34480 41070
rect 34428 41006 34480 41012
rect 34704 40996 34756 41002
rect 34704 40938 34756 40944
rect 34716 40730 34744 40938
rect 34704 40724 34756 40730
rect 34704 40666 34756 40672
rect 33508 39636 33560 39642
rect 33508 39578 33560 39584
rect 32600 39438 32628 39494
rect 32680 39500 32732 39506
rect 32680 39442 32732 39448
rect 32588 39432 32640 39438
rect 32588 39374 32640 39380
rect 32404 38344 32456 38350
rect 32404 38286 32456 38292
rect 32600 38214 32628 39374
rect 32692 38418 32720 39442
rect 33520 38962 33548 39578
rect 34612 39568 34664 39574
rect 34532 39516 34612 39522
rect 34808 39522 34836 41142
rect 35440 41132 35492 41138
rect 35440 41074 35492 41080
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35348 39840 35400 39846
rect 35348 39782 35400 39788
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34888 39636 34940 39642
rect 34888 39578 34940 39584
rect 35256 39636 35308 39642
rect 35256 39578 35308 39584
rect 34532 39510 34664 39516
rect 34532 39494 34652 39510
rect 34716 39494 34836 39522
rect 34244 39432 34296 39438
rect 34244 39374 34296 39380
rect 33968 39092 34020 39098
rect 33968 39034 34020 39040
rect 33980 38962 34008 39034
rect 33508 38956 33560 38962
rect 33508 38898 33560 38904
rect 33968 38956 34020 38962
rect 33968 38898 34020 38904
rect 32680 38412 32732 38418
rect 32680 38354 32732 38360
rect 31944 38208 31996 38214
rect 31944 38150 31996 38156
rect 32588 38208 32640 38214
rect 32588 38150 32640 38156
rect 32036 37324 32088 37330
rect 32036 37266 32088 37272
rect 32048 36922 32076 37266
rect 32772 37188 32824 37194
rect 32772 37130 32824 37136
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32036 36916 32088 36922
rect 32036 36858 32088 36864
rect 32128 36780 32180 36786
rect 32128 36722 32180 36728
rect 31814 36094 31892 36122
rect 31758 36071 31814 36080
rect 31668 36042 31720 36048
rect 31208 36032 31260 36038
rect 31208 35974 31260 35980
rect 31024 35624 31076 35630
rect 31024 35566 31076 35572
rect 31036 35290 31064 35566
rect 31024 35284 31076 35290
rect 31024 35226 31076 35232
rect 31496 35154 31524 36042
rect 31680 35834 31708 36042
rect 31668 35828 31720 35834
rect 31668 35770 31720 35776
rect 31772 35766 31800 36071
rect 31760 35760 31812 35766
rect 31760 35702 31812 35708
rect 32140 35170 32168 36722
rect 32404 36712 32456 36718
rect 32404 36654 32456 36660
rect 32416 36378 32444 36654
rect 32404 36372 32456 36378
rect 32404 36314 32456 36320
rect 32508 36242 32536 37062
rect 32496 36236 32548 36242
rect 32496 36178 32548 36184
rect 32404 35488 32456 35494
rect 32404 35430 32456 35436
rect 32048 35154 32168 35170
rect 32416 35154 32444 35430
rect 31484 35148 31536 35154
rect 31484 35090 31536 35096
rect 32048 35148 32180 35154
rect 32048 35142 32128 35148
rect 31392 34944 31444 34950
rect 31392 34886 31444 34892
rect 31300 34604 31352 34610
rect 31300 34546 31352 34552
rect 31116 34468 31168 34474
rect 31116 34410 31168 34416
rect 31128 33998 31156 34410
rect 31116 33992 31168 33998
rect 31116 33934 31168 33940
rect 31024 32224 31076 32230
rect 31024 32166 31076 32172
rect 31036 31482 31064 32166
rect 31024 31476 31076 31482
rect 31024 31418 31076 31424
rect 30932 31136 30984 31142
rect 30932 31078 30984 31084
rect 30944 30802 30972 31078
rect 30288 30796 30340 30802
rect 30024 30756 30236 30784
rect 30104 30660 30156 30666
rect 30104 30602 30156 30608
rect 30116 29646 30144 30602
rect 30104 29640 30156 29646
rect 30104 29582 30156 29588
rect 30116 29170 30144 29582
rect 30104 29164 30156 29170
rect 30104 29106 30156 29112
rect 30116 28626 30144 29106
rect 30104 28620 30156 28626
rect 30104 28562 30156 28568
rect 29644 28552 29696 28558
rect 29564 28512 29644 28540
rect 29564 28150 29592 28512
rect 29644 28494 29696 28500
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 30012 28552 30064 28558
rect 30012 28494 30064 28500
rect 29932 28150 29960 28494
rect 29552 28144 29604 28150
rect 29552 28086 29604 28092
rect 29920 28144 29972 28150
rect 29920 28086 29972 28092
rect 29460 28076 29512 28082
rect 29460 28018 29512 28024
rect 29276 27532 29328 27538
rect 29276 27474 29328 27480
rect 29184 27464 29236 27470
rect 29184 27406 29236 27412
rect 29196 27130 29224 27406
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 29012 26994 29132 27010
rect 28356 26930 28408 26936
rect 27896 26920 27948 26926
rect 27896 26862 27948 26868
rect 27804 26852 27856 26858
rect 27804 26794 27856 26800
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 27436 25152 27488 25158
rect 27436 25094 27488 25100
rect 27448 24886 27476 25094
rect 27436 24880 27488 24886
rect 27436 24822 27488 24828
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27540 24154 27568 24754
rect 27632 24274 27660 25774
rect 27816 24886 27844 26794
rect 27908 26518 27936 26862
rect 27896 26512 27948 26518
rect 27896 26454 27948 26460
rect 27896 25832 27948 25838
rect 27896 25774 27948 25780
rect 27908 25498 27936 25774
rect 27896 25492 27948 25498
rect 27896 25434 27948 25440
rect 27804 24880 27856 24886
rect 27804 24822 27856 24828
rect 27712 24812 27764 24818
rect 27712 24754 27764 24760
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 27724 24614 27752 24754
rect 27712 24608 27764 24614
rect 27712 24550 27764 24556
rect 27804 24608 27856 24614
rect 28000 24585 28028 24754
rect 28172 24676 28224 24682
rect 28172 24618 28224 24624
rect 27804 24550 27856 24556
rect 27986 24576 28042 24585
rect 27620 24268 27672 24274
rect 27672 24228 27752 24256
rect 27620 24210 27672 24216
rect 27540 24126 27660 24154
rect 27344 23792 27396 23798
rect 27344 23734 27396 23740
rect 27436 23792 27488 23798
rect 27436 23734 27488 23740
rect 27252 23588 27304 23594
rect 27252 23530 27304 23536
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 27172 22642 27200 22918
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 26988 22094 27016 22510
rect 27172 22094 27200 22578
rect 27448 22094 27476 23734
rect 27632 22094 27660 24126
rect 27724 23118 27752 24228
rect 27816 23730 27844 24550
rect 27986 24511 28042 24520
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27908 23662 27936 24346
rect 28184 24274 28212 24618
rect 28368 24410 28396 26930
rect 28828 26926 28856 26982
rect 28908 26988 28960 26994
rect 28908 26930 28960 26936
rect 29000 26988 29132 26994
rect 29052 26982 29132 26988
rect 29000 26930 29052 26936
rect 28816 26920 28868 26926
rect 28816 26862 28868 26868
rect 28724 26784 28776 26790
rect 28724 26726 28776 26732
rect 28448 25832 28500 25838
rect 28448 25774 28500 25780
rect 28356 24404 28408 24410
rect 28356 24346 28408 24352
rect 28172 24268 28224 24274
rect 28172 24210 28224 24216
rect 28460 24206 28488 25774
rect 28540 25152 28592 25158
rect 28540 25094 28592 25100
rect 28632 25152 28684 25158
rect 28632 25094 28684 25100
rect 28552 24834 28580 25094
rect 28644 24954 28672 25094
rect 28632 24948 28684 24954
rect 28632 24890 28684 24896
rect 28552 24818 28672 24834
rect 28552 24812 28684 24818
rect 28552 24806 28632 24812
rect 28632 24754 28684 24760
rect 28644 24342 28672 24754
rect 28632 24336 28684 24342
rect 28632 24278 28684 24284
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 27988 23792 28040 23798
rect 27988 23734 28040 23740
rect 27896 23656 27948 23662
rect 27896 23598 27948 23604
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27724 22642 27752 23054
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27908 22166 27936 22646
rect 27896 22160 27948 22166
rect 27896 22102 27948 22108
rect 26620 22066 26832 22094
rect 26988 22066 27108 22094
rect 27172 22066 27292 22094
rect 27448 22066 27568 22094
rect 27632 22066 27752 22094
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 26620 21486 26648 21830
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 26516 19304 26568 19310
rect 26516 19246 26568 19252
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 25976 17224 26188 17252
rect 25792 16782 25912 16810
rect 25884 16726 25912 16782
rect 25872 16720 25924 16726
rect 25872 16662 25924 16668
rect 25872 15020 25924 15026
rect 25872 14962 25924 14968
rect 25884 14822 25912 14962
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25700 14074 25820 14090
rect 25596 14068 25648 14074
rect 25700 14068 25832 14074
rect 25700 14062 25780 14068
rect 25596 14010 25648 14016
rect 25780 14010 25832 14016
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25608 13394 25636 13874
rect 25884 13870 25912 14758
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25596 13388 25648 13394
rect 25596 13330 25648 13336
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25516 10062 25544 11494
rect 25504 10056 25556 10062
rect 25504 9998 25556 10004
rect 25516 9722 25544 9998
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 25700 9654 25728 13806
rect 25884 13258 25912 13806
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25872 12300 25924 12306
rect 25872 12242 25924 12248
rect 25780 12232 25832 12238
rect 25780 12174 25832 12180
rect 25792 11830 25820 12174
rect 25780 11824 25832 11830
rect 25780 11766 25832 11772
rect 25884 10606 25912 12242
rect 25976 10810 26004 17224
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 26068 16590 26096 17070
rect 26056 16584 26108 16590
rect 26056 16526 26108 16532
rect 26148 16516 26200 16522
rect 26148 16458 26200 16464
rect 26056 15564 26108 15570
rect 26056 15506 26108 15512
rect 26068 15434 26096 15506
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 26160 14906 26188 16458
rect 26424 15904 26476 15910
rect 26424 15846 26476 15852
rect 26332 15632 26384 15638
rect 26332 15574 26384 15580
rect 26344 15434 26372 15574
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26238 15192 26294 15201
rect 26238 15127 26294 15136
rect 26252 15094 26280 15127
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 26436 15026 26464 15846
rect 26528 15570 26556 17818
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26528 15434 26556 15506
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26160 14878 26280 14906
rect 26252 14822 26280 14878
rect 26424 14884 26476 14890
rect 26424 14826 26476 14832
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26056 13796 26108 13802
rect 26056 13738 26108 13744
rect 26068 13258 26096 13738
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 26160 12238 26188 12854
rect 26436 12442 26464 14826
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 26056 12232 26108 12238
rect 26056 12174 26108 12180
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26068 11558 26096 12174
rect 26160 11898 26188 12174
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 26160 10130 26188 11834
rect 26332 11824 26384 11830
rect 26332 11766 26384 11772
rect 26344 11150 26372 11766
rect 26436 11370 26464 12378
rect 26528 12170 26556 14282
rect 26516 12164 26568 12170
rect 26516 12106 26568 12112
rect 26620 11694 26648 21422
rect 26804 19514 26832 22066
rect 26976 21956 27028 21962
rect 26976 21898 27028 21904
rect 26988 21554 27016 21898
rect 27080 21894 27108 22066
rect 27068 21888 27120 21894
rect 27068 21830 27120 21836
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 26988 20942 27016 21490
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 26976 20324 27028 20330
rect 26976 20266 27028 20272
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26896 19786 26924 20198
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 26792 19508 26844 19514
rect 26792 19450 26844 19456
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 26712 18970 26740 19246
rect 26700 18964 26752 18970
rect 26700 18906 26752 18912
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26804 15366 26832 15914
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26712 14278 26740 15302
rect 26792 14884 26844 14890
rect 26792 14826 26844 14832
rect 26804 14414 26832 14826
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26896 14346 26924 16594
rect 26884 14340 26936 14346
rect 26884 14282 26936 14288
rect 26700 14272 26752 14278
rect 26988 14226 27016 20266
rect 26700 14214 26752 14220
rect 26712 13938 26740 14214
rect 26804 14198 27016 14226
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 26804 12434 26832 14198
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 26896 13462 26924 14010
rect 26976 13728 27028 13734
rect 26976 13670 27028 13676
rect 26884 13456 26936 13462
rect 26884 13398 26936 13404
rect 26988 13190 27016 13670
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 26976 12436 27028 12442
rect 26804 12406 26924 12434
rect 26608 11688 26660 11694
rect 26608 11630 26660 11636
rect 26436 11342 26556 11370
rect 26528 11286 26556 11342
rect 26516 11280 26568 11286
rect 26516 11222 26568 11228
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26332 11144 26384 11150
rect 26332 11086 26384 11092
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 25412 9444 25464 9450
rect 25412 9386 25464 9392
rect 25424 9042 25452 9386
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25700 8974 25728 9590
rect 25688 8968 25740 8974
rect 25608 8928 25688 8956
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25424 8498 25452 8570
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 24952 7744 25004 7750
rect 24952 7686 25004 7692
rect 24308 7472 24360 7478
rect 24308 7414 24360 7420
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24768 7472 24820 7478
rect 24768 7414 24820 7420
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24504 6798 24532 7346
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 24216 6724 24268 6730
rect 24216 6666 24268 6672
rect 23756 5772 23808 5778
rect 23756 5714 23808 5720
rect 24228 5710 24256 6666
rect 24964 6662 24992 7686
rect 25412 7200 25464 7206
rect 25412 7142 25464 7148
rect 25424 7002 25452 7142
rect 25412 6996 25464 7002
rect 25412 6938 25464 6944
rect 25608 6730 25636 8928
rect 25688 8910 25740 8916
rect 26344 8498 26372 10406
rect 26436 9042 26464 11154
rect 26516 10464 26568 10470
rect 26516 10406 26568 10412
rect 26528 10130 26556 10406
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26620 9994 26648 11154
rect 26792 11008 26844 11014
rect 26792 10950 26844 10956
rect 26804 10742 26832 10950
rect 26896 10742 26924 12406
rect 26976 12378 27028 12384
rect 26988 11762 27016 12378
rect 27080 11762 27108 21830
rect 27264 17252 27292 22066
rect 27540 21554 27568 22066
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27632 20330 27660 20742
rect 27724 20602 27752 22066
rect 27896 21072 27948 21078
rect 27896 21014 27948 21020
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27620 20324 27672 20330
rect 27620 20266 27672 20272
rect 27724 19718 27752 20538
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27528 18216 27580 18222
rect 27528 18158 27580 18164
rect 27540 17882 27568 18158
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27356 17338 27384 17546
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 27172 17224 27292 17252
rect 27172 12434 27200 17224
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27264 16182 27292 16390
rect 27252 16176 27304 16182
rect 27252 16118 27304 16124
rect 27448 15638 27476 17138
rect 27632 15910 27660 17478
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 27620 15904 27672 15910
rect 27620 15846 27672 15852
rect 27436 15632 27488 15638
rect 27436 15574 27488 15580
rect 27632 15502 27660 15846
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 27264 15337 27292 15370
rect 27528 15360 27580 15366
rect 27250 15328 27306 15337
rect 27528 15302 27580 15308
rect 27250 15263 27306 15272
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27252 14816 27304 14822
rect 27252 14758 27304 14764
rect 27264 13258 27292 14758
rect 27448 14074 27476 14962
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27252 13252 27304 13258
rect 27252 13194 27304 13200
rect 27448 12866 27476 14010
rect 27540 13326 27568 15302
rect 27632 15094 27660 15438
rect 27724 15434 27752 17138
rect 27804 16992 27856 16998
rect 27804 16934 27856 16940
rect 27816 16046 27844 16934
rect 27804 16040 27856 16046
rect 27804 15982 27856 15988
rect 27908 15858 27936 21014
rect 28000 16726 28028 23734
rect 28080 23656 28132 23662
rect 28080 23598 28132 23604
rect 28356 23656 28408 23662
rect 28356 23598 28408 23604
rect 28092 22506 28120 23598
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 28080 22500 28132 22506
rect 28080 22442 28132 22448
rect 28184 21962 28212 22578
rect 28172 21956 28224 21962
rect 28172 21898 28224 21904
rect 28368 21690 28396 23598
rect 28540 22432 28592 22438
rect 28540 22374 28592 22380
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28356 21684 28408 21690
rect 28356 21626 28408 21632
rect 28460 21486 28488 21898
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 28460 21078 28488 21422
rect 28448 21072 28500 21078
rect 28368 21020 28448 21026
rect 28368 21014 28500 21020
rect 28368 20998 28488 21014
rect 28368 20466 28396 20998
rect 28552 20942 28580 22374
rect 28644 22094 28672 24278
rect 28736 23730 28764 26726
rect 28920 26518 28948 26930
rect 28908 26512 28960 26518
rect 28908 26454 28960 26460
rect 29288 26450 29316 27474
rect 29092 26444 29144 26450
rect 29092 26386 29144 26392
rect 29276 26444 29328 26450
rect 29276 26386 29328 26392
rect 28908 25696 28960 25702
rect 28908 25638 28960 25644
rect 28920 25362 28948 25638
rect 29104 25362 29132 26386
rect 29472 26042 29500 28018
rect 29460 26036 29512 26042
rect 29460 25978 29512 25984
rect 29276 25424 29328 25430
rect 29276 25366 29328 25372
rect 28908 25356 28960 25362
rect 28908 25298 28960 25304
rect 29092 25356 29144 25362
rect 29092 25298 29144 25304
rect 29092 25152 29144 25158
rect 29092 25094 29144 25100
rect 28816 24880 28868 24886
rect 28868 24828 29040 24834
rect 28816 24822 29040 24828
rect 28828 24806 29040 24822
rect 29104 24818 29132 25094
rect 29288 24818 29316 25366
rect 28908 24676 28960 24682
rect 28908 24618 28960 24624
rect 28816 24404 28868 24410
rect 28816 24346 28868 24352
rect 28828 24070 28856 24346
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 28736 23322 28764 23666
rect 28724 23316 28776 23322
rect 28724 23258 28776 23264
rect 28920 23118 28948 24618
rect 29012 23254 29040 24806
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29564 24750 29592 28086
rect 30024 28014 30052 28494
rect 30116 28218 30144 28562
rect 30104 28212 30156 28218
rect 30104 28154 30156 28160
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 30012 28008 30064 28014
rect 30012 27950 30064 27956
rect 29656 27130 29684 27950
rect 30208 27946 30236 30756
rect 30288 30738 30340 30744
rect 30932 30796 30984 30802
rect 30932 30738 30984 30744
rect 30472 30116 30524 30122
rect 30472 30058 30524 30064
rect 30484 29714 30512 30058
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30392 29238 30420 29582
rect 30484 29345 30512 29650
rect 31128 29646 31156 33934
rect 31208 31952 31260 31958
rect 31208 31894 31260 31900
rect 31220 30802 31248 31894
rect 31312 31754 31340 34546
rect 31404 33590 31432 34886
rect 31496 34746 31524 35090
rect 31484 34740 31536 34746
rect 31484 34682 31536 34688
rect 32048 34066 32076 35142
rect 32128 35090 32180 35096
rect 32404 35148 32456 35154
rect 32404 35090 32456 35096
rect 32128 34604 32180 34610
rect 32128 34546 32180 34552
rect 31668 34060 31720 34066
rect 31668 34002 31720 34008
rect 32036 34060 32088 34066
rect 32036 34002 32088 34008
rect 31576 33924 31628 33930
rect 31576 33866 31628 33872
rect 31484 33856 31536 33862
rect 31484 33798 31536 33804
rect 31496 33658 31524 33798
rect 31588 33658 31616 33866
rect 31484 33652 31536 33658
rect 31484 33594 31536 33600
rect 31576 33652 31628 33658
rect 31576 33594 31628 33600
rect 31392 33584 31444 33590
rect 31392 33526 31444 33532
rect 31496 32434 31524 33594
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31496 32026 31524 32370
rect 31484 32020 31536 32026
rect 31484 31962 31536 31968
rect 31588 31958 31616 33594
rect 31680 33454 31708 34002
rect 31668 33448 31720 33454
rect 31668 33390 31720 33396
rect 32036 32836 32088 32842
rect 32036 32778 32088 32784
rect 31576 31952 31628 31958
rect 31576 31894 31628 31900
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 31312 31726 31432 31754
rect 31208 30796 31260 30802
rect 31208 30738 31260 30744
rect 31024 29640 31076 29646
rect 31024 29582 31076 29588
rect 31116 29640 31168 29646
rect 31116 29582 31168 29588
rect 30564 29504 30616 29510
rect 30564 29446 30616 29452
rect 30470 29336 30526 29345
rect 30470 29271 30526 29280
rect 30380 29232 30432 29238
rect 30380 29174 30432 29180
rect 30576 29170 30604 29446
rect 31036 29306 31064 29582
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 31024 29300 31076 29306
rect 30944 29260 31024 29288
rect 30656 29232 30708 29238
rect 30656 29174 30708 29180
rect 30564 29164 30616 29170
rect 30564 29106 30616 29112
rect 30380 28960 30432 28966
rect 30380 28902 30432 28908
rect 30288 28552 30340 28558
rect 30288 28494 30340 28500
rect 30196 27940 30248 27946
rect 30196 27882 30248 27888
rect 30104 27872 30156 27878
rect 30104 27814 30156 27820
rect 29920 27532 29972 27538
rect 29920 27474 29972 27480
rect 29644 27124 29696 27130
rect 29644 27066 29696 27072
rect 29736 27056 29788 27062
rect 29736 26998 29788 27004
rect 29748 26382 29776 26998
rect 29932 26994 29960 27474
rect 30116 27441 30144 27814
rect 30102 27432 30158 27441
rect 30102 27367 30158 27376
rect 29920 26988 29972 26994
rect 29920 26930 29972 26936
rect 30012 26784 30064 26790
rect 30012 26726 30064 26732
rect 29736 26376 29788 26382
rect 29736 26318 29788 26324
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 29656 24886 29684 25978
rect 29736 25152 29788 25158
rect 29736 25094 29788 25100
rect 29644 24880 29696 24886
rect 29644 24822 29696 24828
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 29000 23248 29052 23254
rect 29000 23190 29052 23196
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 29092 23044 29144 23050
rect 29092 22986 29144 22992
rect 28644 22066 28764 22094
rect 28736 20942 28764 22066
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28828 21350 28856 21966
rect 29000 21956 29052 21962
rect 29000 21898 29052 21904
rect 28816 21344 28868 21350
rect 28816 21286 28868 21292
rect 28828 20942 28856 21286
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 29012 20602 29040 21898
rect 29104 21146 29132 22986
rect 29564 22094 29592 24686
rect 29656 24342 29684 24822
rect 29644 24336 29696 24342
rect 29644 24278 29696 24284
rect 29748 23594 29776 25094
rect 29828 24812 29880 24818
rect 29828 24754 29880 24760
rect 29840 24614 29868 24754
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 29840 24138 29868 24550
rect 30024 24177 30052 26726
rect 30010 24168 30066 24177
rect 29828 24132 29880 24138
rect 30010 24103 30066 24112
rect 29828 24074 29880 24080
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29564 22066 29684 22094
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29564 21622 29592 21830
rect 29552 21616 29604 21622
rect 29552 21558 29604 21564
rect 29092 21140 29144 21146
rect 29092 21082 29144 21088
rect 29092 20800 29144 20806
rect 29092 20742 29144 20748
rect 29000 20596 29052 20602
rect 29000 20538 29052 20544
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 28080 20392 28132 20398
rect 28080 20334 28132 20340
rect 28092 18834 28120 20334
rect 28368 19922 28396 20402
rect 29012 20058 29040 20538
rect 29104 20398 29132 20742
rect 29184 20528 29236 20534
rect 29184 20470 29236 20476
rect 29092 20392 29144 20398
rect 29092 20334 29144 20340
rect 29000 20052 29052 20058
rect 29000 19994 29052 20000
rect 28356 19916 28408 19922
rect 28356 19858 28408 19864
rect 29196 19786 29224 20470
rect 29276 20256 29328 20262
rect 29276 20198 29328 20204
rect 29000 19780 29052 19786
rect 29000 19722 29052 19728
rect 29184 19780 29236 19786
rect 29184 19722 29236 19728
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 28264 19304 28316 19310
rect 28264 19246 28316 19252
rect 28276 18970 28304 19246
rect 28264 18964 28316 18970
rect 28264 18906 28316 18912
rect 28080 18828 28132 18834
rect 28080 18770 28132 18776
rect 28644 18290 28672 19450
rect 29012 19446 29040 19722
rect 29000 19440 29052 19446
rect 29052 19388 29132 19394
rect 29000 19382 29132 19388
rect 29012 19366 29132 19382
rect 29012 19310 29040 19366
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 28724 17536 28776 17542
rect 28724 17478 28776 17484
rect 28736 17202 28764 17478
rect 28920 17270 28948 18566
rect 29104 18358 29132 19366
rect 29092 18352 29144 18358
rect 29092 18294 29144 18300
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 29012 17338 29040 18158
rect 29104 17610 29132 18294
rect 29092 17604 29144 17610
rect 29092 17546 29144 17552
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 28908 17264 28960 17270
rect 28908 17206 28960 17212
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 28172 17196 28224 17202
rect 28172 17138 28224 17144
rect 28724 17196 28776 17202
rect 28724 17138 28776 17144
rect 28092 16794 28120 17138
rect 28080 16788 28132 16794
rect 28080 16730 28132 16736
rect 28184 16726 28212 17138
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 27988 16720 28040 16726
rect 27988 16662 28040 16668
rect 28172 16720 28224 16726
rect 28172 16662 28224 16668
rect 28540 16584 28592 16590
rect 28540 16526 28592 16532
rect 28552 15910 28580 16526
rect 29012 16250 29040 17070
rect 29104 16794 29132 17546
rect 29092 16788 29144 16794
rect 29092 16730 29144 16736
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 29104 16182 29132 16730
rect 29092 16176 29144 16182
rect 29092 16118 29144 16124
rect 29288 16130 29316 20198
rect 29656 19310 29684 22066
rect 30116 21962 30144 27367
rect 30196 26784 30248 26790
rect 30196 26726 30248 26732
rect 30208 26586 30236 26726
rect 30196 26580 30248 26586
rect 30196 26522 30248 26528
rect 30300 26382 30328 28494
rect 30392 28082 30420 28902
rect 30562 28792 30618 28801
rect 30668 28762 30696 29174
rect 30562 28727 30618 28736
rect 30656 28756 30708 28762
rect 30576 28694 30604 28727
rect 30656 28698 30708 28704
rect 30748 28756 30800 28762
rect 30748 28698 30800 28704
rect 30564 28688 30616 28694
rect 30564 28630 30616 28636
rect 30760 28626 30788 28698
rect 30748 28620 30800 28626
rect 30748 28562 30800 28568
rect 30472 28552 30524 28558
rect 30472 28494 30524 28500
rect 30484 28218 30512 28494
rect 30656 28484 30708 28490
rect 30656 28426 30708 28432
rect 30564 28416 30616 28422
rect 30564 28358 30616 28364
rect 30472 28212 30524 28218
rect 30472 28154 30524 28160
rect 30380 28076 30432 28082
rect 30380 28018 30432 28024
rect 30392 27985 30420 28018
rect 30378 27976 30434 27985
rect 30378 27911 30434 27920
rect 30576 27713 30604 28358
rect 30562 27704 30618 27713
rect 30562 27639 30618 27648
rect 30668 27606 30696 28426
rect 30656 27600 30708 27606
rect 30656 27542 30708 27548
rect 30668 27470 30696 27542
rect 30656 27464 30708 27470
rect 30656 27406 30708 27412
rect 30380 27328 30432 27334
rect 30380 27270 30432 27276
rect 30392 26382 30420 27270
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30668 26790 30696 26998
rect 30656 26784 30708 26790
rect 30656 26726 30708 26732
rect 30760 26382 30788 28562
rect 30944 28490 30972 29260
rect 31024 29242 31076 29248
rect 31312 29170 31340 29446
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 31116 29164 31168 29170
rect 31116 29106 31168 29112
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31036 28762 31064 29106
rect 31024 28756 31076 28762
rect 31024 28698 31076 28704
rect 31128 28626 31156 29106
rect 31208 28688 31260 28694
rect 31208 28630 31260 28636
rect 31116 28620 31168 28626
rect 31116 28562 31168 28568
rect 30932 28484 30984 28490
rect 30932 28426 30984 28432
rect 31128 28150 31156 28562
rect 31116 28144 31168 28150
rect 31116 28086 31168 28092
rect 31220 28082 31248 28630
rect 30840 28076 30892 28082
rect 30840 28018 30892 28024
rect 31208 28076 31260 28082
rect 31208 28018 31260 28024
rect 30852 27674 30880 28018
rect 31312 27962 31340 29106
rect 31128 27934 31340 27962
rect 30930 27704 30986 27713
rect 30840 27668 30892 27674
rect 30930 27639 30986 27648
rect 30840 27610 30892 27616
rect 30944 27470 30972 27639
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 30852 26450 30880 27406
rect 31024 27396 31076 27402
rect 31024 27338 31076 27344
rect 30840 26444 30892 26450
rect 30840 26386 30892 26392
rect 31036 26382 31064 27338
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 30380 26376 30432 26382
rect 30380 26318 30432 26324
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 31024 26376 31076 26382
rect 31024 26318 31076 26324
rect 30564 25696 30616 25702
rect 30564 25638 30616 25644
rect 30472 25424 30524 25430
rect 30472 25366 30524 25372
rect 30288 25288 30340 25294
rect 30288 25230 30340 25236
rect 30300 24954 30328 25230
rect 30288 24948 30340 24954
rect 30288 24890 30340 24896
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 30392 24410 30420 24686
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30484 24206 30512 25366
rect 30576 24410 30604 25638
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 30932 25288 30984 25294
rect 30932 25230 30984 25236
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30472 24200 30524 24206
rect 30472 24142 30524 24148
rect 30576 23186 30604 24346
rect 30668 24206 30696 25094
rect 30656 24200 30708 24206
rect 30656 24142 30708 24148
rect 30760 23866 30788 25230
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30852 24410 30880 25094
rect 30944 24614 30972 25230
rect 30932 24608 30984 24614
rect 30932 24550 30984 24556
rect 30840 24404 30892 24410
rect 30840 24346 30892 24352
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 30852 24070 30880 24142
rect 30944 24138 30972 24550
rect 30932 24132 30984 24138
rect 30932 24074 30984 24080
rect 31024 24132 31076 24138
rect 31024 24074 31076 24080
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30748 23860 30800 23866
rect 30748 23802 30800 23808
rect 30656 23724 30708 23730
rect 30852 23712 30880 24006
rect 31036 23730 31064 24074
rect 30708 23684 30880 23712
rect 31024 23724 31076 23730
rect 30656 23666 30708 23672
rect 31024 23666 31076 23672
rect 30564 23180 30616 23186
rect 30564 23122 30616 23128
rect 31128 23066 31156 27934
rect 31404 27520 31432 31726
rect 31668 31272 31720 31278
rect 31668 31214 31720 31220
rect 31680 30938 31708 31214
rect 31668 30932 31720 30938
rect 31668 30874 31720 30880
rect 31772 30802 31800 31758
rect 31944 31748 31996 31754
rect 31944 31690 31996 31696
rect 31956 31482 31984 31690
rect 32048 31482 32076 32778
rect 32140 32570 32168 34546
rect 32784 34542 32812 37130
rect 33520 36786 33548 38898
rect 33876 38752 33928 38758
rect 33876 38694 33928 38700
rect 33888 38593 33916 38694
rect 33874 38584 33930 38593
rect 33874 38519 33930 38528
rect 33888 38350 33916 38519
rect 33980 38418 34008 38898
rect 34256 38554 34284 39374
rect 34532 39370 34560 39494
rect 34520 39364 34572 39370
rect 34520 39306 34572 39312
rect 34336 39296 34388 39302
rect 34336 39238 34388 39244
rect 34428 39296 34480 39302
rect 34428 39238 34480 39244
rect 34244 38548 34296 38554
rect 34244 38490 34296 38496
rect 33968 38412 34020 38418
rect 33968 38354 34020 38360
rect 33876 38344 33928 38350
rect 33876 38286 33928 38292
rect 33980 37874 34008 38354
rect 34256 38350 34284 38490
rect 34244 38344 34296 38350
rect 34244 38286 34296 38292
rect 34348 38282 34376 39238
rect 34440 38758 34468 39238
rect 34428 38752 34480 38758
rect 34428 38694 34480 38700
rect 34532 38486 34560 39306
rect 34612 38888 34664 38894
rect 34612 38830 34664 38836
rect 34520 38480 34572 38486
rect 34520 38422 34572 38428
rect 34624 38282 34652 38830
rect 34336 38276 34388 38282
rect 34336 38218 34388 38224
rect 34612 38276 34664 38282
rect 34612 38218 34664 38224
rect 33968 37868 34020 37874
rect 33968 37810 34020 37816
rect 33600 37664 33652 37670
rect 33600 37606 33652 37612
rect 33508 36780 33560 36786
rect 33508 36722 33560 36728
rect 32864 36712 32916 36718
rect 32864 36654 32916 36660
rect 32772 34536 32824 34542
rect 32772 34478 32824 34484
rect 32588 32768 32640 32774
rect 32588 32710 32640 32716
rect 32128 32564 32180 32570
rect 32128 32506 32180 32512
rect 32600 31482 32628 32710
rect 32772 32360 32824 32366
rect 32772 32302 32824 32308
rect 32784 31822 32812 32302
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 31944 31476 31996 31482
rect 31944 31418 31996 31424
rect 32036 31476 32088 31482
rect 32036 31418 32088 31424
rect 32588 31476 32640 31482
rect 32588 31418 32640 31424
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32680 31340 32732 31346
rect 32680 31282 32732 31288
rect 31760 30796 31812 30802
rect 31760 30738 31812 30744
rect 31772 30258 31800 30738
rect 32312 30660 32364 30666
rect 32312 30602 32364 30608
rect 32324 30394 32352 30602
rect 32312 30388 32364 30394
rect 32312 30330 32364 30336
rect 31760 30252 31812 30258
rect 31760 30194 31812 30200
rect 31772 29782 31800 30194
rect 31484 29776 31536 29782
rect 31484 29718 31536 29724
rect 31668 29776 31720 29782
rect 31668 29718 31720 29724
rect 31760 29776 31812 29782
rect 31760 29718 31812 29724
rect 31496 29102 31524 29718
rect 31484 29096 31536 29102
rect 31484 29038 31536 29044
rect 31680 27538 31708 29718
rect 32416 29510 32444 31282
rect 32588 29844 32640 29850
rect 32588 29786 32640 29792
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 32036 29300 32088 29306
rect 32036 29242 32088 29248
rect 32048 28694 32076 29242
rect 32220 29164 32272 29170
rect 32220 29106 32272 29112
rect 32232 29073 32260 29106
rect 32218 29064 32274 29073
rect 32218 28999 32274 29008
rect 32036 28688 32088 28694
rect 32036 28630 32088 28636
rect 32048 28558 32076 28630
rect 31852 28552 31904 28558
rect 31852 28494 31904 28500
rect 32036 28552 32088 28558
rect 32036 28494 32088 28500
rect 31864 28014 31892 28494
rect 31852 28008 31904 28014
rect 31852 27950 31904 27956
rect 32128 27872 32180 27878
rect 32128 27814 32180 27820
rect 32140 27674 32168 27814
rect 32128 27668 32180 27674
rect 32128 27610 32180 27616
rect 31668 27532 31720 27538
rect 31404 27492 31524 27520
rect 31496 27402 31524 27492
rect 31668 27474 31720 27480
rect 31484 27396 31536 27402
rect 31484 27338 31536 27344
rect 31208 27328 31260 27334
rect 31208 27270 31260 27276
rect 31220 26790 31248 27270
rect 31208 26784 31260 26790
rect 31208 26726 31260 26732
rect 31496 26586 31524 27338
rect 32128 27124 32180 27130
rect 32128 27066 32180 27072
rect 31668 26784 31720 26790
rect 31668 26726 31720 26732
rect 31300 26580 31352 26586
rect 31300 26522 31352 26528
rect 31484 26580 31536 26586
rect 31484 26522 31536 26528
rect 31312 26228 31340 26522
rect 31484 26376 31536 26382
rect 31536 26336 31616 26364
rect 31484 26318 31536 26324
rect 31312 26200 31432 26228
rect 31404 25974 31432 26200
rect 31392 25968 31444 25974
rect 31392 25910 31444 25916
rect 31404 24886 31432 25910
rect 31588 25158 31616 26336
rect 31680 26246 31708 26726
rect 32140 26518 32168 27066
rect 31760 26512 31812 26518
rect 31760 26454 31812 26460
rect 31944 26512 31996 26518
rect 31944 26454 31996 26460
rect 32128 26512 32180 26518
rect 32128 26454 32180 26460
rect 31772 26382 31800 26454
rect 31760 26376 31812 26382
rect 31956 26353 31984 26454
rect 31760 26318 31812 26324
rect 31942 26344 31998 26353
rect 31942 26279 31998 26288
rect 31668 26240 31720 26246
rect 31668 26182 31720 26188
rect 31680 26042 31708 26182
rect 31668 26036 31720 26042
rect 31668 25978 31720 25984
rect 32140 25838 32168 26454
rect 32128 25832 32180 25838
rect 32128 25774 32180 25780
rect 31576 25152 31628 25158
rect 31576 25094 31628 25100
rect 31392 24880 31444 24886
rect 31392 24822 31444 24828
rect 31484 24608 31536 24614
rect 31484 24550 31536 24556
rect 31208 24200 31260 24206
rect 31392 24200 31444 24206
rect 31260 24160 31392 24188
rect 31208 24142 31260 24148
rect 31392 24142 31444 24148
rect 31300 23792 31352 23798
rect 31298 23760 31300 23769
rect 31352 23760 31354 23769
rect 31298 23695 31354 23704
rect 31312 23186 31340 23695
rect 31300 23180 31352 23186
rect 31300 23122 31352 23128
rect 31128 23038 31340 23066
rect 30288 22976 30340 22982
rect 30288 22918 30340 22924
rect 30300 22710 30328 22918
rect 30288 22704 30340 22710
rect 30288 22646 30340 22652
rect 31208 22092 31260 22098
rect 31208 22034 31260 22040
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30104 21956 30156 21962
rect 30104 21898 30156 21904
rect 29828 21888 29880 21894
rect 29828 21830 29880 21836
rect 29840 21010 29868 21830
rect 30944 21690 30972 21966
rect 31116 21888 31168 21894
rect 31116 21830 31168 21836
rect 30932 21684 30984 21690
rect 30932 21626 30984 21632
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 29920 21344 29972 21350
rect 29920 21286 29972 21292
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 29932 20942 29960 21286
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 30116 20398 30144 21422
rect 31128 20942 31156 21830
rect 31220 21350 31248 22034
rect 31208 21344 31260 21350
rect 31208 21286 31260 21292
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 30104 20392 30156 20398
rect 30156 20352 30236 20380
rect 30104 20334 30156 20340
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 29840 19514 29868 19654
rect 29828 19508 29880 19514
rect 29828 19450 29880 19456
rect 29840 19378 29868 19450
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29656 18766 29684 19246
rect 29644 18760 29696 18766
rect 29644 18702 29696 18708
rect 30208 17746 30236 20352
rect 31220 19496 31248 21286
rect 31128 19468 31248 19496
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30484 18970 30512 19246
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 31024 18828 31076 18834
rect 31024 18770 31076 18776
rect 30932 18624 30984 18630
rect 30932 18566 30984 18572
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 30484 17678 30512 18022
rect 30472 17672 30524 17678
rect 30472 17614 30524 17620
rect 29460 17536 29512 17542
rect 29460 17478 29512 17484
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30656 17536 30708 17542
rect 30656 17478 30708 17484
rect 29472 16590 29500 17478
rect 29748 17270 29776 17478
rect 29736 17264 29788 17270
rect 29736 17206 29788 17212
rect 30208 17202 30236 17478
rect 30668 17270 30696 17478
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30760 17202 30788 18022
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 30196 17196 30248 17202
rect 30196 17138 30248 17144
rect 30564 17196 30616 17202
rect 30564 17138 30616 17144
rect 30748 17196 30800 17202
rect 30748 17138 30800 17144
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 29368 16448 29420 16454
rect 29368 16390 29420 16396
rect 29380 16250 29408 16390
rect 29368 16244 29420 16250
rect 29368 16186 29420 16192
rect 29288 16102 29408 16130
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 28632 15972 28684 15978
rect 28632 15914 28684 15920
rect 27816 15830 27936 15858
rect 28540 15904 28592 15910
rect 28540 15846 28592 15852
rect 27712 15428 27764 15434
rect 27712 15370 27764 15376
rect 27620 15088 27672 15094
rect 27620 15030 27672 15036
rect 27632 14482 27660 15030
rect 27620 14476 27672 14482
rect 27620 14418 27672 14424
rect 27712 13728 27764 13734
rect 27712 13670 27764 13676
rect 27724 13326 27752 13670
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27356 12850 27476 12866
rect 27632 12850 27660 13126
rect 27344 12844 27476 12850
rect 27396 12838 27476 12844
rect 27620 12844 27672 12850
rect 27344 12786 27396 12792
rect 27620 12786 27672 12792
rect 27712 12708 27764 12714
rect 27712 12650 27764 12656
rect 27620 12640 27672 12646
rect 27540 12588 27620 12594
rect 27540 12582 27672 12588
rect 27540 12566 27660 12582
rect 27540 12434 27568 12566
rect 27172 12406 27292 12434
rect 27540 12406 27660 12434
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 27264 11694 27292 12406
rect 27632 11898 27660 12406
rect 27528 11892 27580 11898
rect 27528 11834 27580 11840
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27540 11778 27568 11834
rect 27724 11778 27752 12650
rect 27816 11830 27844 15830
rect 28552 15706 28580 15846
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28172 14952 28224 14958
rect 28172 14894 28224 14900
rect 27896 13932 27948 13938
rect 27896 13874 27948 13880
rect 27908 12288 27936 13874
rect 28078 12880 28134 12889
rect 28184 12850 28212 14894
rect 28368 14278 28396 15302
rect 28552 14890 28580 15642
rect 28644 15502 28672 15914
rect 28632 15496 28684 15502
rect 28632 15438 28684 15444
rect 28540 14884 28592 14890
rect 28540 14826 28592 14832
rect 28644 14618 28672 15438
rect 28736 14958 28764 15982
rect 28816 15904 28868 15910
rect 28816 15846 28868 15852
rect 28828 15026 28856 15846
rect 29288 15638 29316 15982
rect 29276 15632 29328 15638
rect 29276 15574 29328 15580
rect 29092 15156 29144 15162
rect 29092 15098 29144 15104
rect 29104 15026 29132 15098
rect 29380 15026 29408 16102
rect 29472 15570 29500 16526
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 29460 15156 29512 15162
rect 29460 15098 29512 15104
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 29092 15020 29144 15026
rect 29092 14962 29144 14968
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 28724 14952 28776 14958
rect 28724 14894 28776 14900
rect 28632 14612 28684 14618
rect 28632 14554 28684 14560
rect 29092 14340 29144 14346
rect 29092 14282 29144 14288
rect 28356 14272 28408 14278
rect 28356 14214 28408 14220
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28368 13870 28396 14214
rect 28356 13864 28408 13870
rect 28356 13806 28408 13812
rect 28448 13864 28500 13870
rect 28448 13806 28500 13812
rect 28264 13796 28316 13802
rect 28264 13738 28316 13744
rect 28276 13190 28304 13738
rect 28460 13462 28488 13806
rect 28448 13456 28500 13462
rect 28448 13398 28500 13404
rect 28540 13456 28592 13462
rect 28540 13398 28592 13404
rect 28552 13258 28580 13398
rect 28724 13320 28776 13326
rect 28724 13262 28776 13268
rect 28540 13252 28592 13258
rect 28540 13194 28592 13200
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 28736 12986 28764 13262
rect 28724 12980 28776 12986
rect 28724 12922 28776 12928
rect 28078 12815 28080 12824
rect 28132 12815 28134 12824
rect 28172 12844 28224 12850
rect 28080 12786 28132 12792
rect 28172 12786 28224 12792
rect 28724 12844 28776 12850
rect 28724 12786 28776 12792
rect 28000 12714 28212 12730
rect 27988 12708 28224 12714
rect 28040 12702 28172 12708
rect 27988 12650 28040 12656
rect 28172 12650 28224 12656
rect 28736 12646 28764 12786
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28724 12640 28776 12646
rect 28724 12582 28776 12588
rect 27988 12300 28040 12306
rect 27908 12260 27988 12288
rect 27540 11750 27752 11778
rect 27804 11824 27856 11830
rect 27804 11766 27856 11772
rect 27908 11762 27936 12260
rect 27988 12242 28040 12248
rect 28644 12102 28672 12582
rect 28632 12096 28684 12102
rect 28632 12038 28684 12044
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 27252 11688 27304 11694
rect 27252 11630 27304 11636
rect 28724 11552 28776 11558
rect 28724 11494 28776 11500
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27712 11008 27764 11014
rect 27342 10976 27398 10985
rect 27712 10950 27764 10956
rect 27342 10911 27398 10920
rect 26792 10736 26844 10742
rect 26792 10678 26844 10684
rect 26884 10736 26936 10742
rect 26884 10678 26936 10684
rect 27356 10674 27384 10911
rect 27724 10810 27752 10950
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 26700 10532 26752 10538
rect 26700 10474 26752 10480
rect 26608 9988 26660 9994
rect 26608 9930 26660 9936
rect 26620 9654 26648 9930
rect 26608 9648 26660 9654
rect 26608 9590 26660 9596
rect 26712 9586 26740 10474
rect 28000 10198 28028 11086
rect 28736 10810 28764 11494
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 28092 10266 28488 10282
rect 28092 10260 28500 10266
rect 28092 10254 28448 10260
rect 27988 10192 28040 10198
rect 27988 10134 28040 10140
rect 27344 9920 27396 9926
rect 27344 9862 27396 9868
rect 27356 9654 27384 9862
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 26436 7818 26464 8978
rect 26792 8900 26844 8906
rect 26792 8842 26844 8848
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26804 8634 26832 8842
rect 26792 8628 26844 8634
rect 26792 8570 26844 8576
rect 26896 8498 26924 8842
rect 27172 8838 27200 9522
rect 27160 8832 27212 8838
rect 27160 8774 27212 8780
rect 27172 8634 27200 8774
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 26884 8492 26936 8498
rect 26884 8434 26936 8440
rect 26976 8492 27028 8498
rect 26976 8434 27028 8440
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 26988 8090 27016 8434
rect 26792 8084 26844 8090
rect 26792 8026 26844 8032
rect 26976 8084 27028 8090
rect 26976 8026 27028 8032
rect 26804 7886 26832 8026
rect 27172 8022 27200 8434
rect 27160 8016 27212 8022
rect 27160 7958 27212 7964
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 26424 7812 26476 7818
rect 26424 7754 26476 7760
rect 26252 7410 26280 7754
rect 27172 7478 27200 7958
rect 27356 7546 27384 9590
rect 28000 9586 28028 10134
rect 28092 10062 28120 10254
rect 28448 10202 28500 10208
rect 28264 10192 28316 10198
rect 28316 10140 28580 10146
rect 28264 10134 28580 10140
rect 28276 10118 28580 10134
rect 28552 10062 28580 10118
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 28540 10056 28592 10062
rect 28540 9998 28592 10004
rect 28172 9988 28224 9994
rect 28172 9930 28224 9936
rect 28184 9722 28212 9930
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 28276 9450 28304 9998
rect 28828 9738 28856 14214
rect 29104 14006 29132 14282
rect 29276 14272 29328 14278
rect 29276 14214 29328 14220
rect 29288 14006 29316 14214
rect 29092 14000 29144 14006
rect 29092 13942 29144 13948
rect 29276 14000 29328 14006
rect 29276 13942 29328 13948
rect 29000 13456 29052 13462
rect 29000 13398 29052 13404
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28920 12918 28948 13126
rect 28908 12912 28960 12918
rect 28908 12854 28960 12860
rect 28908 12164 28960 12170
rect 28908 12106 28960 12112
rect 28920 11830 28948 12106
rect 29012 11898 29040 13398
rect 29472 12986 29500 15098
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 29460 12980 29512 12986
rect 29460 12922 29512 12928
rect 29104 12220 29132 12922
rect 29368 12912 29420 12918
rect 29368 12854 29420 12860
rect 29276 12844 29328 12850
rect 29276 12786 29328 12792
rect 29288 12238 29316 12786
rect 29184 12232 29236 12238
rect 29104 12192 29184 12220
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 28908 11824 28960 11830
rect 28908 11766 28960 11772
rect 29104 11064 29132 12192
rect 29184 12174 29236 12180
rect 29276 12232 29328 12238
rect 29276 12174 29328 12180
rect 29184 11620 29236 11626
rect 29184 11562 29236 11568
rect 29196 11354 29224 11562
rect 29184 11348 29236 11354
rect 29184 11290 29236 11296
rect 29288 11286 29316 12174
rect 29276 11280 29328 11286
rect 29276 11222 29328 11228
rect 28920 11036 29132 11064
rect 28920 10606 28948 11036
rect 28908 10600 28960 10606
rect 28908 10542 28960 10548
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29104 9994 29132 10542
rect 29092 9988 29144 9994
rect 29092 9930 29144 9936
rect 28736 9722 28856 9738
rect 28724 9716 28856 9722
rect 28776 9710 28856 9716
rect 28776 9664 28856 9674
rect 28724 9658 28856 9664
rect 28736 9654 28856 9658
rect 28736 9648 28868 9654
rect 28736 9646 28816 9648
rect 28816 9590 28868 9596
rect 28264 9444 28316 9450
rect 28264 9386 28316 9392
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27436 7812 27488 7818
rect 27436 7754 27488 7760
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27160 7472 27212 7478
rect 27160 7414 27212 7420
rect 27356 7410 27384 7482
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 25596 6724 25648 6730
rect 25596 6666 25648 6672
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 25608 6390 25636 6666
rect 26068 6458 26096 7278
rect 26252 6866 26280 7346
rect 27448 7274 27476 7754
rect 27632 7342 27660 9318
rect 28828 8634 28856 9590
rect 29104 9382 29132 9930
rect 29092 9376 29144 9382
rect 29092 9318 29144 9324
rect 28816 8628 28868 8634
rect 28816 8570 28868 8576
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 28172 7744 28224 7750
rect 28172 7686 28224 7692
rect 28184 7478 28212 7686
rect 29104 7478 29132 7890
rect 28172 7472 28224 7478
rect 28172 7414 28224 7420
rect 29092 7472 29144 7478
rect 29092 7414 29144 7420
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 27620 7336 27672 7342
rect 27620 7278 27672 7284
rect 27436 7268 27488 7274
rect 27436 7210 27488 7216
rect 26976 7200 27028 7206
rect 26976 7142 27028 7148
rect 26988 7002 27016 7142
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 26240 6860 26292 6866
rect 26240 6802 26292 6808
rect 27448 6458 27476 7210
rect 27816 7002 27844 7346
rect 28908 7336 28960 7342
rect 29276 7336 29328 7342
rect 28960 7284 29040 7290
rect 28908 7278 29040 7284
rect 29276 7278 29328 7284
rect 28448 7268 28500 7274
rect 28920 7262 29040 7278
rect 28448 7210 28500 7216
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27816 6458 27844 6666
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 27436 6452 27488 6458
rect 27436 6394 27488 6400
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 28460 6390 28488 7210
rect 29012 6866 29040 7262
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 28448 6384 28500 6390
rect 28448 6326 28500 6332
rect 28736 6254 28764 6802
rect 28724 6248 28776 6254
rect 28724 6190 28776 6196
rect 28448 6112 28500 6118
rect 28448 6054 28500 6060
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 22928 5568 22980 5574
rect 22928 5510 22980 5516
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 28460 5166 28488 6054
rect 28736 5778 28764 6190
rect 29104 6186 29132 7142
rect 29288 7002 29316 7278
rect 29276 6996 29328 7002
rect 29276 6938 29328 6944
rect 29380 6730 29408 12854
rect 29472 12306 29500 12922
rect 29656 12918 29684 17138
rect 30208 16658 30236 17138
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30576 17082 30604 17138
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 30300 16794 30328 16934
rect 30288 16788 30340 16794
rect 30288 16730 30340 16736
rect 30196 16652 30248 16658
rect 30196 16594 30248 16600
rect 30392 16454 30420 17070
rect 30576 17054 30696 17082
rect 30380 16448 30432 16454
rect 30380 16390 30432 16396
rect 30392 16114 30420 16390
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29748 15366 29776 15438
rect 29736 15360 29788 15366
rect 29736 15302 29788 15308
rect 29828 14884 29880 14890
rect 29828 14826 29880 14832
rect 30472 14884 30524 14890
rect 30524 14844 30604 14872
rect 30472 14826 30524 14832
rect 29840 14482 29868 14826
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 29920 14476 29972 14482
rect 29920 14418 29972 14424
rect 29932 13462 29960 14418
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 29920 13456 29972 13462
rect 29920 13398 29972 13404
rect 30104 13252 30156 13258
rect 30104 13194 30156 13200
rect 29644 12912 29696 12918
rect 29550 12880 29606 12889
rect 29644 12854 29696 12860
rect 29550 12815 29606 12824
rect 29564 12442 29592 12815
rect 29552 12436 29604 12442
rect 30116 12434 30144 13194
rect 30392 12918 30420 14282
rect 30576 14278 30604 14844
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 30472 13864 30524 13870
rect 30472 13806 30524 13812
rect 30484 12986 30512 13806
rect 30576 13394 30604 14214
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30668 13258 30696 17054
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 30116 12406 30236 12434
rect 29552 12378 29604 12384
rect 29460 12300 29512 12306
rect 29460 12242 29512 12248
rect 30208 12238 30236 12406
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30208 11558 30236 12174
rect 30392 12102 30420 12854
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30392 11812 30420 12038
rect 30564 11824 30616 11830
rect 30392 11784 30564 11812
rect 29828 11552 29880 11558
rect 29828 11494 29880 11500
rect 30196 11552 30248 11558
rect 30196 11494 30248 11500
rect 29840 11082 29868 11494
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 29828 11076 29880 11082
rect 29828 11018 29880 11024
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30116 10130 30144 10406
rect 30208 10130 30236 10542
rect 30104 10124 30156 10130
rect 30104 10066 30156 10072
rect 30196 10124 30248 10130
rect 30196 10066 30248 10072
rect 30392 10062 30420 11290
rect 30484 11082 30512 11784
rect 30564 11766 30616 11772
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30472 11076 30524 11082
rect 30472 11018 30524 11024
rect 30576 11014 30604 11630
rect 30564 11008 30616 11014
rect 30564 10950 30616 10956
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 30196 9920 30248 9926
rect 30196 9862 30248 9868
rect 29564 9654 29592 9862
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29840 8974 29868 9318
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 29656 7818 29684 8570
rect 29748 8566 29776 8774
rect 29736 8560 29788 8566
rect 29736 8502 29788 8508
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 29644 7812 29696 7818
rect 29644 7754 29696 7760
rect 29460 7744 29512 7750
rect 29460 7686 29512 7692
rect 29472 7410 29500 7686
rect 29656 7562 29684 7754
rect 29564 7534 29684 7562
rect 29460 7404 29512 7410
rect 29460 7346 29512 7352
rect 29460 6928 29512 6934
rect 29460 6870 29512 6876
rect 29368 6724 29420 6730
rect 29368 6666 29420 6672
rect 29472 6254 29500 6870
rect 29564 6458 29592 7534
rect 29748 7410 29776 8230
rect 29840 8090 29868 8910
rect 29920 8900 29972 8906
rect 29920 8842 29972 8848
rect 29828 8084 29880 8090
rect 29828 8026 29880 8032
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 29656 7002 29684 7346
rect 29644 6996 29696 7002
rect 29644 6938 29696 6944
rect 29932 6798 29960 8842
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 29552 6452 29604 6458
rect 29552 6394 29604 6400
rect 29460 6248 29512 6254
rect 29460 6190 29512 6196
rect 29092 6180 29144 6186
rect 29092 6122 29144 6128
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 28736 5302 28764 5714
rect 29564 5642 29592 6394
rect 30024 6254 30052 8978
rect 30104 8900 30156 8906
rect 30104 8842 30156 8848
rect 30116 8294 30144 8842
rect 30104 8288 30156 8294
rect 30104 8230 30156 8236
rect 30208 6662 30236 9862
rect 30392 9586 30420 9998
rect 30472 9988 30524 9994
rect 30472 9930 30524 9936
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30484 9382 30512 9930
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30288 8900 30340 8906
rect 30288 8842 30340 8848
rect 30300 6934 30328 8842
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30288 6928 30340 6934
rect 30288 6870 30340 6876
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 30208 6390 30236 6598
rect 30196 6384 30248 6390
rect 30300 6361 30328 6870
rect 30484 6866 30512 7482
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30196 6326 30248 6332
rect 30286 6352 30342 6361
rect 30286 6287 30342 6296
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 30012 6248 30064 6254
rect 30576 6202 30604 10950
rect 30760 9364 30788 17138
rect 30944 16250 30972 18566
rect 31036 18222 31064 18770
rect 31024 18216 31076 18222
rect 31024 18158 31076 18164
rect 31128 18034 31156 19468
rect 31036 18006 31156 18034
rect 30932 16244 30984 16250
rect 30932 16186 30984 16192
rect 31036 16130 31064 18006
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 31128 17338 31156 17546
rect 31116 17332 31168 17338
rect 31116 17274 31168 17280
rect 30944 16102 31064 16130
rect 30840 12096 30892 12102
rect 30840 12038 30892 12044
rect 30852 10742 30880 12038
rect 30944 11898 30972 16102
rect 31312 15570 31340 23038
rect 31404 22030 31432 24142
rect 31496 24070 31524 24550
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 31484 23520 31536 23526
rect 31484 23462 31536 23468
rect 31496 23118 31524 23462
rect 31484 23112 31536 23118
rect 31484 23054 31536 23060
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 31484 21956 31536 21962
rect 31484 21898 31536 21904
rect 31496 21622 31524 21898
rect 31484 21616 31536 21622
rect 31484 21558 31536 21564
rect 31496 20806 31524 21558
rect 31484 20800 31536 20806
rect 31484 20742 31536 20748
rect 31588 19514 31616 25094
rect 31852 24948 31904 24954
rect 31852 24890 31904 24896
rect 31668 24404 31720 24410
rect 31668 24346 31720 24352
rect 31680 24138 31708 24346
rect 31864 24206 31892 24890
rect 31852 24200 31904 24206
rect 31852 24142 31904 24148
rect 31668 24132 31720 24138
rect 31668 24074 31720 24080
rect 31668 23860 31720 23866
rect 31668 23802 31720 23808
rect 31680 23594 31708 23802
rect 31760 23724 31812 23730
rect 31760 23666 31812 23672
rect 31668 23588 31720 23594
rect 31668 23530 31720 23536
rect 31772 23050 31800 23666
rect 32232 23186 32260 28999
rect 32312 28416 32364 28422
rect 32312 28358 32364 28364
rect 32324 28082 32352 28358
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32416 27554 32444 29446
rect 32600 27878 32628 29786
rect 32588 27872 32640 27878
rect 32588 27814 32640 27820
rect 32324 27526 32444 27554
rect 32324 23730 32352 27526
rect 32692 26450 32720 31282
rect 32772 29708 32824 29714
rect 32772 29650 32824 29656
rect 32784 28801 32812 29650
rect 32876 29510 32904 36654
rect 33416 36100 33468 36106
rect 33416 36042 33468 36048
rect 33324 35624 33376 35630
rect 33324 35566 33376 35572
rect 33232 35556 33284 35562
rect 33232 35498 33284 35504
rect 33048 34196 33100 34202
rect 33048 34138 33100 34144
rect 33060 33522 33088 34138
rect 33048 33516 33100 33522
rect 33048 33458 33100 33464
rect 33060 31278 33088 33458
rect 33244 33386 33272 35498
rect 33336 33658 33364 35566
rect 33428 35154 33456 36042
rect 33416 35148 33468 35154
rect 33416 35090 33468 35096
rect 33520 35086 33548 36722
rect 33508 35080 33560 35086
rect 33508 35022 33560 35028
rect 33520 34474 33548 35022
rect 33508 34468 33560 34474
rect 33508 34410 33560 34416
rect 33416 33992 33468 33998
rect 33520 33946 33548 34410
rect 33468 33940 33548 33946
rect 33416 33934 33548 33940
rect 33428 33918 33548 33934
rect 33324 33652 33376 33658
rect 33324 33594 33376 33600
rect 33232 33380 33284 33386
rect 33232 33322 33284 33328
rect 33612 32978 33640 37606
rect 33980 37330 34008 37810
rect 34152 37800 34204 37806
rect 34152 37742 34204 37748
rect 34164 37330 34192 37742
rect 33692 37324 33744 37330
rect 33692 37266 33744 37272
rect 33968 37324 34020 37330
rect 33968 37266 34020 37272
rect 34152 37324 34204 37330
rect 34152 37266 34204 37272
rect 33704 36922 33732 37266
rect 33966 37224 34022 37233
rect 33966 37159 33968 37168
rect 34020 37159 34022 37168
rect 33968 37130 34020 37136
rect 33692 36916 33744 36922
rect 33692 36858 33744 36864
rect 33784 36576 33836 36582
rect 33784 36518 33836 36524
rect 33968 36576 34020 36582
rect 33968 36518 34020 36524
rect 33796 36242 33824 36518
rect 33980 36310 34008 36518
rect 34164 36378 34192 37266
rect 34152 36372 34204 36378
rect 34152 36314 34204 36320
rect 33968 36304 34020 36310
rect 33968 36246 34020 36252
rect 33784 36236 33836 36242
rect 33784 36178 33836 36184
rect 33796 36106 33824 36178
rect 33784 36100 33836 36106
rect 33784 36042 33836 36048
rect 34164 35562 34192 36314
rect 34612 36100 34664 36106
rect 34612 36042 34664 36048
rect 34520 36032 34572 36038
rect 34520 35974 34572 35980
rect 34532 35766 34560 35974
rect 34520 35760 34572 35766
rect 34520 35702 34572 35708
rect 34520 35624 34572 35630
rect 34624 35578 34652 36042
rect 34572 35572 34652 35578
rect 34520 35566 34652 35572
rect 34152 35556 34204 35562
rect 34152 35498 34204 35504
rect 34532 35550 34652 35566
rect 34428 35488 34480 35494
rect 34428 35430 34480 35436
rect 33784 35080 33836 35086
rect 33784 35022 33836 35028
rect 33796 34202 33824 35022
rect 34440 35018 34468 35430
rect 34532 35290 34560 35550
rect 34520 35284 34572 35290
rect 34520 35226 34572 35232
rect 34428 35012 34480 35018
rect 34428 34954 34480 34960
rect 34336 34944 34388 34950
rect 34336 34886 34388 34892
rect 34348 34678 34376 34886
rect 34440 34678 34468 34954
rect 34336 34672 34388 34678
rect 34336 34614 34388 34620
rect 34428 34672 34480 34678
rect 34428 34614 34480 34620
rect 34428 34536 34480 34542
rect 34428 34478 34480 34484
rect 33968 34400 34020 34406
rect 33968 34342 34020 34348
rect 33784 34196 33836 34202
rect 33784 34138 33836 34144
rect 33980 34066 34008 34342
rect 33968 34060 34020 34066
rect 33968 34002 34020 34008
rect 34440 33658 34468 34478
rect 34244 33652 34296 33658
rect 34244 33594 34296 33600
rect 34428 33652 34480 33658
rect 34428 33594 34480 33600
rect 34256 33538 34284 33594
rect 34152 33516 34204 33522
rect 34256 33510 34468 33538
rect 34152 33458 34204 33464
rect 33600 32972 33652 32978
rect 33600 32914 33652 32920
rect 33968 32972 34020 32978
rect 33968 32914 34020 32920
rect 33692 32768 33744 32774
rect 33692 32710 33744 32716
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 33336 31482 33364 32370
rect 33704 31822 33732 32710
rect 33980 32026 34008 32914
rect 34164 32570 34192 33458
rect 34440 33454 34468 33510
rect 34428 33448 34480 33454
rect 34428 33390 34480 33396
rect 34244 33312 34296 33318
rect 34244 33254 34296 33260
rect 34256 32978 34284 33254
rect 34244 32972 34296 32978
rect 34244 32914 34296 32920
rect 34336 32836 34388 32842
rect 34336 32778 34388 32784
rect 34152 32564 34204 32570
rect 34152 32506 34204 32512
rect 33968 32020 34020 32026
rect 33968 31962 34020 31968
rect 33692 31816 33744 31822
rect 33692 31758 33744 31764
rect 33508 31680 33560 31686
rect 33508 31622 33560 31628
rect 33324 31476 33376 31482
rect 33324 31418 33376 31424
rect 33140 31408 33192 31414
rect 33140 31350 33192 31356
rect 33048 31272 33100 31278
rect 33048 31214 33100 31220
rect 33152 30598 33180 31350
rect 33416 30728 33468 30734
rect 33520 30682 33548 31622
rect 33784 31476 33836 31482
rect 33784 31418 33836 31424
rect 33468 30676 33548 30682
rect 33416 30670 33548 30676
rect 33428 30654 33548 30670
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 33152 30258 33180 30534
rect 32956 30252 33008 30258
rect 32956 30194 33008 30200
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 32968 29850 32996 30194
rect 33152 29850 33180 30194
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 33140 29844 33192 29850
rect 33140 29786 33192 29792
rect 33048 29572 33100 29578
rect 33048 29514 33100 29520
rect 32864 29504 32916 29510
rect 32864 29446 32916 29452
rect 32876 29306 32904 29446
rect 33060 29306 33088 29514
rect 32864 29300 32916 29306
rect 32864 29242 32916 29248
rect 33048 29300 33100 29306
rect 33048 29242 33100 29248
rect 32954 29200 33010 29209
rect 33152 29170 33180 29786
rect 33416 29640 33468 29646
rect 33336 29600 33416 29628
rect 33232 29300 33284 29306
rect 33232 29242 33284 29248
rect 32954 29135 33010 29144
rect 33048 29164 33100 29170
rect 32770 28792 32826 28801
rect 32770 28727 32826 28736
rect 32784 28150 32812 28727
rect 32772 28144 32824 28150
rect 32772 28086 32824 28092
rect 32772 26920 32824 26926
rect 32772 26862 32824 26868
rect 32680 26444 32732 26450
rect 32680 26386 32732 26392
rect 32692 26042 32720 26386
rect 32784 26314 32812 26862
rect 32968 26586 32996 29135
rect 33048 29106 33100 29112
rect 33140 29164 33192 29170
rect 33140 29106 33192 29112
rect 33060 28994 33088 29106
rect 33060 28966 33180 28994
rect 33152 28218 33180 28966
rect 33140 28212 33192 28218
rect 33140 28154 33192 28160
rect 33152 28121 33180 28154
rect 33138 28112 33194 28121
rect 33138 28047 33194 28056
rect 33244 27470 33272 29242
rect 33336 29073 33364 29600
rect 33416 29582 33468 29588
rect 33416 29504 33468 29510
rect 33416 29446 33468 29452
rect 33428 29102 33456 29446
rect 33416 29096 33468 29102
rect 33322 29064 33378 29073
rect 33416 29038 33468 29044
rect 33322 28999 33378 29008
rect 33520 28234 33548 30654
rect 33692 30184 33744 30190
rect 33692 30126 33744 30132
rect 33704 29850 33732 30126
rect 33692 29844 33744 29850
rect 33692 29786 33744 29792
rect 33598 29744 33654 29753
rect 33598 29679 33654 29688
rect 33612 29646 33640 29679
rect 33600 29640 33652 29646
rect 33600 29582 33652 29588
rect 33598 29472 33654 29481
rect 33598 29407 33654 29416
rect 33612 29034 33640 29407
rect 33796 29152 33824 31418
rect 33980 31278 34008 31962
rect 34164 31754 34192 32506
rect 34348 31754 34376 32778
rect 34440 32230 34468 33390
rect 34716 32910 34744 39494
rect 34796 39432 34848 39438
rect 34796 39374 34848 39380
rect 34808 38554 34836 39374
rect 34900 39030 34928 39578
rect 35164 39364 35216 39370
rect 35164 39306 35216 39312
rect 34888 39024 34940 39030
rect 34888 38966 34940 38972
rect 34900 38758 34928 38966
rect 35176 38865 35204 39306
rect 35268 38894 35296 39578
rect 35360 39506 35388 39782
rect 35348 39500 35400 39506
rect 35348 39442 35400 39448
rect 35452 39386 35480 41074
rect 36004 40594 36032 42026
rect 37476 41614 37504 42094
rect 37740 42016 37792 42022
rect 37740 41958 37792 41964
rect 37464 41608 37516 41614
rect 37516 41556 37596 41562
rect 37464 41550 37596 41556
rect 37476 41534 37596 41550
rect 37464 41472 37516 41478
rect 37464 41414 37516 41420
rect 37372 41200 37424 41206
rect 37372 41142 37424 41148
rect 36820 40928 36872 40934
rect 36820 40870 36872 40876
rect 37188 40928 37240 40934
rect 37188 40870 37240 40876
rect 37280 40928 37332 40934
rect 37280 40870 37332 40876
rect 35992 40588 36044 40594
rect 35992 40530 36044 40536
rect 35594 40284 35902 40293
rect 35594 40282 35600 40284
rect 35656 40282 35680 40284
rect 35736 40282 35760 40284
rect 35816 40282 35840 40284
rect 35896 40282 35902 40284
rect 35656 40230 35658 40282
rect 35838 40230 35840 40282
rect 35594 40228 35600 40230
rect 35656 40228 35680 40230
rect 35736 40228 35760 40230
rect 35816 40228 35840 40230
rect 35896 40228 35902 40230
rect 35594 40219 35902 40228
rect 36832 40118 36860 40870
rect 37200 40610 37228 40870
rect 37292 40730 37320 40870
rect 37384 40730 37412 41142
rect 37280 40724 37332 40730
rect 37280 40666 37332 40672
rect 37372 40724 37424 40730
rect 37372 40666 37424 40672
rect 37200 40582 37412 40610
rect 36820 40112 36872 40118
rect 36820 40054 36872 40060
rect 36832 39438 36860 40054
rect 37384 39438 37412 40582
rect 37476 40050 37504 41414
rect 37568 41206 37596 41534
rect 37648 41540 37700 41546
rect 37648 41482 37700 41488
rect 37556 41200 37608 41206
rect 37556 41142 37608 41148
rect 37660 40934 37688 41482
rect 37752 41274 37780 41958
rect 38016 41676 38068 41682
rect 38016 41618 38068 41624
rect 37832 41540 37884 41546
rect 37832 41482 37884 41488
rect 37740 41268 37792 41274
rect 37740 41210 37792 41216
rect 37844 41206 37872 41482
rect 37924 41472 37976 41478
rect 37924 41414 37976 41420
rect 37936 41206 37964 41414
rect 37832 41200 37884 41206
rect 37832 41142 37884 41148
rect 37924 41200 37976 41206
rect 37924 41142 37976 41148
rect 37832 41064 37884 41070
rect 38028 41018 38056 41618
rect 38108 41540 38160 41546
rect 38108 41482 38160 41488
rect 37884 41012 38056 41018
rect 37832 41006 38056 41012
rect 37844 40990 38056 41006
rect 37648 40928 37700 40934
rect 37648 40870 37700 40876
rect 38028 40662 38056 40990
rect 38016 40656 38068 40662
rect 38016 40598 38068 40604
rect 38120 40458 38148 41482
rect 38580 41206 38608 42094
rect 39488 42016 39540 42022
rect 39488 41958 39540 41964
rect 39028 41676 39080 41682
rect 39028 41618 39080 41624
rect 39040 41414 39068 41618
rect 39396 41540 39448 41546
rect 39396 41482 39448 41488
rect 39040 41386 39252 41414
rect 38568 41200 38620 41206
rect 38568 41142 38620 41148
rect 38292 41132 38344 41138
rect 38292 41074 38344 41080
rect 38304 40730 38332 41074
rect 38844 41064 38896 41070
rect 38844 41006 38896 41012
rect 38292 40724 38344 40730
rect 38292 40666 38344 40672
rect 38108 40452 38160 40458
rect 38108 40394 38160 40400
rect 38856 40118 38884 41006
rect 39224 40526 39252 41386
rect 39408 41274 39436 41482
rect 39500 41274 39528 41958
rect 39396 41268 39448 41274
rect 39396 41210 39448 41216
rect 39488 41268 39540 41274
rect 39488 41210 39540 41216
rect 39580 41132 39632 41138
rect 39580 41074 39632 41080
rect 40224 41132 40276 41138
rect 40224 41074 40276 41080
rect 39304 41064 39356 41070
rect 39304 41006 39356 41012
rect 39212 40520 39264 40526
rect 39212 40462 39264 40468
rect 38292 40112 38344 40118
rect 38292 40054 38344 40060
rect 38844 40112 38896 40118
rect 38844 40054 38896 40060
rect 37464 40044 37516 40050
rect 37464 39986 37516 39992
rect 35360 39358 35480 39386
rect 36820 39432 36872 39438
rect 36820 39374 36872 39380
rect 37372 39432 37424 39438
rect 37372 39374 37424 39380
rect 36636 39364 36688 39370
rect 35256 38888 35308 38894
rect 35162 38856 35218 38865
rect 35256 38830 35308 38836
rect 35162 38791 35218 38800
rect 34888 38752 34940 38758
rect 34888 38694 34940 38700
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34796 38548 34848 38554
rect 34796 38490 34848 38496
rect 35072 38480 35124 38486
rect 35072 38422 35124 38428
rect 35084 38350 35112 38422
rect 35360 38400 35388 39358
rect 36636 39306 36688 39312
rect 35440 39296 35492 39302
rect 35440 39238 35492 39244
rect 35268 38372 35388 38400
rect 34796 38344 34848 38350
rect 34796 38286 34848 38292
rect 34888 38344 34940 38350
rect 34888 38286 34940 38292
rect 35072 38344 35124 38350
rect 35072 38286 35124 38292
rect 34808 37942 34836 38286
rect 34900 38214 34928 38286
rect 34888 38208 34940 38214
rect 34888 38150 34940 38156
rect 34796 37936 34848 37942
rect 34796 37878 34848 37884
rect 34900 37788 34928 38150
rect 34808 37760 34928 37788
rect 34808 37330 34836 37760
rect 35084 37738 35112 38286
rect 35072 37732 35124 37738
rect 35072 37674 35124 37680
rect 35268 37670 35296 38372
rect 35452 38298 35480 39238
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 36176 39092 36228 39098
rect 36176 39034 36228 39040
rect 35714 38856 35770 38865
rect 35714 38791 35716 38800
rect 35768 38791 35770 38800
rect 35716 38762 35768 38768
rect 35624 38752 35676 38758
rect 35624 38694 35676 38700
rect 35992 38752 36044 38758
rect 35992 38694 36044 38700
rect 35636 38536 35664 38694
rect 35636 38508 35756 38536
rect 35360 38270 35480 38298
rect 35728 38282 35756 38508
rect 35716 38276 35768 38282
rect 35256 37664 35308 37670
rect 35256 37606 35308 37612
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37324 34848 37330
rect 34796 37266 34848 37272
rect 34980 37256 35032 37262
rect 34980 37198 35032 37204
rect 35256 37256 35308 37262
rect 35256 37198 35308 37204
rect 34992 36922 35020 37198
rect 34980 36916 35032 36922
rect 34980 36858 35032 36864
rect 35268 36854 35296 37198
rect 35360 37194 35388 38270
rect 35716 38218 35768 38224
rect 35440 38208 35492 38214
rect 35440 38150 35492 38156
rect 35452 38010 35480 38150
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 35440 38004 35492 38010
rect 35440 37946 35492 37952
rect 36004 37874 36032 38694
rect 35992 37868 36044 37874
rect 35992 37810 36044 37816
rect 35348 37188 35400 37194
rect 35348 37130 35400 37136
rect 35256 36848 35308 36854
rect 35256 36790 35308 36796
rect 35360 36786 35388 37130
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 35348 36780 35400 36786
rect 35348 36722 35400 36728
rect 34796 36712 34848 36718
rect 34796 36654 34848 36660
rect 34808 36378 34836 36654
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34796 36372 34848 36378
rect 34796 36314 34848 36320
rect 34888 36304 34940 36310
rect 35360 36258 35388 36722
rect 35716 36644 35768 36650
rect 35716 36586 35768 36592
rect 35992 36644 36044 36650
rect 35992 36586 36044 36592
rect 34888 36246 34940 36252
rect 34796 36100 34848 36106
rect 34796 36042 34848 36048
rect 34808 35766 34836 36042
rect 34900 35834 34928 36246
rect 35268 36230 35388 36258
rect 35268 36174 35296 36230
rect 35256 36168 35308 36174
rect 35256 36110 35308 36116
rect 35728 36020 35756 36586
rect 35452 35992 35756 36020
rect 35452 35834 35480 35992
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 34888 35828 34940 35834
rect 34888 35770 34940 35776
rect 35440 35828 35492 35834
rect 35440 35770 35492 35776
rect 34796 35760 34848 35766
rect 34796 35702 34848 35708
rect 35164 35692 35216 35698
rect 35164 35634 35216 35640
rect 35176 35578 35204 35634
rect 35808 35624 35860 35630
rect 35176 35562 35480 35578
rect 35808 35566 35860 35572
rect 35176 35556 35492 35562
rect 35176 35550 35440 35556
rect 35440 35498 35492 35504
rect 34796 35488 34848 35494
rect 34796 35430 34848 35436
rect 35348 35488 35400 35494
rect 35348 35430 35400 35436
rect 34808 34678 34836 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35360 35290 35388 35430
rect 35348 35284 35400 35290
rect 35348 35226 35400 35232
rect 35820 35222 35848 35566
rect 35808 35216 35860 35222
rect 35808 35158 35860 35164
rect 36004 35154 36032 36586
rect 36188 36242 36216 39034
rect 36648 38962 36676 39306
rect 36636 38956 36688 38962
rect 36636 38898 36688 38904
rect 37384 38826 37412 39374
rect 38200 39364 38252 39370
rect 38200 39306 38252 39312
rect 37648 39296 37700 39302
rect 37648 39238 37700 39244
rect 37660 38962 37688 39238
rect 38212 38962 38240 39306
rect 37648 38956 37700 38962
rect 37648 38898 37700 38904
rect 38108 38956 38160 38962
rect 38108 38898 38160 38904
rect 38200 38956 38252 38962
rect 38200 38898 38252 38904
rect 37372 38820 37424 38826
rect 37372 38762 37424 38768
rect 38016 38820 38068 38826
rect 38016 38762 38068 38768
rect 37832 38752 37884 38758
rect 37832 38694 37884 38700
rect 37740 38344 37792 38350
rect 37740 38286 37792 38292
rect 37188 38208 37240 38214
rect 37188 38150 37240 38156
rect 37200 38010 37228 38150
rect 37188 38004 37240 38010
rect 37188 37946 37240 37952
rect 37464 37256 37516 37262
rect 37648 37256 37700 37262
rect 37516 37216 37596 37244
rect 37464 37198 37516 37204
rect 36360 37120 36412 37126
rect 36360 37062 36412 37068
rect 37280 37120 37332 37126
rect 37280 37062 37332 37068
rect 36372 36786 36400 37062
rect 36360 36780 36412 36786
rect 36360 36722 36412 36728
rect 36452 36712 36504 36718
rect 36452 36654 36504 36660
rect 36464 36378 36492 36654
rect 37188 36576 37240 36582
rect 37188 36518 37240 36524
rect 37200 36378 37228 36518
rect 36452 36372 36504 36378
rect 36452 36314 36504 36320
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 36176 36236 36228 36242
rect 36176 36178 36228 36184
rect 37292 36174 37320 37062
rect 37464 36916 37516 36922
rect 37464 36858 37516 36864
rect 37476 36825 37504 36858
rect 37462 36816 37518 36825
rect 37372 36780 37424 36786
rect 37462 36751 37518 36760
rect 37372 36722 37424 36728
rect 37384 36174 37412 36722
rect 37568 36650 37596 37216
rect 37648 37198 37700 37204
rect 37660 36786 37688 37198
rect 37752 36802 37780 38286
rect 37844 37874 37872 38694
rect 38028 38418 38056 38762
rect 38016 38412 38068 38418
rect 38016 38354 38068 38360
rect 38120 38350 38148 38898
rect 38212 38486 38240 38898
rect 38200 38480 38252 38486
rect 38200 38422 38252 38428
rect 38108 38344 38160 38350
rect 38108 38286 38160 38292
rect 37924 38208 37976 38214
rect 37924 38150 37976 38156
rect 37832 37868 37884 37874
rect 37832 37810 37884 37816
rect 37936 37262 37964 38150
rect 37924 37256 37976 37262
rect 37924 37198 37976 37204
rect 37648 36780 37700 36786
rect 37752 36774 37872 36802
rect 37648 36722 37700 36728
rect 37556 36644 37608 36650
rect 37556 36586 37608 36592
rect 37464 36576 37516 36582
rect 37464 36518 37516 36524
rect 37476 36310 37504 36518
rect 37464 36304 37516 36310
rect 37464 36246 37516 36252
rect 37568 36174 37596 36586
rect 37660 36310 37688 36722
rect 37648 36304 37700 36310
rect 37648 36246 37700 36252
rect 37280 36168 37332 36174
rect 37280 36110 37332 36116
rect 37372 36168 37424 36174
rect 37372 36110 37424 36116
rect 37556 36168 37608 36174
rect 37556 36110 37608 36116
rect 36084 36032 36136 36038
rect 36084 35974 36136 35980
rect 36096 35698 36124 35974
rect 36084 35692 36136 35698
rect 36084 35634 36136 35640
rect 37648 35488 37700 35494
rect 37648 35430 37700 35436
rect 37096 35216 37148 35222
rect 37096 35158 37148 35164
rect 35992 35148 36044 35154
rect 35992 35090 36044 35096
rect 37004 35080 37056 35086
rect 37004 35022 37056 35028
rect 35348 34944 35400 34950
rect 35348 34886 35400 34892
rect 36268 34944 36320 34950
rect 36268 34886 36320 34892
rect 34796 34672 34848 34678
rect 34796 34614 34848 34620
rect 34796 34536 34848 34542
rect 34796 34478 34848 34484
rect 34808 34066 34836 34478
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34796 34060 34848 34066
rect 34796 34002 34848 34008
rect 34704 32904 34756 32910
rect 34704 32846 34756 32852
rect 34612 32836 34664 32842
rect 34612 32778 34664 32784
rect 34428 32224 34480 32230
rect 34428 32166 34480 32172
rect 34440 32026 34468 32166
rect 34428 32020 34480 32026
rect 34428 31962 34480 31968
rect 34164 31726 34284 31754
rect 34348 31726 34468 31754
rect 34256 31346 34284 31726
rect 34244 31340 34296 31346
rect 34244 31282 34296 31288
rect 33968 31272 34020 31278
rect 33968 31214 34020 31220
rect 34336 30252 34388 30258
rect 34336 30194 34388 30200
rect 34242 30152 34298 30161
rect 33968 30116 34020 30122
rect 34242 30087 34298 30096
rect 33968 30058 34020 30064
rect 33874 29608 33930 29617
rect 33874 29543 33876 29552
rect 33928 29543 33930 29552
rect 33876 29514 33928 29520
rect 33876 29164 33928 29170
rect 33796 29124 33876 29152
rect 33876 29106 33928 29112
rect 33600 29028 33652 29034
rect 33600 28970 33652 28976
rect 33520 28206 33732 28234
rect 33888 28218 33916 29106
rect 33600 28076 33652 28082
rect 33600 28018 33652 28024
rect 33508 28008 33560 28014
rect 33508 27950 33560 27956
rect 33520 27606 33548 27950
rect 33612 27674 33640 28018
rect 33600 27668 33652 27674
rect 33600 27610 33652 27616
rect 33508 27600 33560 27606
rect 33508 27542 33560 27548
rect 33048 27464 33100 27470
rect 33048 27406 33100 27412
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33060 26772 33088 27406
rect 33060 26744 33180 26772
rect 33152 26586 33180 26744
rect 32956 26580 33008 26586
rect 32956 26522 33008 26528
rect 33140 26580 33192 26586
rect 33140 26522 33192 26528
rect 32772 26308 32824 26314
rect 32772 26250 32824 26256
rect 32784 26042 32812 26250
rect 33244 26246 33272 27406
rect 33600 26920 33652 26926
rect 33600 26862 33652 26868
rect 33612 26382 33640 26862
rect 33704 26586 33732 28206
rect 33876 28212 33928 28218
rect 33876 28154 33928 28160
rect 33888 28082 33916 28154
rect 33876 28076 33928 28082
rect 33876 28018 33928 28024
rect 33784 27872 33836 27878
rect 33784 27814 33836 27820
rect 33796 27674 33824 27814
rect 33980 27713 34008 30058
rect 34152 29844 34204 29850
rect 34152 29786 34204 29792
rect 34060 29572 34112 29578
rect 34060 29514 34112 29520
rect 34072 29238 34100 29514
rect 34060 29232 34112 29238
rect 34060 29174 34112 29180
rect 34072 28626 34100 29174
rect 34164 29034 34192 29786
rect 34256 29782 34284 30087
rect 34244 29776 34296 29782
rect 34244 29718 34296 29724
rect 34256 29034 34284 29718
rect 34348 29238 34376 30194
rect 34440 30138 34468 31726
rect 34624 30433 34652 32778
rect 34808 32570 34836 34002
rect 35360 33930 35388 34886
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 35532 34672 35584 34678
rect 35532 34614 35584 34620
rect 35544 34542 35572 34614
rect 35532 34536 35584 34542
rect 35532 34478 35584 34484
rect 35624 34536 35676 34542
rect 35624 34478 35676 34484
rect 35544 34406 35572 34478
rect 35532 34400 35584 34406
rect 35532 34342 35584 34348
rect 35544 33930 35572 34342
rect 35636 34066 35664 34478
rect 35624 34060 35676 34066
rect 35624 34002 35676 34008
rect 35348 33924 35400 33930
rect 35348 33866 35400 33872
rect 35532 33924 35584 33930
rect 35532 33866 35584 33872
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 36280 33658 36308 34886
rect 37016 34474 37044 35022
rect 37108 34678 37136 35158
rect 37556 34944 37608 34950
rect 37556 34886 37608 34892
rect 37096 34672 37148 34678
rect 37096 34614 37148 34620
rect 37280 34536 37332 34542
rect 37280 34478 37332 34484
rect 37004 34468 37056 34474
rect 37004 34410 37056 34416
rect 36728 33856 36780 33862
rect 36728 33798 36780 33804
rect 36820 33856 36872 33862
rect 36820 33798 36872 33804
rect 36268 33652 36320 33658
rect 36268 33594 36320 33600
rect 36740 33454 36768 33798
rect 36832 33590 36860 33798
rect 36820 33584 36872 33590
rect 36820 33526 36872 33532
rect 36728 33448 36780 33454
rect 36728 33390 36780 33396
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35440 32904 35492 32910
rect 35440 32846 35492 32852
rect 34888 32768 34940 32774
rect 34888 32710 34940 32716
rect 34980 32768 35032 32774
rect 34980 32710 35032 32716
rect 34900 32570 34928 32710
rect 34796 32564 34848 32570
rect 34796 32506 34848 32512
rect 34888 32564 34940 32570
rect 34888 32506 34940 32512
rect 34808 31890 34836 32506
rect 34992 32502 35020 32710
rect 34980 32496 35032 32502
rect 34980 32438 35032 32444
rect 35452 32314 35480 32846
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 35452 32286 35572 32314
rect 35544 32230 35572 32286
rect 35532 32224 35584 32230
rect 35532 32166 35584 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34796 31884 34848 31890
rect 34796 31826 34848 31832
rect 35348 31748 35400 31754
rect 35348 31690 35400 31696
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30938 35388 31690
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 35348 30932 35400 30938
rect 35348 30874 35400 30880
rect 35716 30796 35768 30802
rect 35716 30738 35768 30744
rect 35072 30728 35124 30734
rect 35532 30728 35584 30734
rect 35072 30670 35124 30676
rect 35452 30676 35532 30682
rect 35728 30705 35756 30738
rect 35452 30670 35584 30676
rect 35714 30696 35770 30705
rect 34610 30424 34666 30433
rect 35084 30394 35112 30670
rect 35348 30660 35400 30666
rect 35348 30602 35400 30608
rect 35452 30654 35572 30670
rect 34610 30359 34666 30368
rect 35072 30388 35124 30394
rect 35072 30330 35124 30336
rect 34704 30320 34756 30326
rect 34704 30262 34756 30268
rect 34612 30184 34664 30190
rect 34440 30110 34560 30138
rect 34612 30126 34664 30132
rect 34428 30048 34480 30054
rect 34428 29990 34480 29996
rect 34440 29714 34468 29990
rect 34428 29708 34480 29714
rect 34428 29650 34480 29656
rect 34336 29232 34388 29238
rect 34336 29174 34388 29180
rect 34152 29028 34204 29034
rect 34152 28970 34204 28976
rect 34244 29028 34296 29034
rect 34244 28970 34296 28976
rect 34242 28928 34298 28937
rect 34242 28863 34298 28872
rect 34060 28620 34112 28626
rect 34060 28562 34112 28568
rect 34152 28484 34204 28490
rect 34152 28426 34204 28432
rect 33966 27704 34022 27713
rect 33784 27668 33836 27674
rect 33966 27639 34022 27648
rect 33784 27610 33836 27616
rect 33980 27606 34008 27639
rect 34164 27606 34192 28426
rect 33876 27600 33928 27606
rect 33782 27568 33838 27577
rect 33876 27542 33928 27548
rect 33968 27600 34020 27606
rect 34152 27600 34204 27606
rect 33968 27542 34020 27548
rect 34058 27568 34114 27577
rect 33782 27503 33838 27512
rect 33796 27470 33824 27503
rect 33784 27464 33836 27470
rect 33784 27406 33836 27412
rect 33888 27418 33916 27542
rect 34152 27542 34204 27548
rect 34058 27503 34114 27512
rect 34072 27418 34100 27503
rect 33692 26580 33744 26586
rect 33692 26522 33744 26528
rect 33796 26450 33824 27406
rect 33888 27390 34100 27418
rect 33876 27328 33928 27334
rect 34060 27328 34112 27334
rect 33928 27288 34008 27316
rect 33876 27270 33928 27276
rect 33876 27056 33928 27062
rect 33876 26998 33928 27004
rect 33888 26586 33916 26998
rect 33876 26580 33928 26586
rect 33876 26522 33928 26528
rect 33784 26444 33836 26450
rect 33784 26386 33836 26392
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 33232 26240 33284 26246
rect 33232 26182 33284 26188
rect 32680 26036 32732 26042
rect 32680 25978 32732 25984
rect 32772 26036 32824 26042
rect 32772 25978 32824 25984
rect 32588 25288 32640 25294
rect 32588 25230 32640 25236
rect 32496 25220 32548 25226
rect 32496 25162 32548 25168
rect 32508 24070 32536 25162
rect 32600 24886 32628 25230
rect 32692 24954 32720 25978
rect 32864 25696 32916 25702
rect 32864 25638 32916 25644
rect 32680 24948 32732 24954
rect 32680 24890 32732 24896
rect 32588 24880 32640 24886
rect 32588 24822 32640 24828
rect 32772 24812 32824 24818
rect 32772 24754 32824 24760
rect 32588 24744 32640 24750
rect 32588 24686 32640 24692
rect 32600 24188 32628 24686
rect 32680 24200 32732 24206
rect 32600 24160 32680 24188
rect 32680 24142 32732 24148
rect 32496 24064 32548 24070
rect 32548 24012 32628 24018
rect 32496 24006 32628 24012
rect 32508 23990 32628 24006
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32036 23180 32088 23186
rect 32036 23122 32088 23128
rect 32220 23180 32272 23186
rect 32220 23122 32272 23128
rect 31760 23044 31812 23050
rect 31760 22986 31812 22992
rect 31772 22778 31800 22986
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 31852 22500 31904 22506
rect 31772 22460 31852 22488
rect 31772 22166 31800 22460
rect 31852 22442 31904 22448
rect 31760 22160 31812 22166
rect 31760 22102 31812 22108
rect 31772 21570 31800 22102
rect 31772 21542 31984 21570
rect 31852 21480 31904 21486
rect 31852 21422 31904 21428
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31772 19718 31800 20878
rect 31864 20806 31892 21422
rect 31852 20800 31904 20806
rect 31852 20742 31904 20748
rect 31956 20058 31984 21542
rect 31944 20052 31996 20058
rect 31944 19994 31996 20000
rect 31760 19712 31812 19718
rect 31760 19654 31812 19660
rect 31576 19508 31628 19514
rect 31576 19450 31628 19456
rect 31588 18766 31616 19450
rect 31772 18766 31800 19654
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 31760 18760 31812 18766
rect 31760 18702 31812 18708
rect 31576 18284 31628 18290
rect 31576 18226 31628 18232
rect 31392 16516 31444 16522
rect 31392 16458 31444 16464
rect 31404 16250 31432 16458
rect 31392 16244 31444 16250
rect 31392 16186 31444 16192
rect 31300 15564 31352 15570
rect 31300 15506 31352 15512
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 31036 15094 31064 15302
rect 31024 15088 31076 15094
rect 31024 15030 31076 15036
rect 31588 14890 31616 18226
rect 31772 17746 31800 18702
rect 31944 18420 31996 18426
rect 31944 18362 31996 18368
rect 31760 17740 31812 17746
rect 31760 17682 31812 17688
rect 31772 16658 31800 17682
rect 31956 17202 31984 18362
rect 32048 17354 32076 23122
rect 32128 22976 32180 22982
rect 32128 22918 32180 22924
rect 32140 22642 32168 22918
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 32140 20942 32168 21966
rect 32404 21956 32456 21962
rect 32404 21898 32456 21904
rect 32416 21690 32444 21898
rect 32508 21894 32536 22714
rect 32496 21888 32548 21894
rect 32496 21830 32548 21836
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 32496 21548 32548 21554
rect 32496 21490 32548 21496
rect 32128 20936 32180 20942
rect 32128 20878 32180 20884
rect 32508 20806 32536 21490
rect 32600 21418 32628 23990
rect 32784 23662 32812 24754
rect 32772 23656 32824 23662
rect 32772 23598 32824 23604
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32588 21412 32640 21418
rect 32588 21354 32640 21360
rect 32312 20800 32364 20806
rect 32312 20742 32364 20748
rect 32496 20800 32548 20806
rect 32496 20742 32548 20748
rect 32128 20392 32180 20398
rect 32128 20334 32180 20340
rect 32140 19514 32168 20334
rect 32128 19508 32180 19514
rect 32128 19450 32180 19456
rect 32048 17326 32168 17354
rect 32036 17264 32088 17270
rect 32036 17206 32088 17212
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 31956 17105 31984 17138
rect 31942 17096 31998 17105
rect 31852 17060 31904 17066
rect 31942 17031 31998 17040
rect 31852 17002 31904 17008
rect 31760 16652 31812 16658
rect 31760 16594 31812 16600
rect 31760 16516 31812 16522
rect 31864 16504 31892 17002
rect 31944 16652 31996 16658
rect 31944 16594 31996 16600
rect 31812 16476 31892 16504
rect 31760 16458 31812 16464
rect 31668 16108 31720 16114
rect 31668 16050 31720 16056
rect 31680 15162 31708 16050
rect 31772 15502 31800 16458
rect 31956 16114 31984 16594
rect 32048 16522 32076 17206
rect 32036 16516 32088 16522
rect 32036 16458 32088 16464
rect 31944 16108 31996 16114
rect 31944 16050 31996 16056
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31852 15496 31904 15502
rect 31852 15438 31904 15444
rect 31864 15162 31892 15438
rect 31668 15156 31720 15162
rect 31668 15098 31720 15104
rect 31852 15156 31904 15162
rect 31852 15098 31904 15104
rect 31576 14884 31628 14890
rect 31496 14844 31576 14872
rect 31116 12776 31168 12782
rect 31116 12718 31168 12724
rect 31128 12442 31156 12718
rect 31496 12646 31524 14844
rect 31576 14826 31628 14832
rect 31956 14482 31984 16050
rect 31944 14476 31996 14482
rect 31944 14418 31996 14424
rect 31852 14340 31904 14346
rect 31852 14282 31904 14288
rect 31864 12782 31892 14282
rect 32140 13870 32168 17326
rect 32220 16448 32272 16454
rect 32220 16390 32272 16396
rect 32232 16182 32260 16390
rect 32220 16176 32272 16182
rect 32220 16118 32272 16124
rect 32220 14816 32272 14822
rect 32220 14758 32272 14764
rect 32232 14482 32260 14758
rect 32220 14476 32272 14482
rect 32220 14418 32272 14424
rect 32128 13864 32180 13870
rect 32128 13806 32180 13812
rect 32140 13274 32168 13806
rect 32324 13802 32352 20742
rect 32404 20596 32456 20602
rect 32404 20538 32456 20544
rect 32416 18290 32444 20538
rect 32588 19508 32640 19514
rect 32588 19450 32640 19456
rect 32600 18766 32628 19450
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 32600 18358 32628 18702
rect 32588 18352 32640 18358
rect 32588 18294 32640 18300
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32416 14074 32444 18226
rect 32496 16992 32548 16998
rect 32496 16934 32548 16940
rect 32508 16794 32536 16934
rect 32496 16788 32548 16794
rect 32496 16730 32548 16736
rect 32404 14068 32456 14074
rect 32404 14010 32456 14016
rect 32312 13796 32364 13802
rect 32312 13738 32364 13744
rect 32416 13530 32444 14010
rect 32404 13524 32456 13530
rect 32404 13466 32456 13472
rect 32140 13246 32260 13274
rect 32128 13184 32180 13190
rect 32128 13126 32180 13132
rect 31576 12776 31628 12782
rect 31576 12718 31628 12724
rect 31852 12776 31904 12782
rect 31852 12718 31904 12724
rect 31484 12640 31536 12646
rect 31484 12582 31536 12588
rect 31116 12436 31168 12442
rect 31588 12434 31616 12718
rect 31588 12406 31708 12434
rect 31116 12378 31168 12384
rect 31680 12306 31708 12406
rect 31668 12300 31720 12306
rect 31668 12242 31720 12248
rect 31024 12164 31076 12170
rect 31024 12106 31076 12112
rect 30932 11892 30984 11898
rect 30932 11834 30984 11840
rect 31036 11762 31064 12106
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 31392 11688 31444 11694
rect 31392 11630 31444 11636
rect 31576 11688 31628 11694
rect 31576 11630 31628 11636
rect 31404 11354 31432 11630
rect 31392 11348 31444 11354
rect 31392 11290 31444 11296
rect 31588 11286 31616 11630
rect 31576 11280 31628 11286
rect 31576 11222 31628 11228
rect 31680 11218 31708 12242
rect 31850 11928 31906 11937
rect 31850 11863 31906 11872
rect 31864 11830 31892 11863
rect 31852 11824 31904 11830
rect 31852 11766 31904 11772
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 31680 11098 31708 11154
rect 31864 11150 31892 11766
rect 32036 11620 32088 11626
rect 32036 11562 32088 11568
rect 31852 11144 31904 11150
rect 31680 11070 31800 11098
rect 31852 11086 31904 11092
rect 32048 11082 32076 11562
rect 30840 10736 30892 10742
rect 30840 10678 30892 10684
rect 30852 9586 30880 10678
rect 31772 10130 31800 11070
rect 32036 11076 32088 11082
rect 32036 11018 32088 11024
rect 31944 11008 31996 11014
rect 31944 10950 31996 10956
rect 31208 10124 31260 10130
rect 31208 10066 31260 10072
rect 31760 10124 31812 10130
rect 31760 10066 31812 10072
rect 31220 9722 31248 10066
rect 31208 9716 31260 9722
rect 31208 9658 31260 9664
rect 31772 9654 31800 10066
rect 31956 9994 31984 10950
rect 31944 9988 31996 9994
rect 31944 9930 31996 9936
rect 31760 9648 31812 9654
rect 31760 9590 31812 9596
rect 30840 9580 30892 9586
rect 30840 9522 30892 9528
rect 30840 9376 30892 9382
rect 30760 9336 30840 9364
rect 30840 9318 30892 9324
rect 31852 8900 31904 8906
rect 31852 8842 31904 8848
rect 31760 8492 31812 8498
rect 31680 8452 31760 8480
rect 31680 8022 31708 8452
rect 31760 8434 31812 8440
rect 31668 8016 31720 8022
rect 31668 7958 31720 7964
rect 31576 7948 31628 7954
rect 31576 7890 31628 7896
rect 31300 7880 31352 7886
rect 31220 7840 31300 7868
rect 31024 7812 31076 7818
rect 31024 7754 31076 7760
rect 31036 7546 31064 7754
rect 31024 7540 31076 7546
rect 31024 7482 31076 7488
rect 30656 7404 30708 7410
rect 30656 7346 30708 7352
rect 30932 7404 30984 7410
rect 30932 7346 30984 7352
rect 30668 6390 30696 7346
rect 30840 6996 30892 7002
rect 30840 6938 30892 6944
rect 30656 6384 30708 6390
rect 30656 6326 30708 6332
rect 30852 6322 30880 6938
rect 30944 6866 30972 7346
rect 31024 7336 31076 7342
rect 31024 7278 31076 7284
rect 31036 7206 31064 7278
rect 31024 7200 31076 7206
rect 31024 7142 31076 7148
rect 30932 6860 30984 6866
rect 30932 6802 30984 6808
rect 31036 6730 31064 7142
rect 31220 6866 31248 7840
rect 31300 7822 31352 7828
rect 31588 7478 31616 7890
rect 31392 7472 31444 7478
rect 31392 7414 31444 7420
rect 31576 7472 31628 7478
rect 31576 7414 31628 7420
rect 31404 7342 31432 7414
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31392 7336 31444 7342
rect 31392 7278 31444 7284
rect 31208 6860 31260 6866
rect 31208 6802 31260 6808
rect 31024 6724 31076 6730
rect 31024 6666 31076 6672
rect 30840 6316 30892 6322
rect 30840 6258 30892 6264
rect 30012 6190 30064 6196
rect 29552 5636 29604 5642
rect 29552 5578 29604 5584
rect 28724 5296 28776 5302
rect 28724 5238 28776 5244
rect 29564 5234 29592 5578
rect 29932 5370 29960 6190
rect 30484 6174 30696 6202
rect 30484 6118 30512 6174
rect 30472 6112 30524 6118
rect 30472 6054 30524 6060
rect 30564 6112 30616 6118
rect 30564 6054 30616 6060
rect 30576 5778 30604 6054
rect 30564 5772 30616 5778
rect 30564 5714 30616 5720
rect 29920 5364 29972 5370
rect 29920 5306 29972 5312
rect 30668 5302 30696 6174
rect 30748 6112 30800 6118
rect 30748 6054 30800 6060
rect 30760 5574 30788 6054
rect 30852 5574 30880 6258
rect 31220 5710 31248 6802
rect 31312 6798 31340 7278
rect 31404 6798 31432 7278
rect 31588 6934 31616 7414
rect 31760 7404 31812 7410
rect 31760 7346 31812 7352
rect 31772 7002 31800 7346
rect 31760 6996 31812 7002
rect 31760 6938 31812 6944
rect 31576 6928 31628 6934
rect 31576 6870 31628 6876
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31392 6792 31444 6798
rect 31392 6734 31444 6740
rect 31312 6662 31340 6734
rect 31300 6656 31352 6662
rect 31300 6598 31352 6604
rect 31312 6322 31340 6598
rect 31864 6458 31892 8842
rect 32140 7886 32168 13126
rect 32232 12986 32260 13246
rect 32220 12980 32272 12986
rect 32220 12922 32272 12928
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32324 12170 32352 12582
rect 32312 12164 32364 12170
rect 32312 12106 32364 12112
rect 32312 11008 32364 11014
rect 32312 10950 32364 10956
rect 32324 10674 32352 10950
rect 32312 10668 32364 10674
rect 32312 10610 32364 10616
rect 32220 10124 32272 10130
rect 32220 10066 32272 10072
rect 32232 9178 32260 10066
rect 32416 9654 32444 13466
rect 32588 12232 32640 12238
rect 32588 12174 32640 12180
rect 32494 12064 32550 12073
rect 32494 11999 32550 12008
rect 32508 11626 32536 11999
rect 32600 11898 32628 12174
rect 32692 12170 32720 22578
rect 32772 20800 32824 20806
rect 32772 20742 32824 20748
rect 32784 20534 32812 20742
rect 32772 20528 32824 20534
rect 32772 20470 32824 20476
rect 32876 19922 32904 25638
rect 33048 24948 33100 24954
rect 33048 24890 33100 24896
rect 32956 24812 33008 24818
rect 32956 24754 33008 24760
rect 32968 24410 32996 24754
rect 32956 24404 33008 24410
rect 32956 24346 33008 24352
rect 33060 24274 33088 24890
rect 33140 24676 33192 24682
rect 33140 24618 33192 24624
rect 33152 24410 33180 24618
rect 33508 24608 33560 24614
rect 33508 24550 33560 24556
rect 33140 24404 33192 24410
rect 33140 24346 33192 24352
rect 33520 24342 33548 24550
rect 33612 24410 33640 26318
rect 33784 26308 33836 26314
rect 33784 26250 33836 26256
rect 33796 26042 33824 26250
rect 33784 26036 33836 26042
rect 33784 25978 33836 25984
rect 33784 25696 33836 25702
rect 33888 25684 33916 26522
rect 33980 26489 34008 27288
rect 34256 27305 34284 28863
rect 34348 28762 34376 29174
rect 34440 29102 34468 29650
rect 34428 29096 34480 29102
rect 34428 29038 34480 29044
rect 34336 28756 34388 28762
rect 34336 28698 34388 28704
rect 34348 28150 34376 28698
rect 34440 28626 34468 29038
rect 34428 28620 34480 28626
rect 34428 28562 34480 28568
rect 34336 28144 34388 28150
rect 34336 28086 34388 28092
rect 34428 28144 34480 28150
rect 34428 28086 34480 28092
rect 34532 28098 34560 30110
rect 34624 29850 34652 30126
rect 34612 29844 34664 29850
rect 34612 29786 34664 29792
rect 34610 29336 34666 29345
rect 34610 29271 34666 29280
rect 34624 28490 34652 29271
rect 34716 28694 34744 30262
rect 35360 30240 35388 30602
rect 35452 30394 35480 30654
rect 35714 30631 35770 30640
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 35440 30388 35492 30394
rect 35440 30330 35492 30336
rect 36360 30388 36412 30394
rect 36360 30330 36412 30336
rect 35992 30252 36044 30258
rect 35360 30212 35572 30240
rect 34796 30048 34848 30054
rect 34796 29990 34848 29996
rect 34799 29832 34827 29990
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34799 29804 34928 29832
rect 34796 29572 34848 29578
rect 34796 29514 34848 29520
rect 34808 29481 34836 29514
rect 34794 29472 34850 29481
rect 34794 29407 34850 29416
rect 34900 29170 34928 29804
rect 34980 29708 35032 29714
rect 35360 29696 35388 30212
rect 35438 30152 35494 30161
rect 35438 30087 35494 30096
rect 34980 29650 35032 29656
rect 35268 29668 35388 29696
rect 34992 29345 35020 29650
rect 35268 29481 35296 29668
rect 35452 29646 35480 30087
rect 35544 29782 35572 30212
rect 35992 30194 36044 30200
rect 36176 30252 36228 30258
rect 36176 30194 36228 30200
rect 36268 30252 36320 30258
rect 36268 30194 36320 30200
rect 35808 30184 35860 30190
rect 35728 30132 35808 30138
rect 35728 30126 35860 30132
rect 35728 30110 35848 30126
rect 35624 30048 35676 30054
rect 35624 29990 35676 29996
rect 35532 29776 35584 29782
rect 35532 29718 35584 29724
rect 35636 29646 35664 29990
rect 35440 29640 35492 29646
rect 35360 29588 35440 29594
rect 35360 29582 35492 29588
rect 35624 29640 35676 29646
rect 35624 29582 35676 29588
rect 35360 29566 35480 29582
rect 35254 29472 35310 29481
rect 35254 29407 35310 29416
rect 34978 29336 35034 29345
rect 34978 29271 35034 29280
rect 34888 29164 34940 29170
rect 34888 29106 34940 29112
rect 35360 29073 35388 29566
rect 35728 29510 35756 30110
rect 35900 30048 35952 30054
rect 35900 29990 35952 29996
rect 35912 29646 35940 29990
rect 36004 29850 36032 30194
rect 35992 29844 36044 29850
rect 35992 29786 36044 29792
rect 36084 29844 36136 29850
rect 36084 29786 36136 29792
rect 35900 29640 35952 29646
rect 35900 29582 35952 29588
rect 35532 29504 35584 29510
rect 35452 29464 35532 29492
rect 35346 29064 35402 29073
rect 35256 29028 35308 29034
rect 35346 28999 35402 29008
rect 35256 28970 35308 28976
rect 34796 28960 34848 28966
rect 34796 28902 34848 28908
rect 35268 28914 35296 28970
rect 34808 28762 34836 28902
rect 35268 28886 35388 28914
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28756 34848 28762
rect 34796 28698 34848 28704
rect 34704 28688 34756 28694
rect 35360 28642 35388 28886
rect 34704 28630 34756 28636
rect 35176 28614 35388 28642
rect 34612 28484 34664 28490
rect 34612 28426 34664 28432
rect 34348 27538 34376 28086
rect 34336 27532 34388 27538
rect 34336 27474 34388 27480
rect 34440 27470 34468 28086
rect 34532 28070 34836 28098
rect 34704 28008 34756 28014
rect 34704 27950 34756 27956
rect 34520 27872 34572 27878
rect 34520 27814 34572 27820
rect 34612 27872 34664 27878
rect 34612 27814 34664 27820
rect 34428 27464 34480 27470
rect 34428 27406 34480 27412
rect 34060 27270 34112 27276
rect 34242 27296 34298 27305
rect 34072 26926 34100 27270
rect 34242 27231 34298 27240
rect 34060 26920 34112 26926
rect 34060 26862 34112 26868
rect 34150 26888 34206 26897
rect 34150 26823 34206 26832
rect 34164 26586 34192 26823
rect 34256 26586 34284 27231
rect 34440 27130 34468 27406
rect 34428 27124 34480 27130
rect 34428 27066 34480 27072
rect 34152 26580 34204 26586
rect 34152 26522 34204 26528
rect 34244 26580 34296 26586
rect 34244 26522 34296 26528
rect 33966 26480 34022 26489
rect 33966 26415 34022 26424
rect 34440 26382 34468 27066
rect 34532 27062 34560 27814
rect 34624 27538 34652 27814
rect 34612 27532 34664 27538
rect 34612 27474 34664 27480
rect 34716 27334 34744 27950
rect 34704 27328 34756 27334
rect 34704 27270 34756 27276
rect 34610 27160 34666 27169
rect 34610 27095 34666 27104
rect 34520 27056 34572 27062
rect 34520 26998 34572 27004
rect 34520 26920 34572 26926
rect 34520 26862 34572 26868
rect 34428 26376 34480 26382
rect 34428 26318 34480 26324
rect 33836 25656 33916 25684
rect 33784 25638 33836 25644
rect 33796 25226 33824 25638
rect 34532 25362 34560 26862
rect 34624 26790 34652 27095
rect 34612 26784 34664 26790
rect 34612 26726 34664 26732
rect 34624 26314 34652 26726
rect 34808 26314 34836 28070
rect 35176 27878 35204 28614
rect 35348 28416 35400 28422
rect 35348 28358 35400 28364
rect 35164 27872 35216 27878
rect 35164 27814 35216 27820
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27606 35388 28358
rect 35348 27600 35400 27606
rect 35348 27542 35400 27548
rect 35256 27464 35308 27470
rect 35256 27406 35308 27412
rect 35268 26858 35296 27406
rect 35256 26852 35308 26858
rect 35256 26794 35308 26800
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34612 26308 34664 26314
rect 34612 26250 34664 26256
rect 34796 26308 34848 26314
rect 34796 26250 34848 26256
rect 34808 25514 34836 26250
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34716 25486 34836 25514
rect 34520 25356 34572 25362
rect 34520 25298 34572 25304
rect 33784 25220 33836 25226
rect 33784 25162 33836 25168
rect 34244 25220 34296 25226
rect 34244 25162 34296 25168
rect 34520 25220 34572 25226
rect 34520 25162 34572 25168
rect 34256 24954 34284 25162
rect 34244 24948 34296 24954
rect 34244 24890 34296 24896
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33704 24682 33732 24754
rect 34532 24750 34560 25162
rect 34520 24744 34572 24750
rect 34520 24686 34572 24692
rect 33692 24676 33744 24682
rect 33692 24618 33744 24624
rect 33600 24404 33652 24410
rect 33600 24346 33652 24352
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 32956 24268 33008 24274
rect 32956 24210 33008 24216
rect 33048 24268 33100 24274
rect 33048 24210 33100 24216
rect 32968 24070 32996 24210
rect 32956 24064 33008 24070
rect 32956 24006 33008 24012
rect 33416 23112 33468 23118
rect 33416 23054 33468 23060
rect 33508 23112 33560 23118
rect 33508 23054 33560 23060
rect 33428 22778 33456 23054
rect 33520 22778 33548 23054
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33508 22772 33560 22778
rect 33508 22714 33560 22720
rect 33232 22704 33284 22710
rect 33232 22646 33284 22652
rect 33140 22024 33192 22030
rect 33140 21966 33192 21972
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 33060 21622 33088 21830
rect 33048 21616 33100 21622
rect 33048 21558 33100 21564
rect 33152 21350 33180 21966
rect 33140 21344 33192 21350
rect 33140 21286 33192 21292
rect 33152 20466 33180 21286
rect 33140 20460 33192 20466
rect 33140 20402 33192 20408
rect 33048 20052 33100 20058
rect 33048 19994 33100 20000
rect 33060 19922 33088 19994
rect 32864 19916 32916 19922
rect 32864 19858 32916 19864
rect 33048 19916 33100 19922
rect 33048 19858 33100 19864
rect 33060 15570 33088 19858
rect 33140 19440 33192 19446
rect 33244 19394 33272 22646
rect 33428 22094 33456 22714
rect 33336 22066 33456 22094
rect 33336 20534 33364 22066
rect 33416 21956 33468 21962
rect 33416 21898 33468 21904
rect 33428 21554 33456 21898
rect 33508 21888 33560 21894
rect 33506 21856 33508 21865
rect 33560 21856 33562 21865
rect 33506 21791 33562 21800
rect 33416 21548 33468 21554
rect 33416 21490 33468 21496
rect 33324 20528 33376 20534
rect 33324 20470 33376 20476
rect 33192 19388 33364 19394
rect 33140 19382 33364 19388
rect 33152 19366 33364 19382
rect 33232 19168 33284 19174
rect 33232 19110 33284 19116
rect 33140 18692 33192 18698
rect 33140 18634 33192 18640
rect 33152 18426 33180 18634
rect 33140 18420 33192 18426
rect 33140 18362 33192 18368
rect 33244 17354 33272 19110
rect 33336 18834 33364 19366
rect 33324 18828 33376 18834
rect 33324 18770 33376 18776
rect 33336 17814 33364 18770
rect 33324 17808 33376 17814
rect 33324 17750 33376 17756
rect 33152 17326 33272 17354
rect 33048 15564 33100 15570
rect 33048 15506 33100 15512
rect 32772 15428 32824 15434
rect 32772 15370 32824 15376
rect 32784 15162 32812 15370
rect 32772 15156 32824 15162
rect 32772 15098 32824 15104
rect 33152 14958 33180 17326
rect 33232 17196 33284 17202
rect 33232 17138 33284 17144
rect 33244 16522 33272 17138
rect 33324 16992 33376 16998
rect 33324 16934 33376 16940
rect 33336 16658 33364 16934
rect 33324 16652 33376 16658
rect 33324 16594 33376 16600
rect 33232 16516 33284 16522
rect 33232 16458 33284 16464
rect 33140 14952 33192 14958
rect 33140 14894 33192 14900
rect 32956 14340 33008 14346
rect 32956 14282 33008 14288
rect 32968 14006 32996 14282
rect 33048 14068 33100 14074
rect 33048 14010 33100 14016
rect 32956 14000 33008 14006
rect 32876 13960 32956 13988
rect 32680 12164 32732 12170
rect 32680 12106 32732 12112
rect 32588 11892 32640 11898
rect 32588 11834 32640 11840
rect 32496 11620 32548 11626
rect 32496 11562 32548 11568
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32508 10810 32536 11086
rect 32692 10810 32720 12106
rect 32876 12102 32904 13960
rect 32956 13942 33008 13948
rect 32956 13796 33008 13802
rect 32956 13738 33008 13744
rect 32968 12442 32996 13738
rect 33060 13394 33088 14010
rect 33048 13388 33100 13394
rect 33048 13330 33100 13336
rect 33152 12782 33180 14894
rect 33428 12986 33456 21490
rect 33508 20392 33560 20398
rect 33508 20334 33560 20340
rect 33520 17678 33548 20334
rect 33612 18970 33640 24346
rect 34532 24070 34560 24686
rect 34612 24404 34664 24410
rect 34612 24346 34664 24352
rect 34624 24206 34652 24346
rect 34612 24200 34664 24206
rect 34612 24142 34664 24148
rect 34520 24064 34572 24070
rect 34520 24006 34572 24012
rect 34716 23798 34744 25486
rect 34796 25356 34848 25362
rect 34796 25298 34848 25304
rect 34808 24138 34836 25298
rect 35256 25288 35308 25294
rect 35162 25256 35218 25265
rect 35256 25230 35308 25236
rect 35162 25191 35218 25200
rect 35176 24818 35204 25191
rect 35268 24954 35296 25230
rect 35348 25152 35400 25158
rect 35348 25094 35400 25100
rect 35256 24948 35308 24954
rect 35256 24890 35308 24896
rect 35164 24812 35216 24818
rect 35164 24754 35216 24760
rect 35268 24562 35296 24890
rect 35360 24818 35388 25094
rect 35348 24812 35400 24818
rect 35452 24808 35480 29464
rect 35532 29446 35584 29452
rect 35716 29504 35768 29510
rect 35716 29446 35768 29452
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 35532 29164 35584 29170
rect 35532 29106 35584 29112
rect 35900 29164 35952 29170
rect 35900 29106 35952 29112
rect 35544 28694 35572 29106
rect 35624 29096 35676 29102
rect 35624 29038 35676 29044
rect 35806 29064 35862 29073
rect 35532 28688 35584 28694
rect 35532 28630 35584 28636
rect 35636 28404 35664 29038
rect 35806 28999 35808 29008
rect 35860 28999 35862 29008
rect 35808 28970 35860 28976
rect 35912 28558 35940 29106
rect 36004 29034 36032 29786
rect 35992 29028 36044 29034
rect 35992 28970 36044 28976
rect 35716 28552 35768 28558
rect 35900 28552 35952 28558
rect 35768 28512 35900 28540
rect 35716 28494 35768 28500
rect 35900 28494 35952 28500
rect 35636 28376 36032 28404
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 35532 27872 35584 27878
rect 35532 27814 35584 27820
rect 35544 27674 35572 27814
rect 36004 27674 36032 28376
rect 36096 28121 36124 29786
rect 36188 29753 36216 30194
rect 36280 30054 36308 30194
rect 36268 30048 36320 30054
rect 36268 29990 36320 29996
rect 36174 29744 36230 29753
rect 36230 29702 36308 29730
rect 36174 29679 36230 29688
rect 36176 29504 36228 29510
rect 36174 29472 36176 29481
rect 36228 29472 36230 29481
rect 36174 29407 36230 29416
rect 36176 29164 36228 29170
rect 36176 29106 36228 29112
rect 36188 28762 36216 29106
rect 36176 28756 36228 28762
rect 36176 28698 36228 28704
rect 36082 28112 36138 28121
rect 36082 28047 36138 28056
rect 35532 27668 35584 27674
rect 35532 27610 35584 27616
rect 35992 27668 36044 27674
rect 35992 27610 36044 27616
rect 35544 27538 35572 27610
rect 36004 27554 36032 27610
rect 35532 27532 35584 27538
rect 35532 27474 35584 27480
rect 35912 27526 36032 27554
rect 35532 27396 35584 27402
rect 35912 27384 35940 27526
rect 35992 27464 36044 27470
rect 35992 27406 36044 27412
rect 35584 27356 35940 27384
rect 35532 27338 35584 27344
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35808 27124 35860 27130
rect 36004 27112 36032 27406
rect 35860 27084 36032 27112
rect 35808 27066 35860 27072
rect 35532 27056 35584 27062
rect 35532 26998 35584 27004
rect 35544 26761 35572 26998
rect 35624 26988 35676 26994
rect 35624 26930 35676 26936
rect 35530 26752 35586 26761
rect 35530 26687 35586 26696
rect 35636 26625 35664 26930
rect 35716 26852 35768 26858
rect 35716 26794 35768 26800
rect 35622 26616 35678 26625
rect 35622 26551 35678 26560
rect 35728 26450 35756 26794
rect 36096 26790 36124 28047
rect 36280 27130 36308 29702
rect 36372 29646 36400 30330
rect 36740 30326 36768 33390
rect 36820 31680 36872 31686
rect 36820 31622 36872 31628
rect 36832 30734 36860 31622
rect 36820 30728 36872 30734
rect 36820 30670 36872 30676
rect 36728 30320 36780 30326
rect 36728 30262 36780 30268
rect 36452 30252 36504 30258
rect 36452 30194 36504 30200
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 36636 30252 36688 30258
rect 36636 30194 36688 30200
rect 36360 29640 36412 29646
rect 36360 29582 36412 29588
rect 36372 29306 36400 29582
rect 36360 29300 36412 29306
rect 36360 29242 36412 29248
rect 36372 28994 36400 29242
rect 36464 29102 36492 30194
rect 36556 30054 36584 30194
rect 36648 30161 36676 30194
rect 36634 30152 36690 30161
rect 36634 30087 36690 30096
rect 36544 30048 36596 30054
rect 36544 29990 36596 29996
rect 36452 29096 36504 29102
rect 36452 29038 36504 29044
rect 36372 28966 36492 28994
rect 36268 27124 36320 27130
rect 36268 27066 36320 27072
rect 36358 27024 36414 27033
rect 36176 26988 36228 26994
rect 36464 26994 36492 28966
rect 36556 28558 36584 29990
rect 36740 29646 36768 30262
rect 36820 29708 36872 29714
rect 36820 29650 36872 29656
rect 36728 29640 36780 29646
rect 36728 29582 36780 29588
rect 36634 29472 36690 29481
rect 36634 29407 36690 29416
rect 36544 28552 36596 28558
rect 36544 28494 36596 28500
rect 36648 27418 36676 29407
rect 36832 29238 36860 29650
rect 36910 29608 36966 29617
rect 36910 29543 36966 29552
rect 36924 29306 36952 29543
rect 36912 29300 36964 29306
rect 36912 29242 36964 29248
rect 36820 29232 36872 29238
rect 36820 29174 36872 29180
rect 36820 29096 36872 29102
rect 36820 29038 36872 29044
rect 36556 27390 36676 27418
rect 36556 27062 36584 27390
rect 36636 27328 36688 27334
rect 36636 27270 36688 27276
rect 36648 27130 36676 27270
rect 36636 27124 36688 27130
rect 36636 27066 36688 27072
rect 36544 27056 36596 27062
rect 36544 26998 36596 27004
rect 36358 26959 36360 26968
rect 36176 26930 36228 26936
rect 36412 26959 36414 26968
rect 36452 26988 36504 26994
rect 36360 26930 36412 26936
rect 36452 26930 36504 26936
rect 36084 26784 36136 26790
rect 36084 26726 36136 26732
rect 35716 26444 35768 26450
rect 35716 26386 35768 26392
rect 36084 26376 36136 26382
rect 36188 26364 36216 26930
rect 36372 26382 36400 26930
rect 36464 26382 36492 26930
rect 36556 26625 36584 26998
rect 36728 26920 36780 26926
rect 36728 26862 36780 26868
rect 36542 26616 36598 26625
rect 36542 26551 36598 26560
rect 36740 26382 36768 26862
rect 36832 26382 36860 29038
rect 36912 29028 36964 29034
rect 36912 28970 36964 28976
rect 36136 26336 36216 26364
rect 36360 26376 36412 26382
rect 36084 26318 36136 26324
rect 36360 26318 36412 26324
rect 36452 26376 36504 26382
rect 36452 26318 36504 26324
rect 36728 26376 36780 26382
rect 36728 26318 36780 26324
rect 36820 26376 36872 26382
rect 36820 26318 36872 26324
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35992 25288 36044 25294
rect 35898 25256 35954 25265
rect 35992 25230 36044 25236
rect 35898 25191 35900 25200
rect 35952 25191 35954 25200
rect 35900 25162 35952 25168
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35636 24818 35940 24834
rect 35624 24812 35940 24818
rect 35348 24754 35400 24760
rect 35440 24802 35492 24808
rect 35676 24806 35940 24812
rect 35624 24754 35676 24760
rect 35440 24744 35492 24750
rect 35624 24608 35676 24614
rect 35268 24534 35388 24562
rect 35624 24550 35676 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24426 35388 24534
rect 35268 24398 35388 24426
rect 34980 24200 35032 24206
rect 35268 24154 35296 24398
rect 35636 24206 35664 24550
rect 35912 24274 35940 24806
rect 36004 24274 36032 25230
rect 35900 24268 35952 24274
rect 35900 24210 35952 24216
rect 35992 24268 36044 24274
rect 35992 24210 36044 24216
rect 34980 24142 35032 24148
rect 34796 24132 34848 24138
rect 34796 24074 34848 24080
rect 34992 23866 35020 24142
rect 35176 24138 35296 24154
rect 35624 24200 35676 24206
rect 35624 24142 35676 24148
rect 35912 24154 35940 24210
rect 35164 24132 35296 24138
rect 35216 24126 35296 24132
rect 35912 24126 36032 24154
rect 36096 24138 36124 26318
rect 36268 26308 36320 26314
rect 36268 26250 36320 26256
rect 36280 26042 36308 26250
rect 36464 26246 36492 26318
rect 36452 26240 36504 26246
rect 36452 26182 36504 26188
rect 36268 26036 36320 26042
rect 36268 25978 36320 25984
rect 36188 25486 36492 25514
rect 36188 25362 36216 25486
rect 36464 25362 36492 25486
rect 36176 25356 36228 25362
rect 36176 25298 36228 25304
rect 36452 25356 36504 25362
rect 36452 25298 36504 25304
rect 36544 25288 36596 25294
rect 36544 25230 36596 25236
rect 36268 25220 36320 25226
rect 36268 25162 36320 25168
rect 36280 24886 36308 25162
rect 36556 24886 36584 25230
rect 36268 24880 36320 24886
rect 36268 24822 36320 24828
rect 36544 24880 36596 24886
rect 36544 24822 36596 24828
rect 36176 24744 36228 24750
rect 36176 24686 36228 24692
rect 36452 24744 36504 24750
rect 36452 24686 36504 24692
rect 35164 24074 35216 24080
rect 34980 23860 35032 23866
rect 34980 23802 35032 23808
rect 35176 23798 35204 24074
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 34704 23792 34756 23798
rect 34704 23734 34756 23740
rect 35164 23792 35216 23798
rect 35164 23734 35216 23740
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 34532 23186 34560 23598
rect 34520 23180 34572 23186
rect 34520 23122 34572 23128
rect 34624 23066 34652 23666
rect 34716 23254 34744 23734
rect 34980 23724 35032 23730
rect 34980 23666 35032 23672
rect 35440 23724 35492 23730
rect 35440 23666 35492 23672
rect 34992 23526 35020 23666
rect 34796 23520 34848 23526
rect 34796 23462 34848 23468
rect 34980 23520 35032 23526
rect 34980 23462 35032 23468
rect 34704 23248 34756 23254
rect 34704 23190 34756 23196
rect 34808 23202 34836 23462
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34532 23038 34652 23066
rect 34716 23066 34744 23190
rect 34808 23174 35112 23202
rect 34716 23038 35020 23066
rect 34060 22228 34112 22234
rect 34060 22170 34112 22176
rect 34072 21554 34100 22170
rect 34532 22094 34560 23038
rect 34992 22982 35020 23038
rect 34612 22976 34664 22982
rect 34612 22918 34664 22924
rect 34888 22976 34940 22982
rect 34888 22918 34940 22924
rect 34980 22976 35032 22982
rect 34980 22918 35032 22924
rect 34624 22234 34652 22918
rect 34900 22710 34928 22918
rect 34888 22704 34940 22710
rect 34888 22646 34940 22652
rect 35084 22658 35112 23174
rect 35256 23112 35308 23118
rect 35256 23054 35308 23060
rect 35268 22778 35296 23054
rect 35256 22772 35308 22778
rect 35256 22714 35308 22720
rect 35084 22630 35388 22658
rect 35452 22642 35480 23666
rect 35716 23588 35768 23594
rect 35716 23530 35768 23536
rect 35530 23216 35586 23225
rect 35728 23186 35756 23530
rect 36004 23186 36032 24126
rect 36084 24132 36136 24138
rect 36084 24074 36136 24080
rect 35530 23151 35532 23160
rect 35584 23151 35586 23160
rect 35716 23180 35768 23186
rect 35532 23122 35584 23128
rect 35716 23122 35768 23128
rect 35992 23180 36044 23186
rect 35992 23122 36044 23128
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35360 22574 35388 22630
rect 35440 22636 35492 22642
rect 35440 22578 35492 22584
rect 34796 22568 34848 22574
rect 34796 22510 34848 22516
rect 35348 22568 35400 22574
rect 35348 22510 35400 22516
rect 34612 22228 34664 22234
rect 34612 22170 34664 22176
rect 34808 22098 34836 22510
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34532 22066 34744 22094
rect 34428 22024 34480 22030
rect 34428 21966 34480 21972
rect 34060 21548 34112 21554
rect 34060 21490 34112 21496
rect 33692 21480 33744 21486
rect 33692 21422 33744 21428
rect 34440 21434 34468 21966
rect 34716 21962 34744 22066
rect 34796 22092 34848 22098
rect 34796 22034 34848 22040
rect 34704 21956 34756 21962
rect 34704 21898 34756 21904
rect 35072 21956 35124 21962
rect 35072 21898 35124 21904
rect 35084 21690 35112 21898
rect 35072 21684 35124 21690
rect 35072 21626 35124 21632
rect 35360 21622 35388 22510
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 35348 21616 35400 21622
rect 35348 21558 35400 21564
rect 34612 21548 34664 21554
rect 34612 21490 34664 21496
rect 34624 21434 34652 21490
rect 33704 20806 33732 21422
rect 34440 21406 34652 21434
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 33784 21344 33836 21350
rect 33782 21312 33784 21321
rect 33876 21344 33928 21350
rect 33836 21312 33838 21321
rect 33876 21286 33928 21292
rect 33782 21247 33838 21256
rect 33888 20942 33916 21286
rect 33876 20936 33928 20942
rect 33876 20878 33928 20884
rect 34336 20868 34388 20874
rect 34336 20810 34388 20816
rect 33692 20800 33744 20806
rect 33692 20742 33744 20748
rect 33600 18964 33652 18970
rect 33600 18906 33652 18912
rect 33612 18426 33640 18906
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 33508 17672 33560 17678
rect 33560 17632 33640 17660
rect 33508 17614 33560 17620
rect 33508 17536 33560 17542
rect 33508 17478 33560 17484
rect 33520 17134 33548 17478
rect 33612 17202 33640 17632
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33508 17128 33560 17134
rect 33508 17070 33560 17076
rect 33520 16726 33548 17070
rect 33508 16720 33560 16726
rect 33508 16662 33560 16668
rect 33416 12980 33468 12986
rect 33416 12922 33468 12928
rect 33140 12776 33192 12782
rect 33140 12718 33192 12724
rect 33508 12776 33560 12782
rect 33508 12718 33560 12724
rect 33600 12776 33652 12782
rect 33600 12718 33652 12724
rect 32956 12436 33008 12442
rect 32956 12378 33008 12384
rect 33324 12300 33376 12306
rect 33324 12242 33376 12248
rect 32956 12232 33008 12238
rect 32954 12200 32956 12209
rect 33008 12200 33010 12209
rect 32954 12135 33010 12144
rect 33336 12102 33364 12242
rect 32864 12096 32916 12102
rect 32864 12038 32916 12044
rect 33048 12096 33100 12102
rect 33048 12038 33100 12044
rect 33232 12096 33284 12102
rect 33232 12038 33284 12044
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 33060 11676 33088 12038
rect 33244 11830 33272 12038
rect 33232 11824 33284 11830
rect 33232 11766 33284 11772
rect 33416 11824 33468 11830
rect 33416 11766 33468 11772
rect 33428 11676 33456 11766
rect 33060 11648 33456 11676
rect 32772 11348 32824 11354
rect 32772 11290 32824 11296
rect 32784 11082 32812 11290
rect 33060 11286 33088 11648
rect 33048 11280 33100 11286
rect 33048 11222 33100 11228
rect 32772 11076 32824 11082
rect 32772 11018 32824 11024
rect 32496 10804 32548 10810
rect 32496 10746 32548 10752
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32784 10606 32812 11018
rect 32772 10600 32824 10606
rect 32772 10542 32824 10548
rect 32680 10192 32732 10198
rect 32680 10134 32732 10140
rect 32588 9920 32640 9926
rect 32588 9862 32640 9868
rect 32404 9648 32456 9654
rect 32404 9590 32456 9596
rect 32220 9172 32272 9178
rect 32220 9114 32272 9120
rect 32232 7954 32260 9114
rect 32600 8838 32628 9862
rect 32692 9450 32720 10134
rect 33060 9994 33088 11222
rect 33520 11218 33548 12718
rect 33508 11212 33560 11218
rect 33508 11154 33560 11160
rect 33612 11098 33640 12718
rect 33704 12434 33732 20742
rect 33876 20256 33928 20262
rect 33876 20198 33928 20204
rect 33968 20256 34020 20262
rect 33968 20198 34020 20204
rect 34152 20256 34204 20262
rect 34152 20198 34204 20204
rect 33888 19922 33916 20198
rect 33876 19916 33928 19922
rect 33876 19858 33928 19864
rect 33980 19446 34008 20198
rect 33968 19440 34020 19446
rect 33968 19382 34020 19388
rect 33784 17604 33836 17610
rect 33784 17546 33836 17552
rect 33796 17202 33824 17546
rect 33784 17196 33836 17202
rect 33784 17138 33836 17144
rect 34060 16992 34112 16998
rect 34060 16934 34112 16940
rect 34072 16590 34100 16934
rect 34060 16584 34112 16590
rect 34060 16526 34112 16532
rect 33784 16448 33836 16454
rect 33784 16390 33836 16396
rect 34060 16448 34112 16454
rect 34060 16390 34112 16396
rect 33796 16182 33824 16390
rect 33784 16176 33836 16182
rect 33784 16118 33836 16124
rect 33876 16040 33928 16046
rect 34072 15994 34100 16390
rect 33928 15988 34100 15994
rect 33876 15982 34100 15988
rect 33888 15966 34100 15982
rect 33876 14952 33928 14958
rect 33876 14894 33928 14900
rect 33888 14278 33916 14894
rect 34072 14822 34100 15966
rect 34060 14816 34112 14822
rect 34060 14758 34112 14764
rect 33876 14272 33928 14278
rect 33876 14214 33928 14220
rect 33968 13864 34020 13870
rect 33968 13806 34020 13812
rect 33980 13462 34008 13806
rect 33968 13456 34020 13462
rect 33968 13398 34020 13404
rect 33704 12406 34008 12434
rect 33690 12336 33746 12345
rect 33980 12306 34008 12406
rect 33690 12271 33692 12280
rect 33744 12271 33746 12280
rect 33876 12300 33928 12306
rect 33692 12242 33744 12248
rect 33876 12242 33928 12248
rect 33968 12300 34020 12306
rect 33968 12242 34020 12248
rect 33520 11070 33640 11098
rect 33888 11082 33916 12242
rect 34164 12102 34192 20198
rect 34348 19310 34376 20810
rect 34440 20466 34468 21406
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35636 20806 35664 21422
rect 35992 21344 36044 21350
rect 35992 21286 36044 21292
rect 36004 20942 36032 21286
rect 35992 20936 36044 20942
rect 35992 20878 36044 20884
rect 34612 20800 34664 20806
rect 34612 20742 34664 20748
rect 35624 20800 35676 20806
rect 35624 20742 35676 20748
rect 34428 20460 34480 20466
rect 34428 20402 34480 20408
rect 34440 19854 34468 20402
rect 34428 19848 34480 19854
rect 34428 19790 34480 19796
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34440 19446 34468 19654
rect 34428 19440 34480 19446
rect 34428 19382 34480 19388
rect 34336 19304 34388 19310
rect 34336 19246 34388 19252
rect 34520 18284 34572 18290
rect 34520 18226 34572 18232
rect 34532 17678 34560 18226
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 34440 16046 34468 17206
rect 34532 17202 34560 17478
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34520 17060 34572 17066
rect 34520 17002 34572 17008
rect 34428 16040 34480 16046
rect 34428 15982 34480 15988
rect 34428 15088 34480 15094
rect 34428 15030 34480 15036
rect 34336 14408 34388 14414
rect 34336 14350 34388 14356
rect 34348 13802 34376 14350
rect 34440 14346 34468 15030
rect 34532 15026 34560 17002
rect 34624 16130 34652 20742
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 34796 20528 34848 20534
rect 34796 20470 34848 20476
rect 34704 19848 34756 19854
rect 34704 19790 34756 19796
rect 34716 19514 34744 19790
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34716 19310 34744 19450
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34716 18834 34744 19246
rect 34704 18828 34756 18834
rect 34704 18770 34756 18776
rect 34808 18154 34836 20470
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20058 35388 20402
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35348 19304 35400 19310
rect 35348 19246 35400 19252
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18426 35388 19246
rect 36096 18630 36124 24074
rect 36188 23662 36216 24686
rect 36464 24342 36492 24686
rect 36636 24676 36688 24682
rect 36636 24618 36688 24624
rect 36452 24336 36504 24342
rect 36452 24278 36504 24284
rect 36176 23656 36228 23662
rect 36176 23598 36228 23604
rect 36464 23225 36492 24278
rect 36544 23520 36596 23526
rect 36544 23462 36596 23468
rect 36450 23216 36506 23225
rect 36450 23151 36506 23160
rect 36268 22976 36320 22982
rect 36188 22936 36268 22964
rect 36188 22778 36216 22936
rect 36268 22918 36320 22924
rect 36176 22772 36228 22778
rect 36176 22714 36228 22720
rect 36268 22704 36320 22710
rect 36268 22646 36320 22652
rect 36280 22098 36308 22646
rect 36464 22574 36492 23151
rect 36556 23117 36584 23462
rect 36544 23111 36596 23117
rect 36544 23053 36596 23059
rect 36452 22568 36504 22574
rect 36452 22510 36504 22516
rect 36648 22420 36676 24618
rect 36740 24596 36768 26318
rect 36740 24568 36860 24596
rect 36728 24064 36780 24070
rect 36728 24006 36780 24012
rect 36372 22392 36676 22420
rect 36268 22092 36320 22098
rect 36268 22034 36320 22040
rect 36176 20256 36228 20262
rect 36176 20198 36228 20204
rect 36188 19922 36216 20198
rect 36176 19916 36228 19922
rect 36176 19858 36228 19864
rect 36372 19514 36400 22392
rect 36740 22250 36768 24006
rect 36832 22982 36860 24568
rect 36924 23032 36952 28970
rect 37016 26761 37044 34410
rect 37292 34066 37320 34478
rect 37280 34060 37332 34066
rect 37280 34002 37332 34008
rect 37568 33930 37596 34886
rect 37660 34678 37688 35430
rect 37648 34672 37700 34678
rect 37648 34614 37700 34620
rect 37556 33924 37608 33930
rect 37556 33866 37608 33872
rect 37188 32904 37240 32910
rect 37240 32852 37320 32858
rect 37188 32846 37320 32852
rect 37200 32830 37320 32846
rect 37292 32366 37320 32830
rect 37372 32428 37424 32434
rect 37372 32370 37424 32376
rect 37280 32360 37332 32366
rect 37280 32302 37332 32308
rect 37384 32026 37412 32370
rect 37372 32020 37424 32026
rect 37372 31962 37424 31968
rect 37740 30728 37792 30734
rect 37740 30670 37792 30676
rect 37556 30388 37608 30394
rect 37556 30330 37608 30336
rect 37568 30258 37596 30330
rect 37372 30252 37424 30258
rect 37372 30194 37424 30200
rect 37556 30252 37608 30258
rect 37556 30194 37608 30200
rect 37096 29640 37148 29646
rect 37096 29582 37148 29588
rect 37108 29209 37136 29582
rect 37384 29578 37412 30194
rect 37372 29572 37424 29578
rect 37372 29514 37424 29520
rect 37094 29200 37150 29209
rect 37094 29135 37150 29144
rect 37646 28656 37702 28665
rect 37646 28591 37702 28600
rect 37660 28558 37688 28591
rect 37648 28552 37700 28558
rect 37648 28494 37700 28500
rect 37752 28218 37780 30670
rect 37844 30546 37872 36774
rect 37924 36780 37976 36786
rect 37924 36722 37976 36728
rect 38108 36780 38160 36786
rect 38108 36722 38160 36728
rect 37936 36378 37964 36722
rect 37924 36372 37976 36378
rect 37924 36314 37976 36320
rect 38016 36168 38068 36174
rect 38120 36156 38148 36722
rect 38068 36128 38148 36156
rect 38016 36110 38068 36116
rect 38108 35624 38160 35630
rect 38108 35566 38160 35572
rect 38120 33658 38148 35566
rect 38304 34746 38332 40054
rect 38568 39568 38620 39574
rect 38568 39510 38620 39516
rect 38580 39030 38608 39510
rect 38568 39024 38620 39030
rect 38568 38966 38620 38972
rect 38384 38956 38436 38962
rect 38384 38898 38436 38904
rect 38396 38486 38424 38898
rect 38384 38480 38436 38486
rect 38384 38422 38436 38428
rect 38660 38344 38712 38350
rect 38660 38286 38712 38292
rect 38568 37800 38620 37806
rect 38568 37742 38620 37748
rect 38580 36582 38608 37742
rect 38672 37738 38700 38286
rect 38660 37732 38712 37738
rect 38660 37674 38712 37680
rect 38672 36922 38700 37674
rect 38660 36916 38712 36922
rect 38660 36858 38712 36864
rect 38568 36576 38620 36582
rect 38568 36518 38620 36524
rect 38658 36272 38714 36281
rect 38658 36207 38714 36216
rect 38672 36174 38700 36207
rect 38660 36168 38712 36174
rect 38660 36110 38712 36116
rect 38476 36100 38528 36106
rect 38476 36042 38528 36048
rect 38568 36100 38620 36106
rect 38568 36042 38620 36048
rect 38488 35630 38516 36042
rect 38580 35986 38608 36042
rect 38752 36032 38804 36038
rect 38580 35958 38700 35986
rect 38752 35974 38804 35980
rect 38672 35766 38700 35958
rect 38660 35760 38712 35766
rect 38660 35702 38712 35708
rect 38476 35624 38528 35630
rect 38476 35566 38528 35572
rect 38764 35562 38792 35974
rect 38752 35556 38804 35562
rect 38752 35498 38804 35504
rect 38660 35284 38712 35290
rect 38660 35226 38712 35232
rect 38292 34740 38344 34746
rect 38292 34682 38344 34688
rect 38672 34610 38700 35226
rect 38660 34604 38712 34610
rect 38660 34546 38712 34552
rect 38672 33998 38700 34546
rect 38660 33992 38712 33998
rect 38660 33934 38712 33940
rect 38108 33652 38160 33658
rect 38108 33594 38160 33600
rect 38292 33516 38344 33522
rect 38292 33458 38344 33464
rect 38660 33516 38712 33522
rect 38660 33458 38712 33464
rect 38304 33114 38332 33458
rect 38292 33108 38344 33114
rect 38292 33050 38344 33056
rect 38108 32836 38160 32842
rect 38108 32778 38160 32784
rect 37924 32224 37976 32230
rect 37924 32166 37976 32172
rect 37936 31414 37964 32166
rect 38120 32026 38148 32778
rect 38568 32768 38620 32774
rect 38568 32710 38620 32716
rect 38108 32020 38160 32026
rect 38108 31962 38160 31968
rect 38580 31890 38608 32710
rect 38672 32570 38700 33458
rect 38660 32564 38712 32570
rect 38660 32506 38712 32512
rect 38752 32224 38804 32230
rect 38752 32166 38804 32172
rect 38764 31958 38792 32166
rect 38752 31952 38804 31958
rect 38752 31894 38804 31900
rect 38568 31884 38620 31890
rect 38568 31826 38620 31832
rect 38476 31680 38528 31686
rect 38476 31622 38528 31628
rect 38660 31680 38712 31686
rect 38660 31622 38712 31628
rect 37924 31408 37976 31414
rect 37924 31350 37976 31356
rect 37936 30734 37964 31350
rect 37924 30728 37976 30734
rect 37924 30670 37976 30676
rect 38200 30660 38252 30666
rect 38200 30602 38252 30608
rect 38292 30660 38344 30666
rect 38292 30602 38344 30608
rect 37844 30518 37964 30546
rect 37936 30326 37964 30518
rect 38212 30394 38240 30602
rect 38200 30388 38252 30394
rect 38200 30330 38252 30336
rect 37924 30320 37976 30326
rect 37924 30262 37976 30268
rect 37832 30252 37884 30258
rect 37832 30194 37884 30200
rect 37844 29646 37872 30194
rect 38016 29708 38068 29714
rect 38016 29650 38068 29656
rect 37832 29640 37884 29646
rect 37832 29582 37884 29588
rect 37924 29096 37976 29102
rect 37924 29038 37976 29044
rect 37936 28626 37964 29038
rect 37924 28620 37976 28626
rect 37924 28562 37976 28568
rect 37832 28484 37884 28490
rect 37832 28426 37884 28432
rect 37844 28218 37872 28426
rect 37740 28212 37792 28218
rect 37740 28154 37792 28160
rect 37832 28212 37884 28218
rect 37832 28154 37884 28160
rect 37372 28144 37424 28150
rect 37372 28086 37424 28092
rect 37280 27600 37332 27606
rect 37278 27568 37280 27577
rect 37332 27568 37334 27577
rect 37278 27503 37334 27512
rect 37002 26752 37058 26761
rect 37002 26687 37058 26696
rect 37016 26382 37044 26687
rect 37096 26512 37148 26518
rect 37096 26454 37148 26460
rect 37004 26376 37056 26382
rect 37004 26318 37056 26324
rect 37004 24880 37056 24886
rect 37004 24822 37056 24828
rect 37016 24274 37044 24822
rect 37004 24268 37056 24274
rect 37004 24210 37056 24216
rect 37016 23730 37044 24210
rect 37004 23724 37056 23730
rect 37004 23666 37056 23672
rect 37108 23050 37136 26454
rect 37186 26344 37242 26353
rect 37186 26279 37188 26288
rect 37240 26279 37242 26288
rect 37188 26250 37240 26256
rect 37280 25832 37332 25838
rect 37280 25774 37332 25780
rect 37292 25430 37320 25774
rect 37280 25424 37332 25430
rect 37280 25366 37332 25372
rect 37292 24886 37320 25366
rect 37280 24880 37332 24886
rect 37280 24822 37332 24828
rect 37280 24608 37332 24614
rect 37280 24550 37332 24556
rect 37292 24274 37320 24550
rect 37280 24268 37332 24274
rect 37280 24210 37332 24216
rect 37004 23044 37056 23050
rect 36924 23004 37004 23032
rect 37004 22986 37056 22992
rect 37096 23044 37148 23050
rect 37096 22986 37148 22992
rect 36820 22976 36872 22982
rect 36820 22918 36872 22924
rect 36648 22222 36768 22250
rect 36544 22092 36596 22098
rect 36544 22034 36596 22040
rect 36452 21684 36504 21690
rect 36452 21626 36504 21632
rect 36464 19768 36492 21626
rect 36556 20942 36584 22034
rect 36544 20936 36596 20942
rect 36544 20878 36596 20884
rect 36648 19854 36676 22222
rect 36728 21344 36780 21350
rect 36728 21286 36780 21292
rect 36636 19848 36688 19854
rect 36636 19790 36688 19796
rect 36544 19780 36596 19786
rect 36464 19740 36544 19768
rect 36544 19722 36596 19728
rect 36360 19508 36412 19514
rect 36360 19450 36412 19456
rect 35440 18624 35492 18630
rect 35440 18566 35492 18572
rect 36084 18624 36136 18630
rect 36084 18566 36136 18572
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 34796 18148 34848 18154
rect 34796 18090 34848 18096
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35452 17882 35480 18566
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35992 18148 36044 18154
rect 35992 18090 36044 18096
rect 35532 18080 35584 18086
rect 35532 18022 35584 18028
rect 35440 17876 35492 17882
rect 35440 17818 35492 17824
rect 35072 17808 35124 17814
rect 35072 17750 35124 17756
rect 34796 17672 34848 17678
rect 34796 17614 34848 17620
rect 34980 17672 35032 17678
rect 34980 17614 35032 17620
rect 34704 17604 34756 17610
rect 34704 17546 34756 17552
rect 34716 16454 34744 17546
rect 34808 17202 34836 17614
rect 34992 17202 35020 17614
rect 34796 17196 34848 17202
rect 34796 17138 34848 17144
rect 34980 17196 35032 17202
rect 34980 17138 35032 17144
rect 34808 16794 34836 17138
rect 35084 17134 35112 17750
rect 35544 17610 35572 18022
rect 35532 17604 35584 17610
rect 35532 17546 35584 17552
rect 35440 17536 35492 17542
rect 35440 17478 35492 17484
rect 35072 17128 35124 17134
rect 35072 17070 35124 17076
rect 35256 17128 35308 17134
rect 35256 17070 35308 17076
rect 35268 16946 35296 17070
rect 35268 16918 35388 16946
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 34888 16788 34940 16794
rect 34888 16730 34940 16736
rect 34808 16522 34836 16730
rect 34900 16658 34928 16730
rect 34888 16652 34940 16658
rect 34888 16594 34940 16600
rect 34980 16584 35032 16590
rect 34980 16526 35032 16532
rect 35256 16584 35308 16590
rect 35256 16526 35308 16532
rect 34796 16516 34848 16522
rect 34796 16458 34848 16464
rect 34704 16448 34756 16454
rect 34704 16390 34756 16396
rect 34716 16250 34744 16390
rect 34704 16244 34756 16250
rect 34704 16186 34756 16192
rect 34624 16102 34744 16130
rect 34520 15020 34572 15026
rect 34520 14962 34572 14968
rect 34428 14340 34480 14346
rect 34428 14282 34480 14288
rect 34336 13796 34388 13802
rect 34336 13738 34388 13744
rect 34440 12918 34468 14282
rect 34612 14272 34664 14278
rect 34612 14214 34664 14220
rect 34624 13870 34652 14214
rect 34612 13864 34664 13870
rect 34612 13806 34664 13812
rect 34428 12912 34480 12918
rect 34428 12854 34480 12860
rect 34520 12776 34572 12782
rect 34520 12718 34572 12724
rect 34152 12096 34204 12102
rect 34152 12038 34204 12044
rect 34164 11354 34192 12038
rect 34532 11626 34560 12718
rect 34612 12640 34664 12646
rect 34612 12582 34664 12588
rect 34624 12306 34652 12582
rect 34716 12442 34744 16102
rect 34992 15978 35020 16526
rect 35164 16516 35216 16522
rect 35164 16458 35216 16464
rect 35176 16046 35204 16458
rect 35268 16250 35296 16526
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 35256 16108 35308 16114
rect 35256 16050 35308 16056
rect 35164 16040 35216 16046
rect 35164 15982 35216 15988
rect 34980 15972 35032 15978
rect 34980 15914 35032 15920
rect 35268 15910 35296 16050
rect 35256 15904 35308 15910
rect 35256 15846 35308 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35256 15564 35308 15570
rect 35360 15552 35388 16918
rect 35452 16522 35480 17478
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35716 16992 35768 16998
rect 35716 16934 35768 16940
rect 35728 16590 35756 16934
rect 35716 16584 35768 16590
rect 35716 16526 35768 16532
rect 35440 16516 35492 16522
rect 35440 16458 35492 16464
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35308 15524 35388 15552
rect 35256 15506 35308 15512
rect 35440 15428 35492 15434
rect 35440 15370 35492 15376
rect 35452 15162 35480 15370
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35440 15156 35492 15162
rect 35440 15098 35492 15104
rect 35440 14952 35492 14958
rect 35440 14894 35492 14900
rect 35348 14884 35400 14890
rect 35348 14826 35400 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35164 14408 35216 14414
rect 35164 14350 35216 14356
rect 35176 14074 35204 14350
rect 35360 14278 35388 14826
rect 35452 14550 35480 14894
rect 35440 14544 35492 14550
rect 35440 14486 35492 14492
rect 35348 14272 35400 14278
rect 35348 14214 35400 14220
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 35164 14068 35216 14074
rect 35164 14010 35216 14016
rect 34808 13410 34836 14010
rect 35348 13932 35400 13938
rect 35348 13874 35400 13880
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34808 13382 34928 13410
rect 34900 13326 34928 13382
rect 34888 13320 34940 13326
rect 34888 13262 34940 13268
rect 35072 13320 35124 13326
rect 35072 13262 35124 13268
rect 35084 13190 35112 13262
rect 35072 13184 35124 13190
rect 35072 13126 35124 13132
rect 35360 12986 35388 13874
rect 35440 13796 35492 13802
rect 35440 13738 35492 13744
rect 35452 13394 35480 13738
rect 35440 13388 35492 13394
rect 35440 13330 35492 13336
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34612 12300 34664 12306
rect 34612 12242 34664 12248
rect 35348 12164 35400 12170
rect 35348 12106 35400 12112
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 34808 11830 34836 12038
rect 35360 11830 35388 12106
rect 34796 11824 34848 11830
rect 34796 11766 34848 11772
rect 35348 11824 35400 11830
rect 35348 11766 35400 11772
rect 34520 11620 34572 11626
rect 34520 11562 34572 11568
rect 34152 11348 34204 11354
rect 34152 11290 34204 11296
rect 34532 11150 34560 11562
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34612 11348 34664 11354
rect 34612 11290 34664 11296
rect 34520 11144 34572 11150
rect 34520 11086 34572 11092
rect 33876 11076 33928 11082
rect 33520 10742 33548 11070
rect 33876 11018 33928 11024
rect 33508 10736 33560 10742
rect 33508 10678 33560 10684
rect 33140 10600 33192 10606
rect 33140 10542 33192 10548
rect 33152 10266 33180 10542
rect 33140 10260 33192 10266
rect 33192 10220 33272 10248
rect 33140 10202 33192 10208
rect 33140 10124 33192 10130
rect 33140 10066 33192 10072
rect 33048 9988 33100 9994
rect 33048 9930 33100 9936
rect 33152 9602 33180 10066
rect 33244 9994 33272 10220
rect 33520 10062 33548 10678
rect 34520 10600 34572 10606
rect 34520 10542 34572 10548
rect 34336 10464 34388 10470
rect 34336 10406 34388 10412
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33232 9988 33284 9994
rect 33232 9930 33284 9936
rect 32968 9574 33180 9602
rect 32680 9444 32732 9450
rect 32680 9386 32732 9392
rect 32588 8832 32640 8838
rect 32588 8774 32640 8780
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 32416 8090 32444 8366
rect 32404 8084 32456 8090
rect 32404 8026 32456 8032
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32128 7880 32180 7886
rect 32128 7822 32180 7828
rect 32140 7750 32168 7822
rect 32128 7744 32180 7750
rect 32128 7686 32180 7692
rect 32692 7546 32720 9386
rect 32968 9042 32996 9574
rect 33048 9512 33100 9518
rect 33048 9454 33100 9460
rect 32956 9036 33008 9042
rect 32956 8978 33008 8984
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 32876 8294 32904 8910
rect 33060 8634 33088 9454
rect 33244 9110 33272 9930
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 33888 9654 33916 9862
rect 33876 9648 33928 9654
rect 33876 9590 33928 9596
rect 33324 9376 33376 9382
rect 33324 9318 33376 9324
rect 33336 9110 33364 9318
rect 34348 9178 34376 10406
rect 34532 10266 34560 10542
rect 34520 10260 34572 10266
rect 34520 10202 34572 10208
rect 34624 10130 34652 11290
rect 35360 11286 35388 11766
rect 35452 11286 35480 13330
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 35532 12980 35584 12986
rect 35532 12922 35584 12928
rect 35544 12170 35572 12922
rect 35716 12844 35768 12850
rect 35716 12786 35768 12792
rect 35728 12209 35756 12786
rect 35900 12640 35952 12646
rect 35900 12582 35952 12588
rect 35912 12306 35940 12582
rect 36004 12374 36032 18090
rect 36096 17610 36124 18566
rect 36372 18426 36400 19450
rect 36544 19304 36596 19310
rect 36544 19246 36596 19252
rect 36556 18970 36584 19246
rect 36544 18964 36596 18970
rect 36544 18906 36596 18912
rect 36556 18698 36584 18906
rect 36544 18692 36596 18698
rect 36544 18634 36596 18640
rect 36360 18420 36412 18426
rect 36360 18362 36412 18368
rect 36452 18216 36504 18222
rect 36452 18158 36504 18164
rect 36360 18080 36412 18086
rect 36360 18022 36412 18028
rect 36084 17604 36136 17610
rect 36084 17546 36136 17552
rect 36372 16590 36400 18022
rect 36464 17746 36492 18158
rect 36452 17740 36504 17746
rect 36452 17682 36504 17688
rect 36360 16584 36412 16590
rect 36360 16526 36412 16532
rect 36372 16114 36400 16526
rect 36360 16108 36412 16114
rect 36360 16050 36412 16056
rect 36464 14940 36492 17682
rect 36556 17270 36584 18634
rect 36544 17264 36596 17270
rect 36544 17206 36596 17212
rect 36556 15910 36584 17206
rect 36544 15904 36596 15910
rect 36544 15846 36596 15852
rect 36556 15366 36584 15846
rect 36544 15360 36596 15366
rect 36544 15302 36596 15308
rect 36544 14952 36596 14958
rect 36464 14912 36544 14940
rect 36544 14894 36596 14900
rect 36452 14816 36504 14822
rect 36452 14758 36504 14764
rect 36464 14006 36492 14758
rect 36452 14000 36504 14006
rect 36452 13942 36504 13948
rect 36084 13252 36136 13258
rect 36084 13194 36136 13200
rect 36268 13252 36320 13258
rect 36268 13194 36320 13200
rect 36096 12986 36124 13194
rect 36084 12980 36136 12986
rect 36084 12922 36136 12928
rect 35992 12368 36044 12374
rect 35992 12310 36044 12316
rect 35900 12300 35952 12306
rect 35900 12242 35952 12248
rect 35714 12200 35770 12209
rect 35532 12164 35584 12170
rect 35714 12135 35770 12144
rect 35532 12106 35584 12112
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 36176 11892 36228 11898
rect 36176 11834 36228 11840
rect 36084 11620 36136 11626
rect 36084 11562 36136 11568
rect 35532 11552 35584 11558
rect 35532 11494 35584 11500
rect 35544 11354 35572 11494
rect 35532 11348 35584 11354
rect 35532 11290 35584 11296
rect 35348 11280 35400 11286
rect 35348 11222 35400 11228
rect 35440 11280 35492 11286
rect 35440 11222 35492 11228
rect 36096 11218 36124 11562
rect 35256 11212 35308 11218
rect 35256 11154 35308 11160
rect 36084 11212 36136 11218
rect 36084 11154 36136 11160
rect 35164 11076 35216 11082
rect 35164 11018 35216 11024
rect 35176 10690 35204 11018
rect 35268 10810 35296 11154
rect 35348 11144 35400 11150
rect 35348 11086 35400 11092
rect 35440 11144 35492 11150
rect 35440 11086 35492 11092
rect 35256 10804 35308 10810
rect 35256 10746 35308 10752
rect 34796 10668 34848 10674
rect 35176 10662 35296 10690
rect 34796 10610 34848 10616
rect 34612 10124 34664 10130
rect 34612 10066 34664 10072
rect 34808 9722 34836 10610
rect 35268 10418 35296 10662
rect 35360 10606 35388 11086
rect 35452 10690 35480 11086
rect 36188 10962 36216 11834
rect 36096 10934 36216 10962
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 35452 10674 35572 10690
rect 36096 10674 36124 10934
rect 35452 10668 35584 10674
rect 35452 10662 35532 10668
rect 35532 10610 35584 10616
rect 36084 10668 36136 10674
rect 36084 10610 36136 10616
rect 35348 10600 35400 10606
rect 35348 10542 35400 10548
rect 35544 10538 35572 10610
rect 35532 10532 35584 10538
rect 35532 10474 35584 10480
rect 35268 10390 35388 10418
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 10130 35388 10390
rect 36096 10146 36124 10610
rect 36176 10600 36228 10606
rect 36176 10542 36228 10548
rect 35348 10124 35400 10130
rect 35348 10066 35400 10072
rect 35440 10124 35492 10130
rect 35440 10066 35492 10072
rect 36004 10118 36124 10146
rect 34796 9716 34848 9722
rect 34796 9658 34848 9664
rect 35452 9602 35480 10066
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 36004 9654 36032 10118
rect 36084 10056 36136 10062
rect 36084 9998 36136 10004
rect 35992 9648 36044 9654
rect 35452 9586 35572 9602
rect 35992 9590 36044 9596
rect 35452 9580 35584 9586
rect 35452 9574 35532 9580
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34336 9172 34388 9178
rect 34336 9114 34388 9120
rect 33232 9104 33284 9110
rect 33232 9046 33284 9052
rect 33324 9104 33376 9110
rect 33324 9046 33376 9052
rect 33232 8968 33284 8974
rect 33232 8910 33284 8916
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 33060 8430 33088 8570
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 32864 8288 32916 8294
rect 32864 8230 32916 8236
rect 32876 7886 32904 8230
rect 33244 8090 33272 8910
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 34256 8566 34284 8774
rect 34244 8560 34296 8566
rect 34244 8502 34296 8508
rect 34336 8424 34388 8430
rect 34336 8366 34388 8372
rect 33876 8288 33928 8294
rect 33876 8230 33928 8236
rect 33232 8084 33284 8090
rect 33232 8026 33284 8032
rect 33888 7954 33916 8230
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 32864 7880 32916 7886
rect 32864 7822 32916 7828
rect 32772 7812 32824 7818
rect 32772 7754 32824 7760
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32680 7540 32732 7546
rect 32680 7482 32732 7488
rect 31852 6452 31904 6458
rect 31852 6394 31904 6400
rect 31864 6322 31892 6394
rect 32416 6322 32444 7482
rect 32784 7426 32812 7754
rect 32600 7398 32812 7426
rect 34152 7404 34204 7410
rect 32600 6361 32628 7398
rect 34152 7346 34204 7352
rect 32772 6996 32824 7002
rect 32772 6938 32824 6944
rect 32680 6384 32732 6390
rect 32586 6352 32642 6361
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31668 6316 31720 6322
rect 31668 6258 31720 6264
rect 31852 6316 31904 6322
rect 31852 6258 31904 6264
rect 31944 6316 31996 6322
rect 31944 6258 31996 6264
rect 32404 6316 32456 6322
rect 32680 6326 32732 6332
rect 32586 6287 32588 6296
rect 32404 6258 32456 6264
rect 32640 6287 32642 6296
rect 32588 6258 32640 6264
rect 31312 5914 31340 6258
rect 31484 6180 31536 6186
rect 31484 6122 31536 6128
rect 31300 5908 31352 5914
rect 31300 5850 31352 5856
rect 31208 5704 31260 5710
rect 31208 5646 31260 5652
rect 30748 5568 30800 5574
rect 30748 5510 30800 5516
rect 30840 5568 30892 5574
rect 30840 5510 30892 5516
rect 30656 5296 30708 5302
rect 30656 5238 30708 5244
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 28448 5160 28500 5166
rect 28448 5102 28500 5108
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 31220 4690 31248 5646
rect 31496 4690 31524 6122
rect 31680 5574 31708 6258
rect 31668 5568 31720 5574
rect 31668 5510 31720 5516
rect 31956 5370 31984 6258
rect 32128 6112 32180 6118
rect 32128 6054 32180 6060
rect 32140 5778 32168 6054
rect 32692 5914 32720 6326
rect 32680 5908 32732 5914
rect 32680 5850 32732 5856
rect 32128 5772 32180 5778
rect 32128 5714 32180 5720
rect 31944 5364 31996 5370
rect 31944 5306 31996 5312
rect 32784 5166 32812 6938
rect 33048 6452 33100 6458
rect 33048 6394 33100 6400
rect 33060 5642 33088 6394
rect 33232 6112 33284 6118
rect 33232 6054 33284 6060
rect 33244 5710 33272 6054
rect 34164 5710 34192 7346
rect 34348 7342 34376 8366
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35348 7948 35400 7954
rect 35348 7890 35400 7896
rect 35164 7812 35216 7818
rect 35164 7754 35216 7760
rect 34888 7744 34940 7750
rect 34888 7686 34940 7692
rect 34704 7540 34756 7546
rect 34704 7482 34756 7488
rect 34336 7336 34388 7342
rect 34336 7278 34388 7284
rect 34348 7206 34376 7278
rect 34336 7200 34388 7206
rect 34336 7142 34388 7148
rect 34716 7002 34744 7482
rect 34796 7472 34848 7478
rect 34796 7414 34848 7420
rect 34704 6996 34756 7002
rect 34704 6938 34756 6944
rect 34612 6792 34664 6798
rect 34612 6734 34664 6740
rect 34336 6724 34388 6730
rect 34336 6666 34388 6672
rect 34348 6458 34376 6666
rect 34336 6452 34388 6458
rect 34336 6394 34388 6400
rect 33232 5704 33284 5710
rect 33232 5646 33284 5652
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 33048 5636 33100 5642
rect 33048 5578 33100 5584
rect 32772 5160 32824 5166
rect 32772 5102 32824 5108
rect 32956 5160 33008 5166
rect 32956 5102 33008 5108
rect 32968 4826 32996 5102
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 31208 4684 31260 4690
rect 31208 4626 31260 4632
rect 31484 4684 31536 4690
rect 31484 4626 31536 4632
rect 33060 4554 33088 5578
rect 34624 5574 34652 6734
rect 34808 6662 34836 7414
rect 34900 7410 34928 7686
rect 34980 7540 35032 7546
rect 34980 7482 35032 7488
rect 34992 7410 35020 7482
rect 35176 7410 35204 7754
rect 34888 7404 34940 7410
rect 34888 7346 34940 7352
rect 34980 7404 35032 7410
rect 34980 7346 35032 7352
rect 35164 7404 35216 7410
rect 35164 7346 35216 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6656 34848 6662
rect 34796 6598 34848 6604
rect 34704 6248 34756 6254
rect 34704 6190 34756 6196
rect 34612 5568 34664 5574
rect 34612 5510 34664 5516
rect 34624 5302 34652 5510
rect 34716 5370 34744 6190
rect 34704 5364 34756 5370
rect 34704 5306 34756 5312
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 34808 5234 34836 6598
rect 35360 6390 35388 7890
rect 35452 7546 35480 9574
rect 35532 9522 35584 9528
rect 36096 9518 36124 9998
rect 36084 9512 36136 9518
rect 36084 9454 36136 9460
rect 36188 9450 36216 10542
rect 36176 9444 36228 9450
rect 36176 9386 36228 9392
rect 36280 9382 36308 13194
rect 36556 12782 36584 14894
rect 36544 12776 36596 12782
rect 36544 12718 36596 12724
rect 36740 12434 36768 21286
rect 36832 13462 36860 22918
rect 36912 22432 36964 22438
rect 36912 22374 36964 22380
rect 36924 22234 36952 22374
rect 36912 22228 36964 22234
rect 36912 22170 36964 22176
rect 37016 22094 37044 22986
rect 37384 22794 37412 28086
rect 38028 28082 38056 29650
rect 38016 28076 38068 28082
rect 38016 28018 38068 28024
rect 37556 28008 37608 28014
rect 37556 27950 37608 27956
rect 37568 26858 37596 27950
rect 38200 27872 38252 27878
rect 38200 27814 38252 27820
rect 37740 27668 37792 27674
rect 37740 27610 37792 27616
rect 37752 27130 37780 27610
rect 37740 27124 37792 27130
rect 37740 27066 37792 27072
rect 37556 26852 37608 26858
rect 37556 26794 37608 26800
rect 37556 26240 37608 26246
rect 37556 26182 37608 26188
rect 37568 25974 37596 26182
rect 37556 25968 37608 25974
rect 37556 25910 37608 25916
rect 37556 24064 37608 24070
rect 37556 24006 37608 24012
rect 37568 23798 37596 24006
rect 37556 23792 37608 23798
rect 37556 23734 37608 23740
rect 37740 22976 37792 22982
rect 37740 22918 37792 22924
rect 37200 22778 37412 22794
rect 37188 22772 37412 22778
rect 37240 22766 37412 22772
rect 37188 22714 37240 22720
rect 37752 22642 37780 22918
rect 38212 22778 38240 27814
rect 38304 26382 38332 30602
rect 38384 30252 38436 30258
rect 38384 30194 38436 30200
rect 38396 27606 38424 30194
rect 38488 29714 38516 31622
rect 38672 30326 38700 31622
rect 38856 30938 38884 40054
rect 39224 39982 39252 40462
rect 39316 40186 39344 41006
rect 39592 40186 39620 41074
rect 40132 41064 40184 41070
rect 40132 41006 40184 41012
rect 39856 40996 39908 41002
rect 39856 40938 39908 40944
rect 39304 40180 39356 40186
rect 39304 40122 39356 40128
rect 39580 40180 39632 40186
rect 39580 40122 39632 40128
rect 39212 39976 39264 39982
rect 39212 39918 39264 39924
rect 39224 38894 39252 39918
rect 39592 39386 39620 40122
rect 39868 39982 39896 40938
rect 40040 40724 40092 40730
rect 40040 40666 40092 40672
rect 39856 39976 39908 39982
rect 39856 39918 39908 39924
rect 39396 39364 39448 39370
rect 39396 39306 39448 39312
rect 39500 39358 39620 39386
rect 39672 39432 39724 39438
rect 39672 39374 39724 39380
rect 39212 38888 39264 38894
rect 39212 38830 39264 38836
rect 39224 38418 39252 38830
rect 39212 38412 39264 38418
rect 39212 38354 39264 38360
rect 39408 38350 39436 39306
rect 39396 38344 39448 38350
rect 39396 38286 39448 38292
rect 39028 36780 39080 36786
rect 39028 36722 39080 36728
rect 39040 36378 39068 36722
rect 39028 36372 39080 36378
rect 39028 36314 39080 36320
rect 38936 36304 38988 36310
rect 38936 36246 38988 36252
rect 38948 36174 38976 36246
rect 38936 36168 38988 36174
rect 39304 36168 39356 36174
rect 38936 36110 38988 36116
rect 39210 36136 39266 36145
rect 38948 35698 38976 36110
rect 39304 36110 39356 36116
rect 39210 36071 39212 36080
rect 39264 36071 39266 36080
rect 39212 36042 39264 36048
rect 39316 35834 39344 36110
rect 39304 35828 39356 35834
rect 39304 35770 39356 35776
rect 39212 35760 39264 35766
rect 39212 35702 39264 35708
rect 38936 35692 38988 35698
rect 38936 35634 38988 35640
rect 38948 34542 38976 35634
rect 39028 34944 39080 34950
rect 39028 34886 39080 34892
rect 38936 34536 38988 34542
rect 38936 34478 38988 34484
rect 39040 33658 39068 34886
rect 39224 34610 39252 35702
rect 39120 34604 39172 34610
rect 39120 34546 39172 34552
rect 39212 34604 39264 34610
rect 39212 34546 39264 34552
rect 39028 33652 39080 33658
rect 39028 33594 39080 33600
rect 38936 31816 38988 31822
rect 38936 31758 38988 31764
rect 38844 30932 38896 30938
rect 38844 30874 38896 30880
rect 38660 30320 38712 30326
rect 38660 30262 38712 30268
rect 38752 30320 38804 30326
rect 38752 30262 38804 30268
rect 38660 30184 38712 30190
rect 38660 30126 38712 30132
rect 38672 29850 38700 30126
rect 38660 29844 38712 29850
rect 38660 29786 38712 29792
rect 38476 29708 38528 29714
rect 38476 29650 38528 29656
rect 38568 29504 38620 29510
rect 38568 29446 38620 29452
rect 38474 28520 38530 28529
rect 38474 28455 38530 28464
rect 38488 28082 38516 28455
rect 38476 28076 38528 28082
rect 38476 28018 38528 28024
rect 38384 27600 38436 27606
rect 38384 27542 38436 27548
rect 38396 27062 38424 27542
rect 38580 27062 38608 29446
rect 38660 28076 38712 28082
rect 38660 28018 38712 28024
rect 38672 27538 38700 28018
rect 38660 27532 38712 27538
rect 38660 27474 38712 27480
rect 38384 27056 38436 27062
rect 38384 26998 38436 27004
rect 38568 27056 38620 27062
rect 38568 26998 38620 27004
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38580 25158 38608 26998
rect 38568 25152 38620 25158
rect 38568 25094 38620 25100
rect 38764 24818 38792 30262
rect 38948 30190 38976 31758
rect 39132 30326 39160 34546
rect 39224 34202 39252 34546
rect 39212 34196 39264 34202
rect 39212 34138 39264 34144
rect 39500 31890 39528 39358
rect 39580 39296 39632 39302
rect 39580 39238 39632 39244
rect 39592 38554 39620 39238
rect 39580 38548 39632 38554
rect 39580 38490 39632 38496
rect 39592 38350 39620 38490
rect 39684 38350 39712 39374
rect 39764 39296 39816 39302
rect 39764 39238 39816 39244
rect 39776 39030 39804 39238
rect 39764 39024 39816 39030
rect 39764 38966 39816 38972
rect 39580 38344 39632 38350
rect 39580 38286 39632 38292
rect 39672 38344 39724 38350
rect 39672 38286 39724 38292
rect 39684 38010 39712 38286
rect 39672 38004 39724 38010
rect 39672 37946 39724 37952
rect 39868 37806 39896 39918
rect 40052 38350 40080 40666
rect 40144 40662 40172 41006
rect 40236 40730 40264 41074
rect 40224 40724 40276 40730
rect 40224 40666 40276 40672
rect 40132 40656 40184 40662
rect 40184 40604 40264 40610
rect 40132 40598 40264 40604
rect 40144 40582 40264 40598
rect 40132 40452 40184 40458
rect 40132 40394 40184 40400
rect 40144 39030 40172 40394
rect 40236 39506 40264 40582
rect 40224 39500 40276 39506
rect 40224 39442 40276 39448
rect 40236 39098 40264 39442
rect 40960 39432 41012 39438
rect 40960 39374 41012 39380
rect 42156 39432 42208 39438
rect 42156 39374 42208 39380
rect 40316 39296 40368 39302
rect 40316 39238 40368 39244
rect 40224 39092 40276 39098
rect 40224 39034 40276 39040
rect 40132 39024 40184 39030
rect 40132 38966 40184 38972
rect 40144 38554 40172 38966
rect 40132 38548 40184 38554
rect 40132 38490 40184 38496
rect 40040 38344 40092 38350
rect 40040 38286 40092 38292
rect 40052 37874 40080 38286
rect 40132 38208 40184 38214
rect 40132 38150 40184 38156
rect 40144 37874 40172 38150
rect 40328 38010 40356 39238
rect 40972 39098 41000 39374
rect 41420 39296 41472 39302
rect 41420 39238 41472 39244
rect 41432 39098 41460 39238
rect 40960 39092 41012 39098
rect 40960 39034 41012 39040
rect 41420 39092 41472 39098
rect 41420 39034 41472 39040
rect 41236 39024 41288 39030
rect 41236 38966 41288 38972
rect 41052 38752 41104 38758
rect 41052 38694 41104 38700
rect 41064 38418 41092 38694
rect 41144 38548 41196 38554
rect 41144 38490 41196 38496
rect 41052 38412 41104 38418
rect 41052 38354 41104 38360
rect 41156 38282 41184 38490
rect 41144 38276 41196 38282
rect 41144 38218 41196 38224
rect 40316 38004 40368 38010
rect 40316 37946 40368 37952
rect 40868 37936 40920 37942
rect 40868 37878 40920 37884
rect 40040 37868 40092 37874
rect 40040 37810 40092 37816
rect 40132 37868 40184 37874
rect 40132 37810 40184 37816
rect 39856 37800 39908 37806
rect 39856 37742 39908 37748
rect 39580 36712 39632 36718
rect 39580 36654 39632 36660
rect 39948 36712 40000 36718
rect 39948 36654 40000 36660
rect 39592 36310 39620 36654
rect 39960 36378 39988 36654
rect 39948 36372 40000 36378
rect 39948 36314 40000 36320
rect 40052 36310 40080 37810
rect 40316 36644 40368 36650
rect 40316 36586 40368 36592
rect 40224 36372 40276 36378
rect 40224 36314 40276 36320
rect 39580 36304 39632 36310
rect 39580 36246 39632 36252
rect 40040 36304 40092 36310
rect 40040 36246 40092 36252
rect 39580 36168 39632 36174
rect 39580 36110 39632 36116
rect 39592 35698 39620 36110
rect 40052 36106 40080 36246
rect 40040 36100 40092 36106
rect 40040 36042 40092 36048
rect 39764 35760 39816 35766
rect 39764 35702 39816 35708
rect 39580 35692 39632 35698
rect 39580 35634 39632 35640
rect 39592 35086 39620 35634
rect 39776 35290 39804 35702
rect 39856 35624 39908 35630
rect 39856 35566 39908 35572
rect 39868 35290 39896 35566
rect 40052 35494 40080 36042
rect 40236 36038 40264 36314
rect 40328 36106 40356 36586
rect 40684 36576 40736 36582
rect 40684 36518 40736 36524
rect 40776 36576 40828 36582
rect 40776 36518 40828 36524
rect 40696 36242 40724 36518
rect 40684 36236 40736 36242
rect 40684 36178 40736 36184
rect 40316 36100 40368 36106
rect 40316 36042 40368 36048
rect 40224 36032 40276 36038
rect 40224 35974 40276 35980
rect 40040 35488 40092 35494
rect 40040 35430 40092 35436
rect 39764 35284 39816 35290
rect 39764 35226 39816 35232
rect 39856 35284 39908 35290
rect 39856 35226 39908 35232
rect 40236 35170 40264 35974
rect 40236 35154 40356 35170
rect 40236 35148 40368 35154
rect 40236 35142 40316 35148
rect 40316 35090 40368 35096
rect 40788 35086 40816 36518
rect 39580 35080 39632 35086
rect 39580 35022 39632 35028
rect 40776 35080 40828 35086
rect 40776 35022 40828 35028
rect 39592 34678 39620 35022
rect 40132 35012 40184 35018
rect 40132 34954 40184 34960
rect 40144 34746 40172 34954
rect 40592 34944 40644 34950
rect 40592 34886 40644 34892
rect 40132 34740 40184 34746
rect 40132 34682 40184 34688
rect 39580 34672 39632 34678
rect 39580 34614 39632 34620
rect 39592 34066 39620 34614
rect 40604 34202 40632 34886
rect 40592 34196 40644 34202
rect 40592 34138 40644 34144
rect 39580 34060 39632 34066
rect 40684 34060 40736 34066
rect 39580 34002 39632 34008
rect 40604 34020 40684 34048
rect 39592 33522 39620 34002
rect 40224 33856 40276 33862
rect 40224 33798 40276 33804
rect 40500 33856 40552 33862
rect 40500 33798 40552 33804
rect 40236 33522 40264 33798
rect 39580 33516 39632 33522
rect 39580 33458 39632 33464
rect 40224 33516 40276 33522
rect 40224 33458 40276 33464
rect 40512 33289 40540 33798
rect 40498 33280 40554 33289
rect 40498 33215 40554 33224
rect 39672 32904 39724 32910
rect 39672 32846 39724 32852
rect 39684 32434 39712 32846
rect 39672 32428 39724 32434
rect 39672 32370 39724 32376
rect 39948 32428 40000 32434
rect 39948 32370 40000 32376
rect 39488 31884 39540 31890
rect 39488 31826 39540 31832
rect 39500 31142 39528 31826
rect 39684 31346 39712 32370
rect 39960 32026 39988 32370
rect 39948 32020 40000 32026
rect 39948 31962 40000 31968
rect 39948 31816 40000 31822
rect 39948 31758 40000 31764
rect 40500 31816 40552 31822
rect 40604 31804 40632 34020
rect 40684 34002 40736 34008
rect 40880 32570 40908 37878
rect 41144 37868 41196 37874
rect 41144 37810 41196 37816
rect 41052 37120 41104 37126
rect 41052 37062 41104 37068
rect 41064 36922 41092 37062
rect 41052 36916 41104 36922
rect 41052 36858 41104 36864
rect 41156 36802 41184 37810
rect 41064 36774 41184 36802
rect 40960 34944 41012 34950
rect 40960 34886 41012 34892
rect 40972 33998 41000 34886
rect 40960 33992 41012 33998
rect 40960 33934 41012 33940
rect 40960 33380 41012 33386
rect 40960 33322 41012 33328
rect 40972 32910 41000 33322
rect 40960 32904 41012 32910
rect 40960 32846 41012 32852
rect 40868 32564 40920 32570
rect 40868 32506 40920 32512
rect 40684 31884 40736 31890
rect 40684 31826 40736 31832
rect 40552 31776 40632 31804
rect 40500 31758 40552 31764
rect 39672 31340 39724 31346
rect 39672 31282 39724 31288
rect 39488 31136 39540 31142
rect 39488 31078 39540 31084
rect 39488 30932 39540 30938
rect 39488 30874 39540 30880
rect 39120 30320 39172 30326
rect 39120 30262 39172 30268
rect 38936 30184 38988 30190
rect 38936 30126 38988 30132
rect 39028 30184 39080 30190
rect 39028 30126 39080 30132
rect 39040 29034 39068 30126
rect 39500 29714 39528 30874
rect 39856 30592 39908 30598
rect 39856 30534 39908 30540
rect 39764 30252 39816 30258
rect 39764 30194 39816 30200
rect 39488 29708 39540 29714
rect 39488 29650 39540 29656
rect 39028 29028 39080 29034
rect 39028 28970 39080 28976
rect 38844 28416 38896 28422
rect 38844 28358 38896 28364
rect 38856 28082 38884 28358
rect 39040 28218 39068 28970
rect 39776 28218 39804 30194
rect 39868 29730 39896 30534
rect 39960 30326 39988 31758
rect 40408 31408 40460 31414
rect 40408 31350 40460 31356
rect 40040 31136 40092 31142
rect 40040 31078 40092 31084
rect 40052 30394 40080 31078
rect 40420 30734 40448 31350
rect 40132 30728 40184 30734
rect 40132 30670 40184 30676
rect 40408 30728 40460 30734
rect 40408 30670 40460 30676
rect 40040 30388 40092 30394
rect 40040 30330 40092 30336
rect 39948 30320 40000 30326
rect 39948 30262 40000 30268
rect 40040 30048 40092 30054
rect 40040 29990 40092 29996
rect 39868 29702 39988 29730
rect 39856 29640 39908 29646
rect 39856 29582 39908 29588
rect 39868 29034 39896 29582
rect 39960 29238 39988 29702
rect 40052 29646 40080 29990
rect 40144 29782 40172 30670
rect 40316 30592 40368 30598
rect 40316 30534 40368 30540
rect 40132 29776 40184 29782
rect 40132 29718 40184 29724
rect 40328 29714 40356 30534
rect 40420 30190 40448 30670
rect 40512 30546 40540 31758
rect 40696 30802 40724 31826
rect 40776 31816 40828 31822
rect 40776 31758 40828 31764
rect 40684 30796 40736 30802
rect 40684 30738 40736 30744
rect 40684 30660 40736 30666
rect 40684 30602 40736 30608
rect 40512 30518 40632 30546
rect 40500 30388 40552 30394
rect 40500 30330 40552 30336
rect 40408 30184 40460 30190
rect 40408 30126 40460 30132
rect 40316 29708 40368 29714
rect 40316 29650 40368 29656
rect 40420 29646 40448 30126
rect 40040 29640 40092 29646
rect 40040 29582 40092 29588
rect 40408 29640 40460 29646
rect 40408 29582 40460 29588
rect 39948 29232 40000 29238
rect 39948 29174 40000 29180
rect 39856 29028 39908 29034
rect 39856 28970 39908 28976
rect 39028 28212 39080 28218
rect 39028 28154 39080 28160
rect 39764 28212 39816 28218
rect 39764 28154 39816 28160
rect 39396 28144 39448 28150
rect 39396 28086 39448 28092
rect 38844 28076 38896 28082
rect 38844 28018 38896 28024
rect 39028 28076 39080 28082
rect 39028 28018 39080 28024
rect 39040 27713 39068 28018
rect 39408 27878 39436 28086
rect 39396 27872 39448 27878
rect 39396 27814 39448 27820
rect 39026 27704 39082 27713
rect 39026 27639 39082 27648
rect 39304 27464 39356 27470
rect 39302 27432 39304 27441
rect 39356 27432 39358 27441
rect 39028 27396 39080 27402
rect 39408 27402 39436 27814
rect 39302 27367 39358 27376
rect 39396 27396 39448 27402
rect 39028 27338 39080 27344
rect 39396 27338 39448 27344
rect 39488 27396 39540 27402
rect 39488 27338 39540 27344
rect 39040 27282 39068 27338
rect 39040 27254 39160 27282
rect 39028 26376 39080 26382
rect 39028 26318 39080 26324
rect 39040 26042 39068 26318
rect 39132 26314 39160 27254
rect 39212 26784 39264 26790
rect 39212 26726 39264 26732
rect 39120 26308 39172 26314
rect 39120 26250 39172 26256
rect 39028 26036 39080 26042
rect 39028 25978 39080 25984
rect 39040 25945 39068 25978
rect 39132 25974 39160 26250
rect 39120 25968 39172 25974
rect 39026 25936 39082 25945
rect 39120 25910 39172 25916
rect 39224 25906 39252 26726
rect 39304 26512 39356 26518
rect 39304 26454 39356 26460
rect 39316 25974 39344 26454
rect 39304 25968 39356 25974
rect 39304 25910 39356 25916
rect 39026 25871 39082 25880
rect 39212 25900 39264 25906
rect 39212 25842 39264 25848
rect 39120 25696 39172 25702
rect 39120 25638 39172 25644
rect 39132 24886 39160 25638
rect 39120 24880 39172 24886
rect 39120 24822 39172 24828
rect 38752 24812 38804 24818
rect 38752 24754 38804 24760
rect 38752 24676 38804 24682
rect 38752 24618 38804 24624
rect 38660 24608 38712 24614
rect 38660 24550 38712 24556
rect 38672 24410 38700 24550
rect 38660 24404 38712 24410
rect 38660 24346 38712 24352
rect 38764 24274 38792 24618
rect 38752 24268 38804 24274
rect 38752 24210 38804 24216
rect 39028 24064 39080 24070
rect 39028 24006 39080 24012
rect 39040 23662 39068 24006
rect 38752 23656 38804 23662
rect 38752 23598 38804 23604
rect 39028 23656 39080 23662
rect 39028 23598 39080 23604
rect 38660 23112 38712 23118
rect 38660 23054 38712 23060
rect 38016 22772 38068 22778
rect 38016 22714 38068 22720
rect 38200 22772 38252 22778
rect 38200 22714 38252 22720
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 37556 22432 37608 22438
rect 37556 22374 37608 22380
rect 37016 22066 37136 22094
rect 36912 20392 36964 20398
rect 36912 20334 36964 20340
rect 36924 19718 36952 20334
rect 36912 19712 36964 19718
rect 36912 19654 36964 19660
rect 36820 13456 36872 13462
rect 36820 13398 36872 13404
rect 36832 12986 36860 13398
rect 36820 12980 36872 12986
rect 36820 12922 36872 12928
rect 36740 12406 36860 12434
rect 36360 12232 36412 12238
rect 36360 12174 36412 12180
rect 36372 11898 36400 12174
rect 36728 12096 36780 12102
rect 36728 12038 36780 12044
rect 36740 11898 36768 12038
rect 36832 11898 36860 12406
rect 36924 12306 36952 19654
rect 37004 17672 37056 17678
rect 37004 17614 37056 17620
rect 37016 16998 37044 17614
rect 37004 16992 37056 16998
rect 37004 16934 37056 16940
rect 37016 16590 37044 16934
rect 37004 16584 37056 16590
rect 37004 16526 37056 16532
rect 37004 15972 37056 15978
rect 37004 15914 37056 15920
rect 36912 12300 36964 12306
rect 36912 12242 36964 12248
rect 36360 11892 36412 11898
rect 36360 11834 36412 11840
rect 36728 11892 36780 11898
rect 36728 11834 36780 11840
rect 36820 11892 36872 11898
rect 36820 11834 36872 11840
rect 36360 11008 36412 11014
rect 36360 10950 36412 10956
rect 36372 10810 36400 10950
rect 36360 10804 36412 10810
rect 36360 10746 36412 10752
rect 36360 10668 36412 10674
rect 36360 10610 36412 10616
rect 36372 9586 36400 10610
rect 36452 10056 36504 10062
rect 36452 9998 36504 10004
rect 36636 10056 36688 10062
rect 36636 9998 36688 10004
rect 36464 9654 36492 9998
rect 36452 9648 36504 9654
rect 36452 9590 36504 9596
rect 36360 9580 36412 9586
rect 36360 9522 36412 9528
rect 36544 9580 36596 9586
rect 36648 9568 36676 9998
rect 37016 9994 37044 15914
rect 37108 15706 37136 22066
rect 37568 20942 37596 22374
rect 37188 20936 37240 20942
rect 37188 20878 37240 20884
rect 37556 20936 37608 20942
rect 37556 20878 37608 20884
rect 37200 20534 37228 20878
rect 37188 20528 37240 20534
rect 37188 20470 37240 20476
rect 37188 19712 37240 19718
rect 37188 19654 37240 19660
rect 37200 18834 37228 19654
rect 37188 18828 37240 18834
rect 37188 18770 37240 18776
rect 37200 18086 37228 18770
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 37188 18080 37240 18086
rect 37188 18022 37240 18028
rect 37476 17678 37504 18158
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37476 16658 37504 17614
rect 37556 17128 37608 17134
rect 37556 17070 37608 17076
rect 37464 16652 37516 16658
rect 37464 16594 37516 16600
rect 37372 16584 37424 16590
rect 37372 16526 37424 16532
rect 37280 15904 37332 15910
rect 37280 15846 37332 15852
rect 37292 15706 37320 15846
rect 37096 15700 37148 15706
rect 37096 15642 37148 15648
rect 37280 15700 37332 15706
rect 37280 15642 37332 15648
rect 37108 15162 37136 15642
rect 37096 15156 37148 15162
rect 37096 15098 37148 15104
rect 37280 15020 37332 15026
rect 37280 14962 37332 14968
rect 37292 14074 37320 14962
rect 37280 14068 37332 14074
rect 37280 14010 37332 14016
rect 37384 13530 37412 16526
rect 37476 16182 37504 16594
rect 37568 16454 37596 17070
rect 37556 16448 37608 16454
rect 37556 16390 37608 16396
rect 37464 16176 37516 16182
rect 37464 16118 37516 16124
rect 37476 15570 37504 16118
rect 37568 15910 37596 16390
rect 37752 16250 37780 22578
rect 38028 22098 38056 22714
rect 38016 22092 38068 22098
rect 38016 22034 38068 22040
rect 38200 21956 38252 21962
rect 38200 21898 38252 21904
rect 37924 20052 37976 20058
rect 37924 19994 37976 20000
rect 37936 19310 37964 19994
rect 38108 19372 38160 19378
rect 38108 19314 38160 19320
rect 37924 19304 37976 19310
rect 37976 19264 38056 19292
rect 37924 19246 37976 19252
rect 37924 18624 37976 18630
rect 37924 18566 37976 18572
rect 37936 18358 37964 18566
rect 37924 18352 37976 18358
rect 37924 18294 37976 18300
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 37844 17338 37872 18158
rect 37832 17332 37884 17338
rect 37832 17274 37884 17280
rect 37936 17134 37964 18294
rect 38028 17762 38056 19264
rect 38120 18970 38148 19314
rect 38108 18964 38160 18970
rect 38108 18906 38160 18912
rect 38028 17734 38148 17762
rect 38016 17604 38068 17610
rect 38016 17546 38068 17552
rect 38028 17338 38056 17546
rect 38016 17332 38068 17338
rect 38016 17274 38068 17280
rect 38016 17196 38068 17202
rect 38016 17138 38068 17144
rect 37924 17128 37976 17134
rect 37924 17070 37976 17076
rect 38028 16794 38056 17138
rect 38016 16788 38068 16794
rect 38016 16730 38068 16736
rect 37740 16244 37792 16250
rect 37740 16186 37792 16192
rect 37556 15904 37608 15910
rect 37556 15846 37608 15852
rect 37464 15564 37516 15570
rect 37464 15506 37516 15512
rect 37476 15162 37504 15506
rect 37464 15156 37516 15162
rect 37464 15098 37516 15104
rect 37476 15026 37504 15098
rect 38028 15094 38056 16730
rect 38120 15978 38148 17734
rect 38212 16590 38240 21898
rect 38672 21146 38700 23054
rect 38764 22030 38792 23598
rect 38752 22024 38804 22030
rect 38752 21966 38804 21972
rect 38660 21140 38712 21146
rect 38660 21082 38712 21088
rect 38764 20890 38792 21966
rect 39224 21010 39252 25842
rect 39408 25838 39436 27338
rect 39500 26246 39528 27338
rect 39580 26308 39632 26314
rect 39580 26250 39632 26256
rect 39488 26240 39540 26246
rect 39488 26182 39540 26188
rect 39396 25832 39448 25838
rect 39396 25774 39448 25780
rect 39592 24886 39620 26250
rect 39580 24880 39632 24886
rect 39580 24822 39632 24828
rect 39592 24750 39620 24822
rect 39580 24744 39632 24750
rect 39580 24686 39632 24692
rect 39592 24206 39620 24686
rect 39672 24608 39724 24614
rect 39672 24550 39724 24556
rect 39580 24200 39632 24206
rect 39486 24168 39542 24177
rect 39304 24132 39356 24138
rect 39580 24142 39632 24148
rect 39486 24103 39488 24112
rect 39304 24074 39356 24080
rect 39540 24103 39542 24112
rect 39488 24074 39540 24080
rect 39316 23322 39344 24074
rect 39304 23316 39356 23322
rect 39304 23258 39356 23264
rect 39394 23216 39450 23225
rect 39394 23151 39450 23160
rect 39408 23118 39436 23151
rect 39396 23112 39448 23118
rect 39396 23054 39448 23060
rect 39396 22500 39448 22506
rect 39396 22442 39448 22448
rect 39408 21010 39436 22442
rect 39212 21004 39264 21010
rect 39212 20946 39264 20952
rect 39396 21004 39448 21010
rect 39396 20946 39448 20952
rect 38672 20862 38792 20890
rect 38476 19780 38528 19786
rect 38476 19722 38528 19728
rect 38488 19514 38516 19722
rect 38672 19718 38700 20862
rect 38752 20800 38804 20806
rect 38752 20742 38804 20748
rect 39580 20800 39632 20806
rect 39580 20742 39632 20748
rect 38764 20466 38792 20742
rect 38752 20460 38804 20466
rect 38752 20402 38804 20408
rect 38844 20460 38896 20466
rect 38844 20402 38896 20408
rect 38856 19922 38884 20402
rect 39028 20256 39080 20262
rect 39028 20198 39080 20204
rect 38844 19916 38896 19922
rect 38844 19858 38896 19864
rect 39040 19854 39068 20198
rect 39028 19848 39080 19854
rect 39028 19790 39080 19796
rect 39592 19718 39620 20742
rect 38660 19712 38712 19718
rect 38660 19654 38712 19660
rect 39580 19712 39632 19718
rect 39580 19654 39632 19660
rect 38476 19508 38528 19514
rect 38476 19450 38528 19456
rect 38672 18426 38700 19654
rect 39592 19446 39620 19654
rect 39580 19440 39632 19446
rect 39580 19382 39632 19388
rect 39304 18760 39356 18766
rect 39304 18702 39356 18708
rect 38660 18420 38712 18426
rect 38660 18362 38712 18368
rect 38672 17610 38700 18362
rect 39316 18086 39344 18702
rect 39304 18080 39356 18086
rect 39304 18022 39356 18028
rect 39580 17808 39632 17814
rect 39580 17750 39632 17756
rect 38660 17604 38712 17610
rect 38660 17546 38712 17552
rect 38476 17196 38528 17202
rect 38476 17138 38528 17144
rect 38568 17196 38620 17202
rect 38568 17138 38620 17144
rect 38488 17066 38516 17138
rect 38476 17060 38528 17066
rect 38476 17002 38528 17008
rect 38200 16584 38252 16590
rect 38200 16526 38252 16532
rect 38108 15972 38160 15978
rect 38108 15914 38160 15920
rect 38016 15088 38068 15094
rect 38016 15030 38068 15036
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37740 14952 37792 14958
rect 37740 14894 37792 14900
rect 37752 14618 37780 14894
rect 38120 14634 38148 15914
rect 38488 15586 38516 17002
rect 38580 16794 38608 17138
rect 38568 16788 38620 16794
rect 38568 16730 38620 16736
rect 38672 15706 38700 17546
rect 38844 17536 38896 17542
rect 38844 17478 38896 17484
rect 38856 17270 38884 17478
rect 38844 17264 38896 17270
rect 38844 17206 38896 17212
rect 39592 17202 39620 17750
rect 39580 17196 39632 17202
rect 39580 17138 39632 17144
rect 39592 16998 39620 17138
rect 39580 16992 39632 16998
rect 39580 16934 39632 16940
rect 39120 16448 39172 16454
rect 39120 16390 39172 16396
rect 38660 15700 38712 15706
rect 38660 15642 38712 15648
rect 38396 15558 38516 15586
rect 38672 15570 38700 15642
rect 38660 15564 38712 15570
rect 37740 14612 37792 14618
rect 38120 14606 38240 14634
rect 37740 14554 37792 14560
rect 38108 14476 38160 14482
rect 38108 14418 38160 14424
rect 37924 14272 37976 14278
rect 37924 14214 37976 14220
rect 37464 13796 37516 13802
rect 37464 13738 37516 13744
rect 37648 13796 37700 13802
rect 37648 13738 37700 13744
rect 37372 13524 37424 13530
rect 37372 13466 37424 13472
rect 37280 13184 37332 13190
rect 37280 13126 37332 13132
rect 37188 12232 37240 12238
rect 37188 12174 37240 12180
rect 37200 11354 37228 12174
rect 37188 11348 37240 11354
rect 37188 11290 37240 11296
rect 37200 10130 37228 11290
rect 37188 10124 37240 10130
rect 37188 10066 37240 10072
rect 37004 9988 37056 9994
rect 37004 9930 37056 9936
rect 36596 9540 36676 9568
rect 36544 9522 36596 9528
rect 36268 9376 36320 9382
rect 36268 9318 36320 9324
rect 36176 8968 36228 8974
rect 36176 8910 36228 8916
rect 35992 8832 36044 8838
rect 35992 8774 36044 8780
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 36004 8378 36032 8774
rect 36084 8492 36136 8498
rect 36084 8434 36136 8440
rect 35912 8350 36032 8378
rect 35912 7818 35940 8350
rect 35992 8288 36044 8294
rect 35992 8230 36044 8236
rect 35900 7812 35952 7818
rect 35900 7754 35952 7760
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 35440 7540 35492 7546
rect 35440 7482 35492 7488
rect 36004 7478 36032 8230
rect 35992 7472 36044 7478
rect 35992 7414 36044 7420
rect 36096 7274 36124 8434
rect 36188 7750 36216 8910
rect 36280 8566 36308 9318
rect 36372 9178 36400 9522
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 36372 9042 36400 9114
rect 36360 9036 36412 9042
rect 36360 8978 36412 8984
rect 36452 9036 36504 9042
rect 36452 8978 36504 8984
rect 36268 8560 36320 8566
rect 36268 8502 36320 8508
rect 36280 7834 36308 8502
rect 36280 7818 36400 7834
rect 36280 7812 36412 7818
rect 36280 7806 36360 7812
rect 36176 7744 36228 7750
rect 36176 7686 36228 7692
rect 36084 7268 36136 7274
rect 36084 7210 36136 7216
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 36004 6798 36032 7142
rect 36188 6866 36216 7686
rect 36176 6860 36228 6866
rect 36176 6802 36228 6808
rect 35992 6792 36044 6798
rect 35992 6734 36044 6740
rect 36280 6730 36308 7806
rect 36360 7754 36412 7760
rect 36464 7698 36492 8978
rect 36544 8492 36596 8498
rect 36544 8434 36596 8440
rect 36372 7670 36492 7698
rect 36372 7410 36400 7670
rect 36556 7478 36584 8434
rect 36544 7472 36596 7478
rect 36544 7414 36596 7420
rect 36360 7404 36412 7410
rect 36360 7346 36412 7352
rect 36452 7404 36504 7410
rect 36452 7346 36504 7352
rect 36372 6798 36400 7346
rect 36464 7002 36492 7346
rect 36544 7336 36596 7342
rect 36544 7278 36596 7284
rect 36452 6996 36504 7002
rect 36452 6938 36504 6944
rect 36360 6792 36412 6798
rect 36360 6734 36412 6740
rect 35440 6724 35492 6730
rect 35440 6666 35492 6672
rect 36268 6724 36320 6730
rect 36268 6666 36320 6672
rect 35452 6390 35480 6666
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 36280 6458 36308 6666
rect 36268 6452 36320 6458
rect 36268 6394 36320 6400
rect 35348 6384 35400 6390
rect 35348 6326 35400 6332
rect 35440 6384 35492 6390
rect 35440 6326 35492 6332
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35256 5568 35308 5574
rect 35256 5510 35308 5516
rect 35268 5234 35296 5510
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 36556 5302 36584 7278
rect 36648 7206 36676 9540
rect 36728 9104 36780 9110
rect 36728 9046 36780 9052
rect 36740 7410 36768 9046
rect 37016 9042 37044 9930
rect 37292 9926 37320 13126
rect 37384 12170 37412 13466
rect 37476 13326 37504 13738
rect 37464 13320 37516 13326
rect 37464 13262 37516 13268
rect 37476 12646 37504 13262
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 37464 12640 37516 12646
rect 37464 12582 37516 12588
rect 37476 12306 37504 12582
rect 37464 12300 37516 12306
rect 37464 12242 37516 12248
rect 37568 12238 37596 12786
rect 37660 12714 37688 13738
rect 37648 12708 37700 12714
rect 37648 12650 37700 12656
rect 37556 12232 37608 12238
rect 37556 12174 37608 12180
rect 37372 12164 37424 12170
rect 37372 12106 37424 12112
rect 37660 11694 37688 12650
rect 37936 12102 37964 14214
rect 38120 13530 38148 14418
rect 38212 13802 38240 14606
rect 38396 14414 38424 15558
rect 38712 15524 38792 15552
rect 38660 15506 38712 15512
rect 38764 15094 38792 15524
rect 39132 15502 39160 16390
rect 39488 16040 39540 16046
rect 39488 15982 39540 15988
rect 39500 15570 39528 15982
rect 39488 15564 39540 15570
rect 39488 15506 39540 15512
rect 39120 15496 39172 15502
rect 39120 15438 39172 15444
rect 39028 15428 39080 15434
rect 39028 15370 39080 15376
rect 38752 15088 38804 15094
rect 38752 15030 38804 15036
rect 38476 14816 38528 14822
rect 38476 14758 38528 14764
rect 38488 14414 38516 14758
rect 38384 14408 38436 14414
rect 38384 14350 38436 14356
rect 38476 14408 38528 14414
rect 38660 14408 38712 14414
rect 38476 14350 38528 14356
rect 38580 14368 38660 14396
rect 38396 14278 38424 14350
rect 38384 14272 38436 14278
rect 38384 14214 38436 14220
rect 38580 14074 38608 14368
rect 38660 14350 38712 14356
rect 38384 14068 38436 14074
rect 38384 14010 38436 14016
rect 38568 14068 38620 14074
rect 38568 14010 38620 14016
rect 38292 13932 38344 13938
rect 38292 13874 38344 13880
rect 38200 13796 38252 13802
rect 38200 13738 38252 13744
rect 38108 13524 38160 13530
rect 38108 13466 38160 13472
rect 38200 12164 38252 12170
rect 38200 12106 38252 12112
rect 37924 12096 37976 12102
rect 37924 12038 37976 12044
rect 37936 11914 37964 12038
rect 37844 11886 37964 11914
rect 37648 11688 37700 11694
rect 37648 11630 37700 11636
rect 37556 11620 37608 11626
rect 37556 11562 37608 11568
rect 37372 10600 37424 10606
rect 37372 10542 37424 10548
rect 37384 10470 37412 10542
rect 37372 10464 37424 10470
rect 37372 10406 37424 10412
rect 37464 10464 37516 10470
rect 37464 10406 37516 10412
rect 37476 9994 37504 10406
rect 37568 10062 37596 11562
rect 37844 11150 37872 11886
rect 37924 11688 37976 11694
rect 37924 11630 37976 11636
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 37832 11008 37884 11014
rect 37832 10950 37884 10956
rect 37844 10606 37872 10950
rect 37936 10674 37964 11630
rect 37924 10668 37976 10674
rect 37924 10610 37976 10616
rect 37832 10600 37884 10606
rect 37832 10542 37884 10548
rect 37648 10532 37700 10538
rect 37648 10474 37700 10480
rect 37660 10062 37688 10474
rect 37556 10056 37608 10062
rect 37556 9998 37608 10004
rect 37648 10056 37700 10062
rect 37648 9998 37700 10004
rect 37464 9988 37516 9994
rect 37464 9930 37516 9936
rect 37280 9920 37332 9926
rect 37280 9862 37332 9868
rect 37004 9036 37056 9042
rect 37004 8978 37056 8984
rect 37292 8974 37320 9862
rect 37660 9722 37688 9998
rect 37648 9716 37700 9722
rect 37648 9658 37700 9664
rect 37096 8968 37148 8974
rect 37096 8910 37148 8916
rect 37280 8968 37332 8974
rect 37280 8910 37332 8916
rect 37464 8968 37516 8974
rect 37464 8910 37516 8916
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 37108 8498 37136 8910
rect 37096 8492 37148 8498
rect 37096 8434 37148 8440
rect 37004 8424 37056 8430
rect 37292 8378 37320 8910
rect 37476 8838 37504 8910
rect 37464 8832 37516 8838
rect 37464 8774 37516 8780
rect 37476 8430 37504 8774
rect 38028 8634 38056 8910
rect 38016 8628 38068 8634
rect 38016 8570 38068 8576
rect 37004 8366 37056 8372
rect 36728 7404 36780 7410
rect 36728 7346 36780 7352
rect 36820 7404 36872 7410
rect 36820 7346 36872 7352
rect 36636 7200 36688 7206
rect 36636 7142 36688 7148
rect 36740 6934 36768 7346
rect 36832 7002 36860 7346
rect 37016 7342 37044 8366
rect 37200 8350 37320 8378
rect 37464 8424 37516 8430
rect 37464 8366 37516 8372
rect 37372 8356 37424 8362
rect 37200 7410 37228 8350
rect 37372 8298 37424 8304
rect 37384 7818 37412 8298
rect 37372 7812 37424 7818
rect 37372 7754 37424 7760
rect 37648 7540 37700 7546
rect 37648 7482 37700 7488
rect 37188 7404 37240 7410
rect 37188 7346 37240 7352
rect 37004 7336 37056 7342
rect 37004 7278 37056 7284
rect 36820 6996 36872 7002
rect 36820 6938 36872 6944
rect 36728 6928 36780 6934
rect 36728 6870 36780 6876
rect 37016 6798 37044 7278
rect 37372 7200 37424 7206
rect 37372 7142 37424 7148
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 37016 5914 37044 6734
rect 37004 5908 37056 5914
rect 37004 5850 37056 5856
rect 37384 5778 37412 7142
rect 37464 6180 37516 6186
rect 37464 6122 37516 6128
rect 37372 5772 37424 5778
rect 37372 5714 37424 5720
rect 36544 5296 36596 5302
rect 36544 5238 36596 5244
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 35256 5228 35308 5234
rect 35256 5170 35308 5176
rect 37476 5166 37504 6122
rect 37660 5778 37688 7482
rect 38212 7478 38240 12106
rect 38304 11014 38332 13874
rect 38396 12442 38424 14010
rect 39040 13530 39068 15370
rect 39132 14414 39160 15438
rect 39212 15360 39264 15366
rect 39212 15302 39264 15308
rect 39304 15360 39356 15366
rect 39304 15302 39356 15308
rect 39224 15094 39252 15302
rect 39212 15088 39264 15094
rect 39212 15030 39264 15036
rect 39224 14414 39252 15030
rect 39120 14408 39172 14414
rect 39120 14350 39172 14356
rect 39212 14408 39264 14414
rect 39212 14350 39264 14356
rect 39132 14278 39160 14350
rect 39120 14272 39172 14278
rect 39120 14214 39172 14220
rect 39316 13938 39344 15302
rect 39500 14414 39528 15506
rect 39580 15496 39632 15502
rect 39580 15438 39632 15444
rect 39592 14618 39620 15438
rect 39580 14612 39632 14618
rect 39580 14554 39632 14560
rect 39592 14482 39620 14554
rect 39580 14476 39632 14482
rect 39580 14418 39632 14424
rect 39488 14408 39540 14414
rect 39488 14350 39540 14356
rect 39500 13938 39528 14350
rect 39120 13932 39172 13938
rect 39120 13874 39172 13880
rect 39304 13932 39356 13938
rect 39304 13874 39356 13880
rect 39488 13932 39540 13938
rect 39488 13874 39540 13880
rect 39028 13524 39080 13530
rect 39028 13466 39080 13472
rect 38476 13252 38528 13258
rect 38476 13194 38528 13200
rect 38488 12646 38516 13194
rect 38568 12980 38620 12986
rect 38568 12922 38620 12928
rect 38476 12640 38528 12646
rect 38476 12582 38528 12588
rect 38384 12436 38436 12442
rect 38384 12378 38436 12384
rect 38488 11694 38516 12582
rect 38476 11688 38528 11694
rect 38476 11630 38528 11636
rect 38580 11626 38608 12922
rect 38844 12776 38896 12782
rect 38844 12718 38896 12724
rect 38856 12306 38884 12718
rect 39040 12306 39068 13466
rect 39132 13326 39160 13874
rect 39212 13864 39264 13870
rect 39212 13806 39264 13812
rect 39224 13326 39252 13806
rect 39396 13728 39448 13734
rect 39396 13670 39448 13676
rect 39408 13530 39436 13670
rect 39396 13524 39448 13530
rect 39396 13466 39448 13472
rect 39120 13320 39172 13326
rect 39120 13262 39172 13268
rect 39212 13320 39264 13326
rect 39212 13262 39264 13268
rect 39132 13190 39160 13262
rect 39120 13184 39172 13190
rect 39120 13126 39172 13132
rect 39408 12986 39436 13466
rect 39488 13320 39540 13326
rect 39488 13262 39540 13268
rect 39396 12980 39448 12986
rect 39396 12922 39448 12928
rect 39212 12776 39264 12782
rect 39132 12736 39212 12764
rect 38844 12300 38896 12306
rect 38844 12242 38896 12248
rect 39028 12300 39080 12306
rect 39028 12242 39080 12248
rect 38934 12200 38990 12209
rect 38934 12135 38936 12144
rect 38988 12135 38990 12144
rect 38936 12106 38988 12112
rect 38384 11620 38436 11626
rect 38384 11562 38436 11568
rect 38568 11620 38620 11626
rect 38568 11562 38620 11568
rect 38396 11218 38424 11562
rect 38384 11212 38436 11218
rect 38384 11154 38436 11160
rect 38292 11008 38344 11014
rect 38292 10950 38344 10956
rect 38396 10690 38424 11154
rect 39132 10810 39160 12736
rect 39212 12718 39264 12724
rect 39212 12640 39264 12646
rect 39212 12582 39264 12588
rect 39304 12640 39356 12646
rect 39304 12582 39356 12588
rect 39224 12238 39252 12582
rect 39212 12232 39264 12238
rect 39212 12174 39264 12180
rect 39316 12170 39344 12582
rect 39500 12442 39528 13262
rect 39396 12436 39448 12442
rect 39396 12378 39448 12384
rect 39488 12436 39540 12442
rect 39488 12378 39540 12384
rect 39408 12322 39436 12378
rect 39580 12368 39632 12374
rect 39408 12316 39580 12322
rect 39408 12310 39632 12316
rect 39408 12294 39620 12310
rect 39580 12232 39632 12238
rect 39408 12192 39580 12220
rect 39304 12164 39356 12170
rect 39304 12106 39356 12112
rect 39212 12096 39264 12102
rect 39408 12050 39436 12192
rect 39580 12174 39632 12180
rect 39264 12044 39436 12050
rect 39212 12038 39436 12044
rect 39224 12022 39436 12038
rect 39120 10804 39172 10810
rect 39120 10746 39172 10752
rect 38476 10736 38528 10742
rect 38396 10684 38476 10690
rect 38396 10678 38528 10684
rect 38396 10662 38516 10678
rect 38396 9722 38424 10662
rect 38568 10600 38620 10606
rect 38568 10542 38620 10548
rect 38936 10600 38988 10606
rect 38936 10542 38988 10548
rect 38580 10266 38608 10542
rect 38844 10464 38896 10470
rect 38844 10406 38896 10412
rect 38568 10260 38620 10266
rect 38568 10202 38620 10208
rect 38856 10062 38884 10406
rect 38948 10062 38976 10542
rect 38844 10056 38896 10062
rect 38844 9998 38896 10004
rect 38936 10056 38988 10062
rect 38936 9998 38988 10004
rect 38660 9920 38712 9926
rect 38660 9862 38712 9868
rect 38384 9716 38436 9722
rect 38384 9658 38436 9664
rect 38396 9602 38424 9658
rect 38672 9654 38700 9862
rect 38304 9574 38424 9602
rect 38660 9648 38712 9654
rect 38660 9590 38712 9596
rect 38304 8566 38332 9574
rect 38660 9512 38712 9518
rect 38712 9472 38884 9500
rect 38660 9454 38712 9460
rect 38568 9444 38620 9450
rect 38568 9386 38620 9392
rect 38580 9330 38608 9386
rect 38580 9302 38700 9330
rect 38672 8974 38700 9302
rect 38660 8968 38712 8974
rect 38660 8910 38712 8916
rect 38476 8832 38528 8838
rect 38476 8774 38528 8780
rect 38488 8634 38516 8774
rect 38476 8628 38528 8634
rect 38476 8570 38528 8576
rect 38292 8560 38344 8566
rect 38292 8502 38344 8508
rect 38200 7472 38252 7478
rect 38200 7414 38252 7420
rect 37740 6792 37792 6798
rect 37740 6734 37792 6740
rect 37752 6458 37780 6734
rect 38304 6730 38332 8502
rect 38672 8090 38700 8910
rect 38856 8548 38884 9472
rect 38948 8906 38976 9998
rect 38936 8900 38988 8906
rect 38936 8842 38988 8848
rect 38936 8560 38988 8566
rect 38856 8520 38936 8548
rect 38936 8502 38988 8508
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 38948 7954 38976 8502
rect 38936 7948 38988 7954
rect 38936 7890 38988 7896
rect 38660 7880 38712 7886
rect 38660 7822 38712 7828
rect 38672 7478 38700 7822
rect 38948 7546 38976 7890
rect 38936 7540 38988 7546
rect 38936 7482 38988 7488
rect 38660 7472 38712 7478
rect 38660 7414 38712 7420
rect 39684 7410 39712 24550
rect 39776 24274 39804 28154
rect 39868 27402 39896 28970
rect 39960 28490 39988 29174
rect 40420 29102 40448 29582
rect 40512 29510 40540 30330
rect 40604 30190 40632 30518
rect 40592 30184 40644 30190
rect 40592 30126 40644 30132
rect 40696 29850 40724 30602
rect 40684 29844 40736 29850
rect 40684 29786 40736 29792
rect 40788 29578 40816 31758
rect 41064 31482 41092 36774
rect 41248 36718 41276 38966
rect 41328 38888 41380 38894
rect 41328 38830 41380 38836
rect 41340 38010 41368 38830
rect 42168 38554 42196 39374
rect 41420 38548 41472 38554
rect 41420 38490 41472 38496
rect 42156 38548 42208 38554
rect 42156 38490 42208 38496
rect 41328 38004 41380 38010
rect 41328 37946 41380 37952
rect 41144 36712 41196 36718
rect 41144 36654 41196 36660
rect 41236 36712 41288 36718
rect 41236 36654 41288 36660
rect 41156 34746 41184 36654
rect 41248 36378 41276 36654
rect 41328 36644 41380 36650
rect 41328 36586 41380 36592
rect 41236 36372 41288 36378
rect 41236 36314 41288 36320
rect 41340 35834 41368 36586
rect 41432 36106 41460 38490
rect 42168 38214 42196 38490
rect 42156 38208 42208 38214
rect 42156 38150 42208 38156
rect 41696 37800 41748 37806
rect 41696 37742 41748 37748
rect 41420 36100 41472 36106
rect 41420 36042 41472 36048
rect 41328 35828 41380 35834
rect 41328 35770 41380 35776
rect 41432 35766 41460 36042
rect 41420 35760 41472 35766
rect 41420 35702 41472 35708
rect 41236 35624 41288 35630
rect 41236 35566 41288 35572
rect 41248 34746 41276 35566
rect 41432 35290 41460 35702
rect 41420 35284 41472 35290
rect 41420 35226 41472 35232
rect 41328 35080 41380 35086
rect 41328 35022 41380 35028
rect 41340 34746 41368 35022
rect 41144 34740 41196 34746
rect 41144 34682 41196 34688
rect 41236 34740 41288 34746
rect 41236 34682 41288 34688
rect 41328 34740 41380 34746
rect 41328 34682 41380 34688
rect 41248 33862 41276 34682
rect 41340 33998 41368 34682
rect 41708 34678 41736 37742
rect 42156 37256 42208 37262
rect 42156 37198 42208 37204
rect 42168 36786 42196 37198
rect 42156 36780 42208 36786
rect 42156 36722 42208 36728
rect 42168 36378 42196 36722
rect 42156 36372 42208 36378
rect 42156 36314 42208 36320
rect 42156 35488 42208 35494
rect 42156 35430 42208 35436
rect 41788 35080 41840 35086
rect 41788 35022 41840 35028
rect 41696 34672 41748 34678
rect 41696 34614 41748 34620
rect 41708 34066 41736 34614
rect 41696 34060 41748 34066
rect 41696 34002 41748 34008
rect 41328 33992 41380 33998
rect 41328 33934 41380 33940
rect 41236 33856 41288 33862
rect 41236 33798 41288 33804
rect 41248 33114 41276 33798
rect 41340 33658 41368 33934
rect 41328 33652 41380 33658
rect 41328 33594 41380 33600
rect 41604 33516 41656 33522
rect 41604 33458 41656 33464
rect 41236 33108 41288 33114
rect 41236 33050 41288 33056
rect 41144 32224 41196 32230
rect 41144 32166 41196 32172
rect 41156 31958 41184 32166
rect 41144 31952 41196 31958
rect 41144 31894 41196 31900
rect 41420 31816 41472 31822
rect 41420 31758 41472 31764
rect 41052 31476 41104 31482
rect 41052 31418 41104 31424
rect 40960 31340 41012 31346
rect 40960 31282 41012 31288
rect 40972 30394 41000 31282
rect 41236 31136 41288 31142
rect 41236 31078 41288 31084
rect 41248 30394 41276 31078
rect 41432 30938 41460 31758
rect 41420 30932 41472 30938
rect 41420 30874 41472 30880
rect 40960 30388 41012 30394
rect 40960 30330 41012 30336
rect 41236 30388 41288 30394
rect 41236 30330 41288 30336
rect 40776 29572 40828 29578
rect 40776 29514 40828 29520
rect 40500 29504 40552 29510
rect 40500 29446 40552 29452
rect 40132 29096 40184 29102
rect 40132 29038 40184 29044
rect 40408 29096 40460 29102
rect 40408 29038 40460 29044
rect 40144 28558 40172 29038
rect 40684 29028 40736 29034
rect 40684 28970 40736 28976
rect 40696 28626 40724 28970
rect 40684 28620 40736 28626
rect 40684 28562 40736 28568
rect 40132 28552 40184 28558
rect 40132 28494 40184 28500
rect 39948 28484 40000 28490
rect 39948 28426 40000 28432
rect 39960 27402 39988 28426
rect 40040 28076 40092 28082
rect 40040 28018 40092 28024
rect 40052 27606 40080 28018
rect 40040 27600 40092 27606
rect 40040 27542 40092 27548
rect 40144 27470 40172 28494
rect 41512 28416 41564 28422
rect 41512 28358 41564 28364
rect 41524 28082 41552 28358
rect 41512 28076 41564 28082
rect 41512 28018 41564 28024
rect 40408 27872 40460 27878
rect 40408 27814 40460 27820
rect 40592 27872 40644 27878
rect 40592 27814 40644 27820
rect 40132 27464 40184 27470
rect 40132 27406 40184 27412
rect 39856 27396 39908 27402
rect 39856 27338 39908 27344
rect 39948 27396 40000 27402
rect 39948 27338 40000 27344
rect 39960 26314 39988 27338
rect 40038 27160 40094 27169
rect 40038 27095 40040 27104
rect 40092 27095 40094 27104
rect 40040 27066 40092 27072
rect 40040 26580 40092 26586
rect 40040 26522 40092 26528
rect 39948 26308 40000 26314
rect 39948 26250 40000 26256
rect 40052 26042 40080 26522
rect 40144 26450 40172 27406
rect 40132 26444 40184 26450
rect 40132 26386 40184 26392
rect 40224 26240 40276 26246
rect 40224 26182 40276 26188
rect 40040 26036 40092 26042
rect 40040 25978 40092 25984
rect 40052 25906 40080 25978
rect 40236 25906 40264 26182
rect 40316 26036 40368 26042
rect 40316 25978 40368 25984
rect 40040 25900 40092 25906
rect 40040 25842 40092 25848
rect 40132 25900 40184 25906
rect 40132 25842 40184 25848
rect 40224 25900 40276 25906
rect 40224 25842 40276 25848
rect 39764 24268 39816 24274
rect 39764 24210 39816 24216
rect 40040 24200 40092 24206
rect 40040 24142 40092 24148
rect 39764 24064 39816 24070
rect 39764 24006 39816 24012
rect 39776 23798 39804 24006
rect 39764 23792 39816 23798
rect 40052 23769 40080 24142
rect 39764 23734 39816 23740
rect 40038 23760 40094 23769
rect 40038 23695 40094 23704
rect 40052 23118 40080 23695
rect 40144 23225 40172 25842
rect 40236 25770 40264 25842
rect 40224 25764 40276 25770
rect 40224 25706 40276 25712
rect 40224 24064 40276 24070
rect 40224 24006 40276 24012
rect 40236 23905 40264 24006
rect 40222 23896 40278 23905
rect 40222 23831 40278 23840
rect 40130 23216 40186 23225
rect 40130 23151 40186 23160
rect 40040 23112 40092 23118
rect 40040 23054 40092 23060
rect 40328 22778 40356 25978
rect 40420 24834 40448 27814
rect 40604 27674 40632 27814
rect 40592 27668 40644 27674
rect 40592 27610 40644 27616
rect 41616 27130 41644 33458
rect 41800 31906 41828 35022
rect 41880 34604 41932 34610
rect 41880 34546 41932 34552
rect 41892 33930 41920 34546
rect 41972 34128 42024 34134
rect 41972 34070 42024 34076
rect 41880 33924 41932 33930
rect 41880 33866 41932 33872
rect 41984 33454 42012 34070
rect 42168 33658 42196 35430
rect 42156 33652 42208 33658
rect 42156 33594 42208 33600
rect 41972 33448 42024 33454
rect 41972 33390 42024 33396
rect 42156 32428 42208 32434
rect 42156 32370 42208 32376
rect 42064 32224 42116 32230
rect 42064 32166 42116 32172
rect 41708 31878 41828 31906
rect 41708 31754 41736 31878
rect 41708 31726 41920 31754
rect 41788 30932 41840 30938
rect 41788 30874 41840 30880
rect 41800 30258 41828 30874
rect 41788 30252 41840 30258
rect 41788 30194 41840 30200
rect 41696 29572 41748 29578
rect 41696 29514 41748 29520
rect 41708 28490 41736 29514
rect 41892 29322 41920 31726
rect 41972 30048 42024 30054
rect 41970 30016 41972 30025
rect 42024 30016 42026 30025
rect 41970 29951 42026 29960
rect 42076 29345 42104 32166
rect 42168 31822 42196 32370
rect 42156 31816 42208 31822
rect 42156 31758 42208 31764
rect 42168 29850 42196 31758
rect 42156 29844 42208 29850
rect 42156 29786 42208 29792
rect 42062 29336 42118 29345
rect 41892 29294 42012 29322
rect 41880 29164 41932 29170
rect 41880 29106 41932 29112
rect 41892 28762 41920 29106
rect 41880 28756 41932 28762
rect 41880 28698 41932 28704
rect 41696 28484 41748 28490
rect 41696 28426 41748 28432
rect 41708 28098 41736 28426
rect 41708 28070 41828 28098
rect 41694 27976 41750 27985
rect 41694 27911 41696 27920
rect 41748 27911 41750 27920
rect 41696 27882 41748 27888
rect 40868 27124 40920 27130
rect 40868 27066 40920 27072
rect 41604 27124 41656 27130
rect 41604 27066 41656 27072
rect 40592 26988 40644 26994
rect 40592 26930 40644 26936
rect 40776 26988 40828 26994
rect 40776 26930 40828 26936
rect 40604 26042 40632 26930
rect 40788 26897 40816 26930
rect 40774 26888 40830 26897
rect 40774 26823 40830 26832
rect 40684 26784 40736 26790
rect 40684 26726 40736 26732
rect 40696 26450 40724 26726
rect 40684 26444 40736 26450
rect 40684 26386 40736 26392
rect 40880 26330 40908 27066
rect 41052 26988 41104 26994
rect 41052 26930 41104 26936
rect 41064 26450 41092 26930
rect 41236 26852 41288 26858
rect 41236 26794 41288 26800
rect 41052 26444 41104 26450
rect 41052 26386 41104 26392
rect 40696 26302 40908 26330
rect 40592 26036 40644 26042
rect 40592 25978 40644 25984
rect 40500 25900 40552 25906
rect 40552 25860 40632 25888
rect 40500 25842 40552 25848
rect 40604 25294 40632 25860
rect 40592 25288 40644 25294
rect 40592 25230 40644 25236
rect 40500 25220 40552 25226
rect 40500 25162 40552 25168
rect 40512 24954 40540 25162
rect 40500 24948 40552 24954
rect 40500 24890 40552 24896
rect 40420 24806 40540 24834
rect 40408 24200 40460 24206
rect 40408 24142 40460 24148
rect 40420 23866 40448 24142
rect 40408 23860 40460 23866
rect 40408 23802 40460 23808
rect 40408 23112 40460 23118
rect 40408 23054 40460 23060
rect 40316 22772 40368 22778
rect 40316 22714 40368 22720
rect 40132 22432 40184 22438
rect 40132 22374 40184 22380
rect 40144 21962 40172 22374
rect 40420 22030 40448 23054
rect 40408 22024 40460 22030
rect 40408 21966 40460 21972
rect 40132 21956 40184 21962
rect 40132 21898 40184 21904
rect 40420 21622 40448 21966
rect 40408 21616 40460 21622
rect 40408 21558 40460 21564
rect 40224 21344 40276 21350
rect 40224 21286 40276 21292
rect 40040 21004 40092 21010
rect 40040 20946 40092 20952
rect 40052 20754 40080 20946
rect 39960 20726 40080 20754
rect 39960 20534 39988 20726
rect 40236 20602 40264 21286
rect 40420 21010 40448 21558
rect 40408 21004 40460 21010
rect 40408 20946 40460 20952
rect 40408 20868 40460 20874
rect 40408 20810 40460 20816
rect 40224 20596 40276 20602
rect 40224 20538 40276 20544
rect 39948 20528 40000 20534
rect 39948 20470 40000 20476
rect 40420 20398 40448 20810
rect 40512 20534 40540 24806
rect 40604 24750 40632 25230
rect 40592 24744 40644 24750
rect 40592 24686 40644 24692
rect 40696 24138 40724 26302
rect 40776 25968 40828 25974
rect 40776 25910 40828 25916
rect 40788 25838 40816 25910
rect 41064 25906 41092 26386
rect 40868 25900 40920 25906
rect 40868 25842 40920 25848
rect 41052 25900 41104 25906
rect 41052 25842 41104 25848
rect 40776 25832 40828 25838
rect 40776 25774 40828 25780
rect 40880 25770 40908 25842
rect 40868 25764 40920 25770
rect 40868 25706 40920 25712
rect 40776 25152 40828 25158
rect 40776 25094 40828 25100
rect 40788 24274 40816 25094
rect 40880 24954 40908 25706
rect 40960 25696 41012 25702
rect 40960 25638 41012 25644
rect 40972 25226 41000 25638
rect 40960 25220 41012 25226
rect 40960 25162 41012 25168
rect 40868 24948 40920 24954
rect 40868 24890 40920 24896
rect 40958 24848 41014 24857
rect 40868 24812 40920 24818
rect 40958 24783 40960 24792
rect 40868 24754 40920 24760
rect 41012 24783 41014 24792
rect 40960 24754 41012 24760
rect 40880 24721 40908 24754
rect 40866 24712 40922 24721
rect 40866 24647 40922 24656
rect 40776 24268 40828 24274
rect 40776 24210 40828 24216
rect 40684 24132 40736 24138
rect 40684 24074 40736 24080
rect 41052 23792 41104 23798
rect 41052 23734 41104 23740
rect 41142 23760 41198 23769
rect 41064 23032 41092 23734
rect 41142 23695 41144 23704
rect 41196 23695 41198 23704
rect 41248 23712 41276 26794
rect 41800 25498 41828 28070
rect 41880 28076 41932 28082
rect 41880 28018 41932 28024
rect 41892 27674 41920 28018
rect 41880 27668 41932 27674
rect 41880 27610 41932 27616
rect 41878 25936 41934 25945
rect 41878 25871 41880 25880
rect 41932 25871 41934 25880
rect 41880 25842 41932 25848
rect 41788 25492 41840 25498
rect 41788 25434 41840 25440
rect 41510 25256 41566 25265
rect 41510 25191 41566 25200
rect 41524 25158 41552 25191
rect 41512 25152 41564 25158
rect 41512 25094 41564 25100
rect 41604 25152 41656 25158
rect 41604 25094 41656 25100
rect 41328 24812 41380 24818
rect 41328 24754 41380 24760
rect 41340 24410 41368 24754
rect 41616 24698 41644 25094
rect 41800 24886 41828 25434
rect 41984 25226 42012 29294
rect 42062 29271 42118 29280
rect 42064 29028 42116 29034
rect 42064 28970 42116 28976
rect 42076 28665 42104 28970
rect 42062 28656 42118 28665
rect 42062 28591 42118 28600
rect 42064 27872 42116 27878
rect 42064 27814 42116 27820
rect 42076 27305 42104 27814
rect 42062 27296 42118 27305
rect 42062 27231 42118 27240
rect 42064 26784 42116 26790
rect 42064 26726 42116 26732
rect 42076 26625 42104 26726
rect 42062 26616 42118 26625
rect 42062 26551 42118 26560
rect 42064 26036 42116 26042
rect 42064 25978 42116 25984
rect 42076 25945 42104 25978
rect 42062 25936 42118 25945
rect 42062 25871 42118 25880
rect 41972 25220 42024 25226
rect 41972 25162 42024 25168
rect 41696 24880 41748 24886
rect 41696 24822 41748 24828
rect 41788 24880 41840 24886
rect 41788 24822 41840 24828
rect 41432 24670 41644 24698
rect 41432 24614 41460 24670
rect 41420 24608 41472 24614
rect 41512 24608 41564 24614
rect 41420 24550 41472 24556
rect 41510 24576 41512 24585
rect 41564 24576 41566 24585
rect 41510 24511 41566 24520
rect 41328 24404 41380 24410
rect 41328 24346 41380 24352
rect 41708 23798 41736 24822
rect 41788 24676 41840 24682
rect 41788 24618 41840 24624
rect 41800 24206 41828 24618
rect 41788 24200 41840 24206
rect 41788 24142 41840 24148
rect 41696 23792 41748 23798
rect 41696 23734 41748 23740
rect 41420 23724 41472 23730
rect 41144 23666 41196 23672
rect 41248 23684 41420 23712
rect 41144 23044 41196 23050
rect 41064 23004 41144 23032
rect 41144 22986 41196 22992
rect 40960 22636 41012 22642
rect 40960 22578 41012 22584
rect 40972 22438 41000 22578
rect 41156 22522 41184 22986
rect 41248 22778 41276 23684
rect 41420 23666 41472 23672
rect 41604 23724 41656 23730
rect 41604 23666 41656 23672
rect 41328 23520 41380 23526
rect 41328 23462 41380 23468
rect 41340 22982 41368 23462
rect 41616 23225 41644 23666
rect 41708 23322 41736 23734
rect 42064 23724 42116 23730
rect 42064 23666 42116 23672
rect 41696 23316 41748 23322
rect 41696 23258 41748 23264
rect 41602 23216 41658 23225
rect 41602 23151 41658 23160
rect 42076 22982 42104 23666
rect 42154 23216 42210 23225
rect 42154 23151 42210 23160
rect 41328 22976 41380 22982
rect 41328 22918 41380 22924
rect 42064 22976 42116 22982
rect 42064 22918 42116 22924
rect 41236 22772 41288 22778
rect 41236 22714 41288 22720
rect 42076 22710 42104 22918
rect 42064 22704 42116 22710
rect 42064 22646 42116 22652
rect 41972 22636 42024 22642
rect 41972 22578 42024 22584
rect 41328 22568 41380 22574
rect 41156 22494 41276 22522
rect 41328 22510 41380 22516
rect 40684 22432 40736 22438
rect 40684 22374 40736 22380
rect 40960 22432 41012 22438
rect 40960 22374 41012 22380
rect 41144 22432 41196 22438
rect 41144 22374 41196 22380
rect 40696 21554 40724 22374
rect 40684 21548 40736 21554
rect 40684 21490 40736 21496
rect 40960 21344 41012 21350
rect 40960 21286 41012 21292
rect 40684 20868 40736 20874
rect 40684 20810 40736 20816
rect 40696 20602 40724 20810
rect 40684 20596 40736 20602
rect 40684 20538 40736 20544
rect 40500 20528 40552 20534
rect 40500 20470 40552 20476
rect 40972 20466 41000 21286
rect 40960 20460 41012 20466
rect 40960 20402 41012 20408
rect 40408 20392 40460 20398
rect 40408 20334 40460 20340
rect 40224 19780 40276 19786
rect 40224 19722 40276 19728
rect 40236 19514 40264 19722
rect 40868 19712 40920 19718
rect 40868 19654 40920 19660
rect 40224 19508 40276 19514
rect 40224 19450 40276 19456
rect 40880 19378 40908 19654
rect 40972 19514 41000 20402
rect 40960 19508 41012 19514
rect 40960 19450 41012 19456
rect 40592 19372 40644 19378
rect 40592 19314 40644 19320
rect 40868 19372 40920 19378
rect 40868 19314 40920 19320
rect 40604 18970 40632 19314
rect 40592 18964 40644 18970
rect 40592 18906 40644 18912
rect 40880 18766 40908 19314
rect 41052 19236 41104 19242
rect 41052 19178 41104 19184
rect 40868 18760 40920 18766
rect 40868 18702 40920 18708
rect 41064 18698 41092 19178
rect 41052 18692 41104 18698
rect 41052 18634 41104 18640
rect 40224 18624 40276 18630
rect 40224 18566 40276 18572
rect 40236 18358 40264 18566
rect 41064 18426 41092 18634
rect 41052 18420 41104 18426
rect 41052 18362 41104 18368
rect 40224 18352 40276 18358
rect 40224 18294 40276 18300
rect 41064 17746 41092 18362
rect 39948 17740 40000 17746
rect 39948 17682 40000 17688
rect 41052 17740 41104 17746
rect 41052 17682 41104 17688
rect 39856 17672 39908 17678
rect 39856 17614 39908 17620
rect 39868 17202 39896 17614
rect 39960 17202 39988 17682
rect 40052 17462 40264 17490
rect 40052 17338 40080 17462
rect 40040 17332 40092 17338
rect 40040 17274 40092 17280
rect 40132 17332 40184 17338
rect 40132 17274 40184 17280
rect 39856 17196 39908 17202
rect 39856 17138 39908 17144
rect 39948 17196 40000 17202
rect 39948 17138 40000 17144
rect 39868 15570 39896 17138
rect 40144 16590 40172 17274
rect 40132 16584 40184 16590
rect 40132 16526 40184 16532
rect 40040 16448 40092 16454
rect 40040 16390 40092 16396
rect 40052 16114 40080 16390
rect 40144 16114 40172 16526
rect 40040 16108 40092 16114
rect 40040 16050 40092 16056
rect 40132 16108 40184 16114
rect 40132 16050 40184 16056
rect 40236 16046 40264 17462
rect 40408 16992 40460 16998
rect 40408 16934 40460 16940
rect 40500 16992 40552 16998
rect 40500 16934 40552 16940
rect 40224 16040 40276 16046
rect 40224 15982 40276 15988
rect 39856 15564 39908 15570
rect 39856 15506 39908 15512
rect 40420 15502 40448 16934
rect 40512 16658 40540 16934
rect 40500 16652 40552 16658
rect 40500 16594 40552 16600
rect 40500 16516 40552 16522
rect 40500 16458 40552 16464
rect 40512 16046 40540 16458
rect 40500 16040 40552 16046
rect 40500 15982 40552 15988
rect 40040 15496 40092 15502
rect 40408 15496 40460 15502
rect 40092 15456 40172 15484
rect 40040 15438 40092 15444
rect 40040 15360 40092 15366
rect 40040 15302 40092 15308
rect 39856 15088 39908 15094
rect 39856 15030 39908 15036
rect 39868 14414 39896 15030
rect 40052 14482 40080 15302
rect 40144 14890 40172 15456
rect 40408 15438 40460 15444
rect 40132 14884 40184 14890
rect 40132 14826 40184 14832
rect 40040 14476 40092 14482
rect 40040 14418 40092 14424
rect 39764 14408 39816 14414
rect 39764 14350 39816 14356
rect 39856 14408 39908 14414
rect 39856 14350 39908 14356
rect 39776 14006 39804 14350
rect 39764 14000 39816 14006
rect 39764 13942 39816 13948
rect 39764 13864 39816 13870
rect 39868 13818 39896 14350
rect 39948 14068 40000 14074
rect 39948 14010 40000 14016
rect 39816 13812 39896 13818
rect 39764 13806 39896 13812
rect 39776 13790 39896 13806
rect 39960 12306 39988 14010
rect 40224 13184 40276 13190
rect 40224 13126 40276 13132
rect 39948 12300 40000 12306
rect 39948 12242 40000 12248
rect 40236 12238 40264 13126
rect 40420 12850 40448 15438
rect 40868 14952 40920 14958
rect 40868 14894 40920 14900
rect 40880 14618 40908 14894
rect 40868 14612 40920 14618
rect 40868 14554 40920 14560
rect 41156 14074 41184 22374
rect 41248 20874 41276 22494
rect 41340 22234 41368 22510
rect 41328 22228 41380 22234
rect 41328 22170 41380 22176
rect 41984 22098 42012 22578
rect 42168 22506 42196 23151
rect 42156 22500 42208 22506
rect 42156 22442 42208 22448
rect 41972 22092 42024 22098
rect 41972 22034 42024 22040
rect 41328 22024 41380 22030
rect 41328 21966 41380 21972
rect 41340 21690 41368 21966
rect 41328 21684 41380 21690
rect 41328 21626 41380 21632
rect 41236 20868 41288 20874
rect 41236 20810 41288 20816
rect 41248 19786 41276 20810
rect 41984 20602 42012 22034
rect 42156 20800 42208 20806
rect 42156 20742 42208 20748
rect 41972 20596 42024 20602
rect 41972 20538 42024 20544
rect 41512 20460 41564 20466
rect 41512 20402 41564 20408
rect 41236 19780 41288 19786
rect 41236 19722 41288 19728
rect 41248 19334 41276 19722
rect 41524 19514 41552 20402
rect 41696 20392 41748 20398
rect 41696 20334 41748 20340
rect 41708 20058 41736 20334
rect 41696 20052 41748 20058
rect 41696 19994 41748 20000
rect 41512 19508 41564 19514
rect 41512 19450 41564 19456
rect 41248 19306 41552 19334
rect 42168 19310 42196 20742
rect 41328 19168 41380 19174
rect 41328 19110 41380 19116
rect 41340 18222 41368 19110
rect 41328 18216 41380 18222
rect 41328 18158 41380 18164
rect 41340 16114 41368 18158
rect 41420 18080 41472 18086
rect 41420 18022 41472 18028
rect 41432 17678 41460 18022
rect 41420 17672 41472 17678
rect 41420 17614 41472 17620
rect 41328 16108 41380 16114
rect 41328 16050 41380 16056
rect 41420 15496 41472 15502
rect 41420 15438 41472 15444
rect 41432 15162 41460 15438
rect 41420 15156 41472 15162
rect 41420 15098 41472 15104
rect 41144 14068 41196 14074
rect 41144 14010 41196 14016
rect 41432 14006 41460 15098
rect 41524 14414 41552 19306
rect 42156 19304 42208 19310
rect 42156 19246 42208 19252
rect 42064 18896 42116 18902
rect 42064 18838 42116 18844
rect 41604 18760 41656 18766
rect 41604 18702 41656 18708
rect 41616 17882 41644 18702
rect 42076 18358 42104 18838
rect 42064 18352 42116 18358
rect 42064 18294 42116 18300
rect 41696 18080 41748 18086
rect 41696 18022 41748 18028
rect 41604 17876 41656 17882
rect 41604 17818 41656 17824
rect 41708 17066 41736 18022
rect 42168 17202 42196 19246
rect 42248 18352 42300 18358
rect 42248 18294 42300 18300
rect 41972 17196 42024 17202
rect 41972 17138 42024 17144
rect 42156 17196 42208 17202
rect 42156 17138 42208 17144
rect 41696 17060 41748 17066
rect 41696 17002 41748 17008
rect 41604 16584 41656 16590
rect 41604 16526 41656 16532
rect 41616 15706 41644 16526
rect 41984 16454 42012 17138
rect 42168 16776 42196 17138
rect 42076 16748 42196 16776
rect 41972 16448 42024 16454
rect 41972 16390 42024 16396
rect 41984 16182 42012 16390
rect 41972 16176 42024 16182
rect 41972 16118 42024 16124
rect 42076 16114 42104 16748
rect 42064 16108 42116 16114
rect 42064 16050 42116 16056
rect 42260 16046 42288 18294
rect 42248 16040 42300 16046
rect 42248 15982 42300 15988
rect 41604 15700 41656 15706
rect 41604 15642 41656 15648
rect 41616 14958 41644 15642
rect 41788 15428 41840 15434
rect 41788 15370 41840 15376
rect 41604 14952 41656 14958
rect 41604 14894 41656 14900
rect 41800 14618 41828 15370
rect 41788 14612 41840 14618
rect 41788 14554 41840 14560
rect 41512 14408 41564 14414
rect 41512 14350 41564 14356
rect 41420 14000 41472 14006
rect 41420 13942 41472 13948
rect 40776 13796 40828 13802
rect 40776 13738 40828 13744
rect 40684 13728 40736 13734
rect 40684 13670 40736 13676
rect 40696 13394 40724 13670
rect 40684 13388 40736 13394
rect 40684 13330 40736 13336
rect 40500 12912 40552 12918
rect 40500 12854 40552 12860
rect 40408 12844 40460 12850
rect 40408 12786 40460 12792
rect 40512 12306 40540 12854
rect 40684 12776 40736 12782
rect 40684 12718 40736 12724
rect 40696 12306 40724 12718
rect 40500 12300 40552 12306
rect 40500 12242 40552 12248
rect 40684 12300 40736 12306
rect 40684 12242 40736 12248
rect 40224 12232 40276 12238
rect 39762 12200 39818 12209
rect 40224 12174 40276 12180
rect 39762 12135 39764 12144
rect 39816 12135 39818 12144
rect 39764 12106 39816 12112
rect 40592 12096 40644 12102
rect 40592 12038 40644 12044
rect 40604 11898 40632 12038
rect 40696 11898 40724 12242
rect 40592 11892 40644 11898
rect 40592 11834 40644 11840
rect 40684 11892 40736 11898
rect 40684 11834 40736 11840
rect 39948 10804 40000 10810
rect 39948 10746 40000 10752
rect 39960 9994 39988 10746
rect 40788 10674 40816 13738
rect 41144 13252 41196 13258
rect 41144 13194 41196 13200
rect 41156 11762 41184 13194
rect 41524 13002 41552 14350
rect 42156 13864 42208 13870
rect 42156 13806 42208 13812
rect 42168 13530 42196 13806
rect 42156 13524 42208 13530
rect 42156 13466 42208 13472
rect 41432 12974 41552 13002
rect 41144 11756 41196 11762
rect 41144 11698 41196 11704
rect 40776 10668 40828 10674
rect 40776 10610 40828 10616
rect 40408 10056 40460 10062
rect 40408 9998 40460 10004
rect 39948 9988 40000 9994
rect 39948 9930 40000 9936
rect 40420 9518 40448 9998
rect 40408 9512 40460 9518
rect 40408 9454 40460 9460
rect 39764 8424 39816 8430
rect 39764 8366 39816 8372
rect 39776 8022 39804 8366
rect 39764 8016 39816 8022
rect 39764 7958 39816 7964
rect 41432 7546 41460 12974
rect 42168 12850 42196 13466
rect 41512 12844 41564 12850
rect 41512 12786 41564 12792
rect 42156 12844 42208 12850
rect 42156 12786 42208 12792
rect 41524 12238 41552 12786
rect 41512 12232 41564 12238
rect 41512 12174 41564 12180
rect 41420 7540 41472 7546
rect 41420 7482 41472 7488
rect 38752 7404 38804 7410
rect 38752 7346 38804 7352
rect 39672 7404 39724 7410
rect 39672 7346 39724 7352
rect 38292 6724 38344 6730
rect 38292 6666 38344 6672
rect 37740 6452 37792 6458
rect 37740 6394 37792 6400
rect 37648 5772 37700 5778
rect 37648 5714 37700 5720
rect 38304 5642 38332 6666
rect 38764 6186 38792 7346
rect 38844 7268 38896 7274
rect 38844 7210 38896 7216
rect 38856 6798 38884 7210
rect 38844 6792 38896 6798
rect 38844 6734 38896 6740
rect 41972 6316 42024 6322
rect 41972 6258 42024 6264
rect 38752 6180 38804 6186
rect 38752 6122 38804 6128
rect 41984 5914 42012 6258
rect 41972 5908 42024 5914
rect 41972 5850 42024 5856
rect 38292 5636 38344 5642
rect 38292 5578 38344 5584
rect 42064 5636 42116 5642
rect 42064 5578 42116 5584
rect 42076 5545 42104 5578
rect 42062 5536 42118 5545
rect 42062 5471 42118 5480
rect 37464 5160 37516 5166
rect 37464 5102 37516 5108
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 33048 4548 33100 4554
rect 33048 4490 33100 4496
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 11440 2746 11560 2774
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 11440 2446 11468 2746
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 11624 800 11652 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 11610 0 11666 800
<< via2 >>
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 35600 43546 35656 43548
rect 35680 43546 35736 43548
rect 35760 43546 35816 43548
rect 35840 43546 35896 43548
rect 35600 43494 35646 43546
rect 35646 43494 35656 43546
rect 35680 43494 35710 43546
rect 35710 43494 35722 43546
rect 35722 43494 35736 43546
rect 35760 43494 35774 43546
rect 35774 43494 35786 43546
rect 35786 43494 35816 43546
rect 35840 43494 35850 43546
rect 35850 43494 35896 43546
rect 35600 43492 35656 43494
rect 35680 43492 35736 43494
rect 35760 43492 35816 43494
rect 35840 43492 35896 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 110 41928 166 41984
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 3146 32952 3202 33008
rect 2410 31356 2412 31376
rect 2412 31356 2464 31376
rect 2464 31356 2466 31376
rect 2410 31320 2466 31356
rect 2778 31320 2834 31376
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 846 27820 848 27840
rect 848 27820 900 27840
rect 900 27820 902 27840
rect 846 27784 902 27820
rect 5446 32952 5502 33008
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 5262 30252 5318 30288
rect 5262 30232 5264 30252
rect 5264 30232 5316 30252
rect 5316 30232 5318 30252
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 846 26036 902 26072
rect 846 26016 848 26036
rect 848 26016 900 26036
rect 900 26016 902 26036
rect 1306 25200 1362 25256
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4526 27396 4582 27432
rect 4526 27376 4528 27396
rect 4528 27376 4580 27396
rect 4580 27376 4582 27396
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4710 26580 4766 26616
rect 4710 26560 4712 26580
rect 4712 26560 4764 26580
rect 4764 26560 4766 26580
rect 4710 26288 4766 26344
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 5078 26324 5080 26344
rect 5080 26324 5132 26344
rect 5132 26324 5134 26344
rect 5078 26288 5134 26324
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 5906 31356 5908 31376
rect 5908 31356 5960 31376
rect 5960 31356 5962 31376
rect 5906 31320 5962 31356
rect 5722 27396 5778 27432
rect 5722 27376 5724 27396
rect 5724 27376 5776 27396
rect 5776 27376 5778 27396
rect 5354 26424 5410 26480
rect 7654 30232 7710 30288
rect 5998 26560 6054 26616
rect 5814 26424 5870 26480
rect 6182 26324 6184 26344
rect 6184 26324 6236 26344
rect 6236 26324 6238 26344
rect 6182 26288 6238 26324
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 1582 23160 1638 23216
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 1306 22480 1362 22536
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 1398 17720 1454 17776
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 846 17196 902 17232
rect 846 17176 848 17196
rect 848 17176 900 17196
rect 900 17176 902 17196
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 6090 24148 6092 24168
rect 6092 24148 6144 24168
rect 6144 24148 6146 24168
rect 6090 24112 6146 24148
rect 5998 21936 6054 21992
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 846 15816 902 15872
rect 1398 15000 1454 15056
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4894 17196 4950 17232
rect 4894 17176 4896 17196
rect 4896 17176 4948 17196
rect 4948 17176 4950 17196
rect 4986 16904 5042 16960
rect 5538 17176 5594 17232
rect 5354 17040 5410 17096
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 1490 12960 1546 13016
rect 1214 12280 1270 12336
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 3330 11600 3386 11656
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 7010 24248 7066 24304
rect 7654 24112 7710 24168
rect 11978 26288 12034 26344
rect 12898 28484 12954 28520
rect 12898 28464 12900 28484
rect 12900 28464 12952 28484
rect 12952 28464 12954 28484
rect 7470 21972 7472 21992
rect 7472 21972 7524 21992
rect 7524 21972 7526 21992
rect 7470 21936 7526 21972
rect 9218 24248 9274 24304
rect 6734 17040 6790 17096
rect 6458 16904 6514 16960
rect 12714 24812 12770 24848
rect 12714 24792 12716 24812
rect 12716 24792 12768 24812
rect 12768 24792 12770 24812
rect 13450 25236 13452 25256
rect 13452 25236 13504 25256
rect 13504 25236 13506 25256
rect 13450 25200 13506 25236
rect 14370 27376 14426 27432
rect 16854 32444 16856 32464
rect 16856 32444 16908 32464
rect 16908 32444 16910 32464
rect 16854 32408 16910 32444
rect 15014 26968 15070 27024
rect 14462 26152 14518 26208
rect 14738 26036 14794 26072
rect 14738 26016 14740 26036
rect 14740 26016 14792 26036
rect 14792 26016 14794 26036
rect 16118 27512 16174 27568
rect 15474 26444 15530 26480
rect 15474 26424 15476 26444
rect 15476 26424 15528 26444
rect 15528 26424 15530 26444
rect 15750 26016 15806 26072
rect 5906 12180 5908 12200
rect 5908 12180 5960 12200
rect 5960 12180 5962 12200
rect 5906 12144 5962 12180
rect 6642 12164 6698 12200
rect 6642 12144 6644 12164
rect 6644 12144 6696 12164
rect 6696 12144 6698 12164
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 16302 27124 16358 27160
rect 16302 27104 16304 27124
rect 16304 27104 16356 27124
rect 16356 27104 16358 27124
rect 16394 26444 16450 26480
rect 16394 26424 16396 26444
rect 16396 26424 16448 26444
rect 16448 26424 16450 26444
rect 18786 37168 18842 37224
rect 19338 36644 19394 36680
rect 19338 36624 19340 36644
rect 19340 36624 19392 36644
rect 19392 36624 19394 36644
rect 18786 36488 18842 36544
rect 17406 31084 17408 31104
rect 17408 31084 17460 31104
rect 17460 31084 17462 31104
rect 17406 31048 17462 31084
rect 16946 26868 16948 26888
rect 16948 26868 17000 26888
rect 17000 26868 17002 26888
rect 16946 26832 17002 26868
rect 16946 25200 17002 25256
rect 18050 29688 18106 29744
rect 17774 29452 17776 29472
rect 17776 29452 17828 29472
rect 17828 29452 17830 29472
rect 17774 29416 17830 29452
rect 17682 27648 17738 27704
rect 17314 27104 17370 27160
rect 17222 26968 17278 27024
rect 17498 26852 17554 26888
rect 17498 26832 17500 26852
rect 17500 26832 17552 26852
rect 17552 26832 17554 26852
rect 17866 27104 17922 27160
rect 17222 26324 17224 26344
rect 17224 26324 17276 26344
rect 17276 26324 17278 26344
rect 17222 26288 17278 26324
rect 16670 24792 16726 24848
rect 17130 23704 17186 23760
rect 17866 23840 17922 23896
rect 18694 30116 18750 30152
rect 18694 30096 18696 30116
rect 18696 30096 18748 30116
rect 18748 30096 18750 30116
rect 18694 28328 18750 28384
rect 18418 26152 18474 26208
rect 18418 24520 18474 24576
rect 17590 23432 17646 23488
rect 16026 21004 16082 21040
rect 16026 20984 16028 21004
rect 16028 20984 16080 21004
rect 16080 20984 16082 21004
rect 18510 24148 18512 24168
rect 18512 24148 18564 24168
rect 18564 24148 18566 24168
rect 18510 24112 18566 24148
rect 19890 36624 19946 36680
rect 20166 36524 20168 36544
rect 20168 36524 20220 36544
rect 20220 36524 20222 36544
rect 20166 36488 20222 36524
rect 19062 26832 19118 26888
rect 19154 26152 19210 26208
rect 19706 30812 19708 30832
rect 19708 30812 19760 30832
rect 19760 30812 19762 30832
rect 19706 30776 19762 30812
rect 19982 30796 20038 30832
rect 19982 30776 19984 30796
rect 19984 30776 20036 30796
rect 20036 30776 20038 30796
rect 19522 29416 19578 29472
rect 19430 28328 19486 28384
rect 19522 24384 19578 24440
rect 19430 24148 19432 24168
rect 19432 24148 19484 24168
rect 19484 24148 19486 24168
rect 19430 24112 19486 24148
rect 17130 16108 17186 16144
rect 17130 16088 17132 16108
rect 17132 16088 17184 16108
rect 17184 16088 17186 16108
rect 18050 15136 18106 15192
rect 20258 27512 20314 27568
rect 20258 26852 20314 26888
rect 20258 26832 20260 26852
rect 20260 26832 20312 26852
rect 20312 26832 20314 26852
rect 19706 18536 19762 18592
rect 22190 38256 22246 38312
rect 22098 34176 22154 34232
rect 20718 29588 20720 29608
rect 20720 29588 20772 29608
rect 20772 29588 20774 29608
rect 20718 29552 20774 29588
rect 20994 29164 21050 29200
rect 20994 29144 20996 29164
rect 20996 29144 21048 29164
rect 21048 29144 21050 29164
rect 20810 27376 20866 27432
rect 21638 29824 21694 29880
rect 21178 26868 21180 26888
rect 21180 26868 21232 26888
rect 21232 26868 21234 26888
rect 21178 26832 21234 26868
rect 22190 29824 22246 29880
rect 23018 38276 23074 38312
rect 23018 38256 23020 38276
rect 23020 38256 23072 38276
rect 23072 38256 23074 38276
rect 22374 30540 22376 30560
rect 22376 30540 22428 30560
rect 22428 30540 22430 30560
rect 22374 30504 22430 30540
rect 22098 29164 22154 29200
rect 22098 29144 22100 29164
rect 22100 29144 22152 29164
rect 22152 29144 22154 29164
rect 22466 29844 22522 29880
rect 22466 29824 22468 29844
rect 22468 29824 22520 29844
rect 22520 29824 22522 29844
rect 20442 23860 20498 23896
rect 20442 23840 20444 23860
rect 20444 23840 20496 23860
rect 20496 23840 20498 23860
rect 22374 27668 22430 27704
rect 22374 27648 22376 27668
rect 22376 27648 22428 27668
rect 22428 27648 22430 27668
rect 22098 25100 22100 25120
rect 22100 25100 22152 25120
rect 22152 25100 22154 25120
rect 22098 25064 22154 25100
rect 22466 24792 22522 24848
rect 21822 15544 21878 15600
rect 22742 28464 22798 28520
rect 22834 27240 22890 27296
rect 23386 40976 23442 41032
rect 23202 29280 23258 29336
rect 23478 29416 23534 29472
rect 23018 27532 23074 27568
rect 23018 27512 23020 27532
rect 23020 27512 23072 27532
rect 23072 27512 23074 27532
rect 23938 29416 23994 29472
rect 23754 26968 23810 27024
rect 23570 25064 23626 25120
rect 22466 15580 22468 15600
rect 22468 15580 22520 15600
rect 22520 15580 22522 15600
rect 22466 15544 22522 15580
rect 24214 31220 24216 31240
rect 24216 31220 24268 31240
rect 24268 31220 24270 31240
rect 24214 31184 24270 31220
rect 24490 29416 24546 29472
rect 24950 29416 25006 29472
rect 25318 27648 25374 27704
rect 25686 29280 25742 29336
rect 26146 29416 26202 29472
rect 26238 29144 26294 29200
rect 25226 24384 25282 24440
rect 25594 24656 25650 24712
rect 26514 28364 26516 28384
rect 26516 28364 26568 28384
rect 26568 28364 26570 28384
rect 26514 28328 26570 28364
rect 26514 26988 26570 27024
rect 27526 38256 27582 38312
rect 27802 40840 27858 40896
rect 28078 40468 28080 40488
rect 28080 40468 28132 40488
rect 28132 40468 28134 40488
rect 27802 40296 27858 40352
rect 28078 40432 28134 40468
rect 26790 28464 26846 28520
rect 26514 26968 26516 26988
rect 26516 26968 26568 26988
rect 26568 26968 26570 26988
rect 26882 27648 26938 27704
rect 26514 24384 26570 24440
rect 25594 15136 25650 15192
rect 28630 40876 28632 40896
rect 28632 40876 28684 40896
rect 28684 40876 28686 40896
rect 28630 40840 28686 40876
rect 28446 40296 28502 40352
rect 28906 40468 28908 40488
rect 28908 40468 28960 40488
rect 28960 40468 28962 40488
rect 28906 40432 28962 40468
rect 28906 40332 28908 40352
rect 28908 40332 28960 40352
rect 28960 40332 28962 40352
rect 28906 40296 28962 40332
rect 29090 36216 29146 36272
rect 30930 40976 30986 41032
rect 30930 40024 30986 40080
rect 28170 28600 28226 28656
rect 28630 29180 28632 29200
rect 28632 29180 28684 29200
rect 28684 29180 28686 29200
rect 28630 29144 28686 29180
rect 28906 27920 28962 27976
rect 28998 27104 29054 27160
rect 31482 36796 31484 36816
rect 31484 36796 31536 36816
rect 31536 36796 31538 36816
rect 31482 36760 31538 36796
rect 31758 40024 31814 40080
rect 31758 36080 31814 36136
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 35600 42458 35656 42460
rect 35680 42458 35736 42460
rect 35760 42458 35816 42460
rect 35840 42458 35896 42460
rect 35600 42406 35646 42458
rect 35646 42406 35656 42458
rect 35680 42406 35710 42458
rect 35710 42406 35722 42458
rect 35722 42406 35736 42458
rect 35760 42406 35774 42458
rect 35774 42406 35786 42458
rect 35786 42406 35816 42458
rect 35840 42406 35850 42458
rect 35850 42406 35896 42458
rect 35600 42404 35656 42406
rect 35680 42404 35736 42406
rect 35760 42404 35816 42406
rect 35840 42404 35896 42406
rect 35600 41370 35656 41372
rect 35680 41370 35736 41372
rect 35760 41370 35816 41372
rect 35840 41370 35896 41372
rect 35600 41318 35646 41370
rect 35646 41318 35656 41370
rect 35680 41318 35710 41370
rect 35710 41318 35722 41370
rect 35722 41318 35736 41370
rect 35760 41318 35774 41370
rect 35774 41318 35786 41370
rect 35786 41318 35816 41370
rect 35840 41318 35850 41370
rect 35850 41318 35896 41370
rect 35600 41316 35656 41318
rect 35680 41316 35736 41318
rect 35760 41316 35816 41318
rect 35840 41316 35896 41318
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 27986 24520 28042 24576
rect 26238 15136 26294 15192
rect 27250 15272 27306 15328
rect 30470 29280 30526 29336
rect 30102 27376 30158 27432
rect 30010 24112 30066 24168
rect 30562 28736 30618 28792
rect 30378 27920 30434 27976
rect 30562 27648 30618 27704
rect 30930 27648 30986 27704
rect 33874 38528 33930 38584
rect 32218 29008 32274 29064
rect 31942 26288 31998 26344
rect 31298 23740 31300 23760
rect 31300 23740 31352 23760
rect 31352 23740 31354 23760
rect 31298 23704 31354 23740
rect 28078 12844 28134 12880
rect 28078 12824 28080 12844
rect 28080 12824 28132 12844
rect 28132 12824 28134 12844
rect 27342 10920 27398 10976
rect 29550 12824 29606 12880
rect 30286 6296 30342 6352
rect 33966 37188 34022 37224
rect 33966 37168 33968 37188
rect 33968 37168 34020 37188
rect 34020 37168 34022 37188
rect 32954 29144 33010 29200
rect 32770 28736 32826 28792
rect 33138 28056 33194 28112
rect 33322 29008 33378 29064
rect 33598 29688 33654 29744
rect 33598 29416 33654 29472
rect 35600 40282 35656 40284
rect 35680 40282 35736 40284
rect 35760 40282 35816 40284
rect 35840 40282 35896 40284
rect 35600 40230 35646 40282
rect 35646 40230 35656 40282
rect 35680 40230 35710 40282
rect 35710 40230 35722 40282
rect 35722 40230 35736 40282
rect 35760 40230 35774 40282
rect 35774 40230 35786 40282
rect 35786 40230 35816 40282
rect 35840 40230 35850 40282
rect 35850 40230 35896 40282
rect 35600 40228 35656 40230
rect 35680 40228 35736 40230
rect 35760 40228 35816 40230
rect 35840 40228 35896 40230
rect 35162 38800 35218 38856
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 35714 38820 35770 38856
rect 35714 38800 35716 38820
rect 35716 38800 35768 38820
rect 35768 38800 35770 38820
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 37462 36760 37518 36816
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34242 30096 34298 30152
rect 33874 29572 33930 29608
rect 33874 29552 33876 29572
rect 33876 29552 33928 29572
rect 33928 29552 33930 29572
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34610 30368 34666 30424
rect 34242 28872 34298 28928
rect 33966 27648 34022 27704
rect 33782 27512 33838 27568
rect 34058 27512 34114 27568
rect 31942 17040 31998 17096
rect 31850 11872 31906 11928
rect 32494 12008 32550 12064
rect 34610 29280 34666 29336
rect 35714 30640 35770 30696
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34794 29416 34850 29472
rect 35438 30096 35494 30152
rect 35254 29416 35310 29472
rect 34978 29280 35034 29336
rect 35346 29008 35402 29064
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34242 27240 34298 27296
rect 34150 26832 34206 26888
rect 33966 26424 34022 26480
rect 34610 27104 34666 27160
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 33506 21836 33508 21856
rect 33508 21836 33560 21856
rect 33560 21836 33562 21856
rect 33506 21800 33562 21836
rect 35162 25200 35218 25256
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 35806 29028 35862 29064
rect 35806 29008 35808 29028
rect 35808 29008 35860 29028
rect 35860 29008 35862 29028
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 36174 29688 36230 29744
rect 36174 29452 36176 29472
rect 36176 29452 36228 29472
rect 36228 29452 36230 29472
rect 36174 29416 36230 29452
rect 36082 28056 36138 28112
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 35530 26696 35586 26752
rect 35622 26560 35678 26616
rect 36634 30096 36690 30152
rect 36358 26988 36414 27024
rect 36634 29416 36690 29472
rect 36910 29552 36966 29608
rect 36358 26968 36360 26988
rect 36360 26968 36412 26988
rect 36412 26968 36414 26988
rect 36542 26560 36598 26616
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 35898 25220 35954 25256
rect 35898 25200 35900 25220
rect 35900 25200 35952 25220
rect 35952 25200 35954 25220
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35530 23180 35586 23216
rect 35530 23160 35532 23180
rect 35532 23160 35584 23180
rect 35584 23160 35586 23180
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 33782 21292 33784 21312
rect 33784 21292 33836 21312
rect 33836 21292 33838 21312
rect 33782 21256 33838 21292
rect 32954 12180 32956 12200
rect 32956 12180 33008 12200
rect 33008 12180 33010 12200
rect 32954 12144 33010 12180
rect 33690 12300 33746 12336
rect 33690 12280 33692 12300
rect 33692 12280 33744 12300
rect 33744 12280 33746 12300
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 36450 23160 36506 23216
rect 37094 29144 37150 29200
rect 37646 28600 37702 28656
rect 38658 36216 38714 36272
rect 37278 27548 37280 27568
rect 37280 27548 37332 27568
rect 37332 27548 37334 27568
rect 37278 27512 37334 27548
rect 37002 26696 37058 26752
rect 37186 26308 37242 26344
rect 37186 26288 37188 26308
rect 37188 26288 37240 26308
rect 37240 26288 37242 26308
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 35714 12144 35770 12200
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 32586 6316 32642 6352
rect 32586 6296 32588 6316
rect 32588 6296 32640 6316
rect 32640 6296 32642 6316
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 39210 36100 39266 36136
rect 39210 36080 39212 36100
rect 39212 36080 39264 36100
rect 39264 36080 39266 36100
rect 38474 28464 38530 28520
rect 40498 33224 40554 33280
rect 39026 27648 39082 27704
rect 39302 27412 39304 27432
rect 39304 27412 39356 27432
rect 39356 27412 39358 27432
rect 39302 27376 39358 27412
rect 39026 25880 39082 25936
rect 39486 24132 39542 24168
rect 39486 24112 39488 24132
rect 39488 24112 39540 24132
rect 39540 24112 39542 24132
rect 39394 23160 39450 23216
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 38934 12164 38990 12200
rect 38934 12144 38936 12164
rect 38936 12144 38988 12164
rect 38988 12144 38990 12164
rect 40038 27124 40094 27160
rect 40038 27104 40040 27124
rect 40040 27104 40092 27124
rect 40092 27104 40094 27124
rect 40038 23704 40094 23760
rect 40222 23840 40278 23896
rect 40130 23160 40186 23216
rect 41970 29996 41972 30016
rect 41972 29996 42024 30016
rect 42024 29996 42026 30016
rect 41970 29960 42026 29996
rect 41694 27940 41750 27976
rect 41694 27920 41696 27940
rect 41696 27920 41748 27940
rect 41748 27920 41750 27940
rect 40774 26832 40830 26888
rect 40958 24812 41014 24848
rect 40958 24792 40960 24812
rect 40960 24792 41012 24812
rect 41012 24792 41014 24812
rect 40866 24656 40922 24712
rect 41142 23724 41198 23760
rect 41142 23704 41144 23724
rect 41144 23704 41196 23724
rect 41196 23704 41198 23724
rect 41878 25900 41934 25936
rect 41878 25880 41880 25900
rect 41880 25880 41932 25900
rect 41932 25880 41934 25900
rect 41510 25200 41566 25256
rect 42062 29280 42118 29336
rect 42062 28600 42118 28656
rect 42062 27240 42118 27296
rect 42062 26560 42118 26616
rect 42062 25880 42118 25936
rect 41510 24556 41512 24576
rect 41512 24556 41564 24576
rect 41564 24556 41566 24576
rect 41510 24520 41566 24556
rect 41602 23160 41658 23216
rect 42154 23160 42210 23216
rect 39762 12164 39818 12200
rect 39762 12144 39764 12164
rect 39764 12144 39816 12164
rect 39816 12144 39818 12164
rect 42062 5480 42118 5536
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 35590 43552 35906 43553
rect 35590 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35906 43552
rect 35590 43487 35906 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 35590 42464 35906 42465
rect 35590 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35906 42464
rect 35590 42399 35906 42400
rect 0 42258 800 42288
rect 0 42198 1042 42258
rect 0 42168 800 42198
rect 105 41986 171 41989
rect 982 41986 1042 42198
rect 105 41984 1042 41986
rect 105 41928 110 41984
rect 166 41928 1042 41984
rect 105 41926 1042 41928
rect 105 41923 171 41926
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 35590 41376 35906 41377
rect 35590 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35906 41376
rect 35590 41311 35906 41312
rect 23381 41034 23447 41037
rect 30925 41034 30991 41037
rect 23381 41032 30991 41034
rect 23381 40976 23386 41032
rect 23442 40976 30930 41032
rect 30986 40976 30991 41032
rect 23381 40974 30991 40976
rect 23381 40971 23447 40974
rect 30925 40971 30991 40974
rect 27797 40898 27863 40901
rect 28625 40898 28691 40901
rect 27797 40896 28691 40898
rect 27797 40840 27802 40896
rect 27858 40840 28630 40896
rect 28686 40840 28691 40896
rect 27797 40838 28691 40840
rect 27797 40835 27863 40838
rect 28625 40835 28691 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 28073 40490 28139 40493
rect 28901 40490 28967 40493
rect 28073 40488 28967 40490
rect 28073 40432 28078 40488
rect 28134 40432 28906 40488
rect 28962 40432 28967 40488
rect 28073 40430 28967 40432
rect 28073 40427 28139 40430
rect 28901 40427 28967 40430
rect 27797 40354 27863 40357
rect 28441 40354 28507 40357
rect 28901 40354 28967 40357
rect 27797 40352 28967 40354
rect 27797 40296 27802 40352
rect 27858 40296 28446 40352
rect 28502 40296 28906 40352
rect 28962 40296 28967 40352
rect 27797 40294 28967 40296
rect 27797 40291 27863 40294
rect 28441 40291 28507 40294
rect 28901 40291 28967 40294
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 35590 40288 35906 40289
rect 35590 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35906 40288
rect 35590 40223 35906 40224
rect 30925 40082 30991 40085
rect 31753 40082 31819 40085
rect 30925 40080 31819 40082
rect 30925 40024 30930 40080
rect 30986 40024 31758 40080
rect 31814 40024 31819 40080
rect 30925 40022 31819 40024
rect 30925 40019 30991 40022
rect 31753 40019 31819 40022
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 34646 38796 34652 38860
rect 34716 38858 34722 38860
rect 35157 38858 35223 38861
rect 35709 38858 35775 38861
rect 34716 38856 35775 38858
rect 34716 38800 35162 38856
rect 35218 38800 35714 38856
rect 35770 38800 35775 38856
rect 34716 38798 35775 38800
rect 34716 38796 34722 38798
rect 35157 38795 35223 38798
rect 35709 38795 35775 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 33869 38588 33935 38589
rect 33869 38586 33916 38588
rect 33824 38584 33916 38586
rect 33824 38528 33874 38584
rect 33824 38526 33916 38528
rect 33869 38524 33916 38526
rect 33980 38524 33986 38588
rect 33869 38523 33935 38524
rect 22185 38314 22251 38317
rect 23013 38314 23079 38317
rect 27521 38314 27587 38317
rect 22185 38312 27587 38314
rect 22185 38256 22190 38312
rect 22246 38256 23018 38312
rect 23074 38256 27526 38312
rect 27582 38256 27587 38312
rect 22185 38254 27587 38256
rect 22185 38251 22251 38254
rect 23013 38251 23079 38254
rect 27521 38251 27587 38254
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 18781 37226 18847 37229
rect 33961 37226 34027 37229
rect 18781 37224 34027 37226
rect 18781 37168 18786 37224
rect 18842 37168 33966 37224
rect 34022 37168 34027 37224
rect 18781 37166 34027 37168
rect 18781 37163 18847 37166
rect 33961 37163 34027 37166
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 31477 36818 31543 36821
rect 37457 36818 37523 36821
rect 31477 36816 37523 36818
rect 31477 36760 31482 36816
rect 31538 36760 37462 36816
rect 37518 36760 37523 36816
rect 31477 36758 37523 36760
rect 31477 36755 31543 36758
rect 37457 36755 37523 36758
rect 19333 36682 19399 36685
rect 19885 36682 19951 36685
rect 19333 36680 19951 36682
rect 19333 36624 19338 36680
rect 19394 36624 19890 36680
rect 19946 36624 19951 36680
rect 19333 36622 19951 36624
rect 19333 36619 19399 36622
rect 19885 36619 19951 36622
rect 18781 36546 18847 36549
rect 20161 36546 20227 36549
rect 18781 36544 20227 36546
rect 18781 36488 18786 36544
rect 18842 36488 20166 36544
rect 20222 36488 20227 36544
rect 18781 36486 20227 36488
rect 18781 36483 18847 36486
rect 20161 36483 20227 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 29085 36274 29151 36277
rect 38653 36274 38719 36277
rect 29085 36272 38719 36274
rect 29085 36216 29090 36272
rect 29146 36216 38658 36272
rect 38714 36216 38719 36272
rect 29085 36214 38719 36216
rect 29085 36211 29151 36214
rect 38653 36211 38719 36214
rect 31753 36138 31819 36141
rect 39205 36138 39271 36141
rect 31753 36136 39271 36138
rect 31753 36080 31758 36136
rect 31814 36080 39210 36136
rect 39266 36080 39271 36136
rect 31753 36078 39271 36080
rect 31753 36075 31819 36078
rect 39205 36075 39271 36078
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 22093 34236 22159 34237
rect 22093 34232 22140 34236
rect 22204 34234 22210 34236
rect 22093 34176 22098 34232
rect 22093 34172 22140 34176
rect 22204 34174 22250 34234
rect 22204 34172 22210 34174
rect 22093 34171 22159 34172
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 40166 33220 40172 33284
rect 40236 33282 40242 33284
rect 40493 33282 40559 33285
rect 40236 33280 40559 33282
rect 40236 33224 40498 33280
rect 40554 33224 40559 33280
rect 40236 33222 40559 33224
rect 40236 33220 40242 33222
rect 40493 33219 40559 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 3141 33010 3207 33013
rect 5441 33010 5507 33013
rect 3141 33008 5507 33010
rect 3141 32952 3146 33008
rect 3202 32952 5446 33008
rect 5502 32952 5507 33008
rect 3141 32950 5507 32952
rect 3141 32947 3207 32950
rect 5441 32947 5507 32950
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 16849 32466 16915 32469
rect 17718 32466 17724 32468
rect 16849 32464 17724 32466
rect 16849 32408 16854 32464
rect 16910 32408 17724 32464
rect 16849 32406 17724 32408
rect 16849 32403 16915 32406
rect 17718 32404 17724 32406
rect 17788 32404 17794 32468
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 2405 31378 2471 31381
rect 2773 31378 2839 31381
rect 5901 31378 5967 31381
rect 2405 31376 5967 31378
rect 2405 31320 2410 31376
rect 2466 31320 2778 31376
rect 2834 31320 5906 31376
rect 5962 31320 5967 31376
rect 2405 31318 5967 31320
rect 2405 31315 2471 31318
rect 2773 31315 2839 31318
rect 5901 31315 5967 31318
rect 24209 31242 24275 31245
rect 24894 31242 24900 31244
rect 24209 31240 24900 31242
rect 24209 31184 24214 31240
rect 24270 31184 24900 31240
rect 24209 31182 24900 31184
rect 24209 31179 24275 31182
rect 24894 31180 24900 31182
rect 24964 31180 24970 31244
rect 17401 31106 17467 31109
rect 17534 31106 17540 31108
rect 17401 31104 17540 31106
rect 17401 31048 17406 31104
rect 17462 31048 17540 31104
rect 17401 31046 17540 31048
rect 17401 31043 17467 31046
rect 17534 31044 17540 31046
rect 17604 31044 17610 31108
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19701 30834 19767 30837
rect 19977 30834 20043 30837
rect 19701 30832 20043 30834
rect 19701 30776 19706 30832
rect 19762 30776 19982 30832
rect 20038 30776 20043 30832
rect 19701 30774 20043 30776
rect 19701 30771 19767 30774
rect 19977 30771 20043 30774
rect 35709 30698 35775 30701
rect 36118 30698 36124 30700
rect 35709 30696 36124 30698
rect 35709 30640 35714 30696
rect 35770 30640 36124 30696
rect 35709 30638 36124 30640
rect 35709 30635 35775 30638
rect 36118 30636 36124 30638
rect 36188 30636 36194 30700
rect 22369 30564 22435 30565
rect 22318 30500 22324 30564
rect 22388 30562 22435 30564
rect 22388 30560 22480 30562
rect 22430 30504 22480 30560
rect 22388 30502 22480 30504
rect 22388 30500 22435 30502
rect 22369 30499 22435 30500
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 34462 30364 34468 30428
rect 34532 30426 34538 30428
rect 34605 30426 34671 30429
rect 34532 30424 34671 30426
rect 34532 30368 34610 30424
rect 34666 30368 34671 30424
rect 34532 30366 34671 30368
rect 34532 30364 34538 30366
rect 34605 30363 34671 30366
rect 5257 30290 5323 30293
rect 7649 30290 7715 30293
rect 5257 30288 7715 30290
rect 5257 30232 5262 30288
rect 5318 30232 7654 30288
rect 7710 30232 7715 30288
rect 5257 30230 7715 30232
rect 5257 30227 5323 30230
rect 7649 30227 7715 30230
rect 18689 30154 18755 30157
rect 34237 30154 34303 30157
rect 18689 30152 34303 30154
rect 18689 30096 18694 30152
rect 18750 30096 34242 30152
rect 34298 30096 34303 30152
rect 18689 30094 34303 30096
rect 18689 30091 18755 30094
rect 34237 30091 34303 30094
rect 35433 30154 35499 30157
rect 36629 30154 36695 30157
rect 35433 30152 36695 30154
rect 35433 30096 35438 30152
rect 35494 30096 36634 30152
rect 36690 30096 36695 30152
rect 35433 30094 36695 30096
rect 35433 30091 35499 30094
rect 36629 30091 36695 30094
rect 41965 30018 42031 30021
rect 42813 30018 43613 30048
rect 41965 30016 43613 30018
rect 41965 29960 41970 30016
rect 42026 29960 43613 30016
rect 41965 29958 43613 29960
rect 41965 29955 42031 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 42813 29928 43613 29958
rect 34930 29887 35246 29888
rect 21633 29882 21699 29885
rect 22185 29882 22251 29885
rect 22461 29882 22527 29885
rect 21633 29880 22527 29882
rect 21633 29824 21638 29880
rect 21694 29824 22190 29880
rect 22246 29824 22466 29880
rect 22522 29824 22527 29880
rect 21633 29822 22527 29824
rect 21633 29819 21699 29822
rect 22185 29819 22251 29822
rect 22461 29819 22527 29822
rect 18045 29746 18111 29749
rect 33593 29746 33659 29749
rect 36169 29746 36235 29749
rect 18045 29744 36235 29746
rect 18045 29688 18050 29744
rect 18106 29688 33598 29744
rect 33654 29688 36174 29744
rect 36230 29688 36235 29744
rect 18045 29686 36235 29688
rect 18045 29683 18111 29686
rect 33593 29683 33659 29686
rect 36169 29683 36235 29686
rect 20713 29610 20779 29613
rect 33869 29610 33935 29613
rect 36905 29610 36971 29613
rect 20713 29608 33935 29610
rect 20713 29552 20718 29608
rect 20774 29552 33874 29608
rect 33930 29552 33935 29608
rect 20713 29550 33935 29552
rect 20713 29547 20779 29550
rect 33869 29547 33935 29550
rect 34102 29608 36971 29610
rect 34102 29552 36910 29608
rect 36966 29552 36971 29608
rect 34102 29550 36971 29552
rect 17166 29412 17172 29476
rect 17236 29474 17242 29476
rect 17769 29474 17835 29477
rect 19517 29474 19583 29477
rect 17236 29472 19583 29474
rect 17236 29416 17774 29472
rect 17830 29416 19522 29472
rect 19578 29416 19583 29472
rect 17236 29414 19583 29416
rect 17236 29412 17242 29414
rect 17769 29411 17835 29414
rect 19517 29411 19583 29414
rect 23473 29474 23539 29477
rect 23933 29474 23999 29477
rect 23473 29472 23999 29474
rect 23473 29416 23478 29472
rect 23534 29416 23938 29472
rect 23994 29416 23999 29472
rect 23473 29414 23999 29416
rect 23473 29411 23539 29414
rect 23933 29411 23999 29414
rect 24485 29474 24551 29477
rect 24945 29474 25011 29477
rect 26141 29474 26207 29477
rect 24485 29472 26207 29474
rect 24485 29416 24490 29472
rect 24546 29416 24950 29472
rect 25006 29416 26146 29472
rect 26202 29416 26207 29472
rect 24485 29414 26207 29416
rect 24485 29411 24551 29414
rect 24945 29411 25011 29414
rect 26141 29411 26207 29414
rect 33593 29474 33659 29477
rect 34102 29474 34162 29550
rect 36905 29547 36971 29550
rect 33593 29472 34162 29474
rect 33593 29416 33598 29472
rect 33654 29416 34162 29472
rect 33593 29414 34162 29416
rect 34789 29474 34855 29477
rect 35249 29474 35315 29477
rect 34789 29472 35315 29474
rect 34789 29416 34794 29472
rect 34850 29416 35254 29472
rect 35310 29416 35315 29472
rect 34789 29414 35315 29416
rect 33593 29411 33659 29414
rect 34789 29411 34855 29414
rect 35249 29411 35315 29414
rect 36169 29474 36235 29477
rect 36629 29474 36695 29477
rect 36169 29472 36695 29474
rect 36169 29416 36174 29472
rect 36230 29416 36634 29472
rect 36690 29416 36695 29472
rect 36169 29414 36695 29416
rect 36169 29411 36235 29414
rect 36629 29411 36695 29414
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 23197 29338 23263 29341
rect 25681 29338 25747 29341
rect 23197 29336 25747 29338
rect 23197 29280 23202 29336
rect 23258 29280 25686 29336
rect 25742 29280 25747 29336
rect 23197 29278 25747 29280
rect 23197 29275 23263 29278
rect 25681 29275 25747 29278
rect 30465 29338 30531 29341
rect 34605 29338 34671 29341
rect 34973 29338 35039 29341
rect 30465 29336 35039 29338
rect 30465 29280 30470 29336
rect 30526 29280 34610 29336
rect 34666 29280 34978 29336
rect 35034 29280 35039 29336
rect 30465 29278 35039 29280
rect 30465 29275 30531 29278
rect 34605 29275 34671 29278
rect 34973 29275 35039 29278
rect 42057 29338 42123 29341
rect 42813 29338 43613 29368
rect 42057 29336 43613 29338
rect 42057 29280 42062 29336
rect 42118 29280 43613 29336
rect 42057 29278 43613 29280
rect 42057 29275 42123 29278
rect 42813 29248 43613 29278
rect 20989 29202 21055 29205
rect 22093 29202 22159 29205
rect 20989 29200 22159 29202
rect 20989 29144 20994 29200
rect 21050 29144 22098 29200
rect 22154 29144 22159 29200
rect 20989 29142 22159 29144
rect 20989 29139 21055 29142
rect 22093 29139 22159 29142
rect 26233 29202 26299 29205
rect 28625 29202 28691 29205
rect 26233 29200 28691 29202
rect 26233 29144 26238 29200
rect 26294 29144 28630 29200
rect 28686 29144 28691 29200
rect 26233 29142 28691 29144
rect 26233 29139 26299 29142
rect 28625 29139 28691 29142
rect 32949 29202 33015 29205
rect 37089 29202 37155 29205
rect 32949 29200 37155 29202
rect 32949 29144 32954 29200
rect 33010 29144 37094 29200
rect 37150 29144 37155 29200
rect 32949 29142 37155 29144
rect 32949 29139 33015 29142
rect 37089 29139 37155 29142
rect 32213 29066 32279 29069
rect 33317 29066 33383 29069
rect 35341 29066 35407 29069
rect 32213 29064 33383 29066
rect 32213 29008 32218 29064
rect 32274 29008 33322 29064
rect 33378 29008 33383 29064
rect 32213 29006 33383 29008
rect 32213 29003 32279 29006
rect 33317 29003 33383 29006
rect 34700 29064 35407 29066
rect 34700 29008 35346 29064
rect 35402 29008 35407 29064
rect 34700 29006 35407 29008
rect 34237 28930 34303 28933
rect 34700 28930 34760 29006
rect 35341 29003 35407 29006
rect 35801 29066 35867 29069
rect 36118 29066 36124 29068
rect 35801 29064 36124 29066
rect 35801 29008 35806 29064
rect 35862 29008 36124 29064
rect 35801 29006 36124 29008
rect 35801 29003 35867 29006
rect 36118 29004 36124 29006
rect 36188 29004 36194 29068
rect 34237 28928 34760 28930
rect 34237 28872 34242 28928
rect 34298 28872 34760 28928
rect 34237 28870 34760 28872
rect 34237 28867 34303 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 30557 28794 30623 28797
rect 32765 28794 32831 28797
rect 30557 28792 32831 28794
rect 30557 28736 30562 28792
rect 30618 28736 32770 28792
rect 32826 28736 32831 28792
rect 30557 28734 32831 28736
rect 30557 28731 30623 28734
rect 32765 28731 32831 28734
rect 28165 28658 28231 28661
rect 37641 28658 37707 28661
rect 28165 28656 37707 28658
rect 28165 28600 28170 28656
rect 28226 28600 37646 28656
rect 37702 28600 37707 28656
rect 28165 28598 37707 28600
rect 28165 28595 28231 28598
rect 37641 28595 37707 28598
rect 42057 28658 42123 28661
rect 42813 28658 43613 28688
rect 42057 28656 43613 28658
rect 42057 28600 42062 28656
rect 42118 28600 43613 28656
rect 42057 28598 43613 28600
rect 42057 28595 42123 28598
rect 42813 28568 43613 28598
rect 12893 28522 12959 28525
rect 22134 28522 22140 28524
rect 12893 28520 22140 28522
rect 12893 28464 12898 28520
rect 12954 28464 22140 28520
rect 12893 28462 22140 28464
rect 12893 28459 12959 28462
rect 22134 28460 22140 28462
rect 22204 28522 22210 28524
rect 22737 28522 22803 28525
rect 22204 28520 22803 28522
rect 22204 28464 22742 28520
rect 22798 28464 22803 28520
rect 22204 28462 22803 28464
rect 22204 28460 22210 28462
rect 22737 28459 22803 28462
rect 26785 28522 26851 28525
rect 38469 28522 38535 28525
rect 26785 28520 38535 28522
rect 26785 28464 26790 28520
rect 26846 28464 38474 28520
rect 38530 28464 38535 28520
rect 26785 28462 38535 28464
rect 26785 28459 26851 28462
rect 38469 28459 38535 28462
rect 18689 28386 18755 28389
rect 19425 28386 19491 28389
rect 26509 28386 26575 28389
rect 18689 28384 26575 28386
rect 18689 28328 18694 28384
rect 18750 28328 19430 28384
rect 19486 28328 26514 28384
rect 26570 28328 26575 28384
rect 18689 28326 26575 28328
rect 18689 28323 18755 28326
rect 19425 28323 19491 28326
rect 26509 28323 26575 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 33133 28114 33199 28117
rect 36077 28114 36143 28117
rect 33133 28112 36143 28114
rect 33133 28056 33138 28112
rect 33194 28056 36082 28112
rect 36138 28056 36143 28112
rect 33133 28054 36143 28056
rect 33133 28051 33199 28054
rect 36077 28051 36143 28054
rect 0 27978 800 28008
rect 28901 27978 28967 27981
rect 30373 27978 30439 27981
rect 0 27888 858 27978
rect 28901 27976 30439 27978
rect 28901 27920 28906 27976
rect 28962 27920 30378 27976
rect 30434 27920 30439 27976
rect 28901 27918 30439 27920
rect 28901 27915 28967 27918
rect 30373 27915 30439 27918
rect 41689 27978 41755 27981
rect 42813 27978 43613 28008
rect 41689 27976 43613 27978
rect 41689 27920 41694 27976
rect 41750 27920 43613 27976
rect 41689 27918 43613 27920
rect 41689 27915 41755 27918
rect 42813 27888 43613 27918
rect 798 27845 858 27888
rect 798 27840 907 27845
rect 798 27784 846 27840
rect 902 27784 907 27840
rect 798 27782 907 27784
rect 841 27779 907 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 17677 27706 17743 27709
rect 22369 27708 22435 27709
rect 22318 27706 22324 27708
rect 17677 27704 17786 27706
rect 17677 27648 17682 27704
rect 17738 27648 17786 27704
rect 17677 27643 17786 27648
rect 22278 27646 22324 27706
rect 22388 27704 22435 27708
rect 22430 27648 22435 27704
rect 22318 27644 22324 27646
rect 22388 27644 22435 27648
rect 24894 27644 24900 27708
rect 24964 27706 24970 27708
rect 25313 27706 25379 27709
rect 26877 27706 26943 27709
rect 24964 27704 26943 27706
rect 24964 27648 25318 27704
rect 25374 27648 26882 27704
rect 26938 27648 26943 27704
rect 24964 27646 26943 27648
rect 24964 27644 24970 27646
rect 22369 27643 22435 27644
rect 25313 27643 25379 27646
rect 26877 27643 26943 27646
rect 30557 27706 30623 27709
rect 30925 27706 30991 27709
rect 33961 27706 34027 27709
rect 30557 27704 34027 27706
rect 30557 27648 30562 27704
rect 30618 27648 30930 27704
rect 30986 27648 33966 27704
rect 34022 27648 34027 27704
rect 30557 27646 34027 27648
rect 30557 27643 30623 27646
rect 30925 27643 30991 27646
rect 33961 27643 34027 27646
rect 38694 27644 38700 27708
rect 38764 27706 38770 27708
rect 39021 27706 39087 27709
rect 38764 27704 39087 27706
rect 38764 27648 39026 27704
rect 39082 27648 39087 27704
rect 38764 27646 39087 27648
rect 38764 27644 38770 27646
rect 39021 27643 39087 27646
rect 16113 27570 16179 27573
rect 17726 27570 17786 27643
rect 20253 27570 20319 27573
rect 23013 27572 23079 27573
rect 23013 27570 23060 27572
rect 16113 27568 20319 27570
rect 16113 27512 16118 27568
rect 16174 27512 20258 27568
rect 20314 27512 20319 27568
rect 16113 27510 20319 27512
rect 22968 27568 23060 27570
rect 22968 27512 23018 27568
rect 22968 27510 23060 27512
rect 16113 27507 16179 27510
rect 20253 27507 20319 27510
rect 23013 27508 23060 27510
rect 23124 27508 23130 27572
rect 33777 27570 33843 27573
rect 33910 27570 33916 27572
rect 33777 27568 33916 27570
rect 33777 27512 33782 27568
rect 33838 27512 33916 27568
rect 33777 27510 33916 27512
rect 23013 27507 23079 27508
rect 33777 27507 33843 27510
rect 33910 27508 33916 27510
rect 33980 27508 33986 27572
rect 34053 27570 34119 27573
rect 37273 27570 37339 27573
rect 34053 27568 37339 27570
rect 34053 27512 34058 27568
rect 34114 27512 37278 27568
rect 37334 27512 37339 27568
rect 34053 27510 37339 27512
rect 34053 27507 34119 27510
rect 37273 27507 37339 27510
rect 4521 27434 4587 27437
rect 5717 27434 5783 27437
rect 4521 27432 5783 27434
rect 4521 27376 4526 27432
rect 4582 27376 5722 27432
rect 5778 27376 5783 27432
rect 4521 27374 5783 27376
rect 4521 27371 4587 27374
rect 5717 27371 5783 27374
rect 14365 27434 14431 27437
rect 20805 27434 20871 27437
rect 14365 27432 20871 27434
rect 14365 27376 14370 27432
rect 14426 27376 20810 27432
rect 20866 27376 20871 27432
rect 14365 27374 20871 27376
rect 14365 27371 14431 27374
rect 20805 27371 20871 27374
rect 30097 27434 30163 27437
rect 39297 27434 39363 27437
rect 30097 27432 39363 27434
rect 30097 27376 30102 27432
rect 30158 27376 39302 27432
rect 39358 27376 39363 27432
rect 30097 27374 39363 27376
rect 30097 27371 30163 27374
rect 39297 27371 39363 27374
rect 22829 27298 22895 27301
rect 34237 27298 34303 27301
rect 22829 27296 34303 27298
rect 22829 27240 22834 27296
rect 22890 27240 34242 27296
rect 34298 27240 34303 27296
rect 22829 27238 34303 27240
rect 22829 27235 22895 27238
rect 34237 27235 34303 27238
rect 42057 27298 42123 27301
rect 42813 27298 43613 27328
rect 42057 27296 43613 27298
rect 42057 27240 42062 27296
rect 42118 27240 43613 27296
rect 42057 27238 43613 27240
rect 42057 27235 42123 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 42813 27208 43613 27238
rect 35590 27167 35906 27168
rect 16297 27162 16363 27165
rect 17309 27162 17375 27165
rect 16297 27160 17375 27162
rect 16297 27104 16302 27160
rect 16358 27104 17314 27160
rect 17370 27104 17375 27160
rect 16297 27102 17375 27104
rect 16297 27099 16363 27102
rect 17309 27099 17375 27102
rect 17861 27162 17927 27165
rect 28993 27162 29059 27165
rect 17861 27160 29059 27162
rect 17861 27104 17866 27160
rect 17922 27104 28998 27160
rect 29054 27104 29059 27160
rect 17861 27102 29059 27104
rect 17861 27099 17927 27102
rect 28993 27099 29059 27102
rect 34462 27100 34468 27164
rect 34532 27162 34538 27164
rect 34605 27162 34671 27165
rect 34532 27160 34671 27162
rect 34532 27104 34610 27160
rect 34666 27104 34671 27160
rect 34532 27102 34671 27104
rect 34532 27100 34538 27102
rect 34605 27099 34671 27102
rect 40033 27162 40099 27165
rect 40166 27162 40172 27164
rect 40033 27160 40172 27162
rect 40033 27104 40038 27160
rect 40094 27104 40172 27160
rect 40033 27102 40172 27104
rect 40033 27099 40099 27102
rect 40166 27100 40172 27102
rect 40236 27100 40242 27164
rect 15009 27026 15075 27029
rect 17217 27026 17283 27029
rect 15009 27024 17283 27026
rect 15009 26968 15014 27024
rect 15070 26968 17222 27024
rect 17278 26968 17283 27024
rect 15009 26966 17283 26968
rect 15009 26963 15075 26966
rect 17217 26963 17283 26966
rect 23749 27026 23815 27029
rect 26509 27026 26575 27029
rect 23749 27024 26575 27026
rect 23749 26968 23754 27024
rect 23810 26968 26514 27024
rect 26570 26968 26575 27024
rect 23749 26966 26575 26968
rect 23749 26963 23815 26966
rect 26509 26963 26575 26966
rect 34646 26964 34652 27028
rect 34716 27026 34722 27028
rect 36353 27026 36419 27029
rect 34716 27024 36419 27026
rect 34716 26968 36358 27024
rect 36414 26968 36419 27024
rect 34716 26966 36419 26968
rect 34716 26964 34722 26966
rect 36353 26963 36419 26966
rect 16941 26890 17007 26893
rect 17493 26890 17559 26893
rect 19057 26890 19123 26893
rect 16941 26888 19123 26890
rect 16941 26832 16946 26888
rect 17002 26832 17498 26888
rect 17554 26832 19062 26888
rect 19118 26832 19123 26888
rect 16941 26830 19123 26832
rect 16941 26827 17007 26830
rect 17493 26827 17559 26830
rect 19057 26827 19123 26830
rect 20253 26890 20319 26893
rect 21173 26890 21239 26893
rect 20253 26888 21239 26890
rect 20253 26832 20258 26888
rect 20314 26832 21178 26888
rect 21234 26832 21239 26888
rect 20253 26830 21239 26832
rect 20253 26827 20319 26830
rect 21173 26827 21239 26830
rect 34145 26890 34211 26893
rect 40769 26890 40835 26893
rect 34145 26888 40835 26890
rect 34145 26832 34150 26888
rect 34206 26832 40774 26888
rect 40830 26832 40835 26888
rect 34145 26830 40835 26832
rect 34145 26827 34211 26830
rect 40769 26827 40835 26830
rect 35525 26754 35591 26757
rect 36997 26754 37063 26757
rect 35525 26752 37063 26754
rect 35525 26696 35530 26752
rect 35586 26696 37002 26752
rect 37058 26696 37063 26752
rect 35525 26694 37063 26696
rect 35525 26691 35591 26694
rect 36997 26691 37063 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4705 26618 4771 26621
rect 5993 26618 6059 26621
rect 35617 26618 35683 26621
rect 36537 26618 36603 26621
rect 4705 26616 6059 26618
rect 4705 26560 4710 26616
rect 4766 26560 5998 26616
rect 6054 26560 6059 26616
rect 4705 26558 6059 26560
rect 4705 26555 4771 26558
rect 5993 26555 6059 26558
rect 35344 26616 36603 26618
rect 35344 26560 35622 26616
rect 35678 26560 36542 26616
rect 36598 26560 36603 26616
rect 35344 26558 36603 26560
rect 5349 26482 5415 26485
rect 5809 26482 5875 26485
rect 5349 26480 5875 26482
rect 5349 26424 5354 26480
rect 5410 26424 5814 26480
rect 5870 26424 5875 26480
rect 5349 26422 5875 26424
rect 5349 26419 5415 26422
rect 5809 26419 5875 26422
rect 15469 26482 15535 26485
rect 16389 26482 16455 26485
rect 15469 26480 16455 26482
rect 15469 26424 15474 26480
rect 15530 26424 16394 26480
rect 16450 26424 16455 26480
rect 15469 26422 16455 26424
rect 15469 26419 15535 26422
rect 16389 26419 16455 26422
rect 33961 26482 34027 26485
rect 35344 26482 35404 26558
rect 35617 26555 35683 26558
rect 36537 26555 36603 26558
rect 42057 26618 42123 26621
rect 42813 26618 43613 26648
rect 42057 26616 43613 26618
rect 42057 26560 42062 26616
rect 42118 26560 43613 26616
rect 42057 26558 43613 26560
rect 42057 26555 42123 26558
rect 42813 26528 43613 26558
rect 33961 26480 35404 26482
rect 33961 26424 33966 26480
rect 34022 26424 35404 26480
rect 33961 26422 35404 26424
rect 33961 26419 34027 26422
rect 4705 26346 4771 26349
rect 5073 26346 5139 26349
rect 6177 26346 6243 26349
rect 4705 26344 6243 26346
rect 4705 26288 4710 26344
rect 4766 26288 5078 26344
rect 5134 26288 6182 26344
rect 6238 26288 6243 26344
rect 4705 26286 6243 26288
rect 4705 26283 4771 26286
rect 5073 26283 5139 26286
rect 6177 26283 6243 26286
rect 11973 26346 12039 26349
rect 17217 26346 17283 26349
rect 11973 26344 17283 26346
rect 11973 26288 11978 26344
rect 12034 26288 17222 26344
rect 17278 26288 17283 26344
rect 11973 26286 17283 26288
rect 11973 26283 12039 26286
rect 17217 26283 17283 26286
rect 31937 26346 32003 26349
rect 37181 26346 37247 26349
rect 31937 26344 37247 26346
rect 31937 26288 31942 26344
rect 31998 26288 37186 26344
rect 37242 26288 37247 26344
rect 31937 26286 37247 26288
rect 31937 26283 32003 26286
rect 37181 26283 37247 26286
rect 14457 26210 14523 26213
rect 18413 26210 18479 26213
rect 19149 26210 19215 26213
rect 14457 26208 19215 26210
rect 14457 26152 14462 26208
rect 14518 26152 18418 26208
rect 18474 26152 19154 26208
rect 19210 26152 19215 26208
rect 14457 26150 19215 26152
rect 14457 26147 14523 26150
rect 18413 26147 18479 26150
rect 19149 26147 19215 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 841 26074 907 26077
rect 798 26072 907 26074
rect 798 26016 846 26072
rect 902 26016 907 26072
rect 798 26011 907 26016
rect 14733 26074 14799 26077
rect 15745 26074 15811 26077
rect 14733 26072 15811 26074
rect 14733 26016 14738 26072
rect 14794 26016 15750 26072
rect 15806 26016 15811 26072
rect 14733 26014 15811 26016
rect 14733 26011 14799 26014
rect 15745 26011 15811 26014
rect 798 25968 858 26011
rect 0 25878 858 25968
rect 39021 25938 39087 25941
rect 41873 25938 41939 25941
rect 39021 25936 41939 25938
rect 39021 25880 39026 25936
rect 39082 25880 41878 25936
rect 41934 25880 41939 25936
rect 39021 25878 41939 25880
rect 0 25848 800 25878
rect 39021 25875 39087 25878
rect 41873 25875 41939 25878
rect 42057 25938 42123 25941
rect 42813 25938 43613 25968
rect 42057 25936 43613 25938
rect 42057 25880 42062 25936
rect 42118 25880 43613 25936
rect 42057 25878 43613 25880
rect 42057 25875 42123 25878
rect 42813 25848 43613 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25288
rect 1301 25258 1367 25261
rect 0 25256 1367 25258
rect 0 25200 1306 25256
rect 1362 25200 1367 25256
rect 0 25198 1367 25200
rect 0 25168 800 25198
rect 1301 25195 1367 25198
rect 13445 25258 13511 25261
rect 16941 25258 17007 25261
rect 13445 25256 17007 25258
rect 13445 25200 13450 25256
rect 13506 25200 16946 25256
rect 17002 25200 17007 25256
rect 13445 25198 17007 25200
rect 13445 25195 13511 25198
rect 16941 25195 17007 25198
rect 35157 25258 35223 25261
rect 35893 25258 35959 25261
rect 35157 25256 35959 25258
rect 35157 25200 35162 25256
rect 35218 25200 35898 25256
rect 35954 25200 35959 25256
rect 35157 25198 35959 25200
rect 35157 25195 35223 25198
rect 35893 25195 35959 25198
rect 41505 25258 41571 25261
rect 42813 25258 43613 25288
rect 41505 25256 43613 25258
rect 41505 25200 41510 25256
rect 41566 25200 43613 25256
rect 41505 25198 43613 25200
rect 41505 25195 41571 25198
rect 42813 25168 43613 25198
rect 22093 25122 22159 25125
rect 23565 25122 23631 25125
rect 22093 25120 23631 25122
rect 22093 25064 22098 25120
rect 22154 25064 23570 25120
rect 23626 25064 23631 25120
rect 22093 25062 23631 25064
rect 22093 25059 22159 25062
rect 23565 25059 23631 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 12709 24850 12775 24853
rect 16665 24850 16731 24853
rect 12709 24848 16731 24850
rect 12709 24792 12714 24848
rect 12770 24792 16670 24848
rect 16726 24792 16731 24848
rect 12709 24790 16731 24792
rect 12709 24787 12775 24790
rect 16665 24787 16731 24790
rect 22461 24850 22527 24853
rect 40953 24850 41019 24853
rect 22461 24848 41019 24850
rect 22461 24792 22466 24848
rect 22522 24792 40958 24848
rect 41014 24792 41019 24848
rect 22461 24790 41019 24792
rect 22461 24787 22527 24790
rect 40953 24787 41019 24790
rect 25589 24714 25655 24717
rect 40861 24714 40927 24717
rect 25589 24712 40927 24714
rect 25589 24656 25594 24712
rect 25650 24656 40866 24712
rect 40922 24656 40927 24712
rect 25589 24654 40927 24656
rect 25589 24651 25655 24654
rect 40861 24651 40927 24654
rect 18413 24578 18479 24581
rect 27981 24578 28047 24581
rect 18413 24576 28047 24578
rect 18413 24520 18418 24576
rect 18474 24520 27986 24576
rect 28042 24520 28047 24576
rect 18413 24518 28047 24520
rect 18413 24515 18479 24518
rect 27981 24515 28047 24518
rect 41505 24578 41571 24581
rect 42813 24578 43613 24608
rect 41505 24576 43613 24578
rect 41505 24520 41510 24576
rect 41566 24520 43613 24576
rect 41505 24518 43613 24520
rect 41505 24515 41571 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 42813 24488 43613 24518
rect 34930 24447 35246 24448
rect 19517 24442 19583 24445
rect 25221 24442 25287 24445
rect 26509 24442 26575 24445
rect 19517 24440 26575 24442
rect 19517 24384 19522 24440
rect 19578 24384 25226 24440
rect 25282 24384 26514 24440
rect 26570 24384 26575 24440
rect 19517 24382 26575 24384
rect 19517 24379 19583 24382
rect 25221 24379 25287 24382
rect 26509 24379 26575 24382
rect 7005 24306 7071 24309
rect 9213 24306 9279 24309
rect 7005 24304 9279 24306
rect 7005 24248 7010 24304
rect 7066 24248 9218 24304
rect 9274 24248 9279 24304
rect 7005 24246 9279 24248
rect 7005 24243 7071 24246
rect 9213 24243 9279 24246
rect 6085 24170 6151 24173
rect 7649 24170 7715 24173
rect 6085 24168 7715 24170
rect 6085 24112 6090 24168
rect 6146 24112 7654 24168
rect 7710 24112 7715 24168
rect 6085 24110 7715 24112
rect 6085 24107 6151 24110
rect 7649 24107 7715 24110
rect 18505 24170 18571 24173
rect 19425 24170 19491 24173
rect 18505 24168 19491 24170
rect 18505 24112 18510 24168
rect 18566 24112 19430 24168
rect 19486 24112 19491 24168
rect 18505 24110 19491 24112
rect 18505 24107 18571 24110
rect 19425 24107 19491 24110
rect 30005 24170 30071 24173
rect 39481 24170 39547 24173
rect 30005 24168 39547 24170
rect 30005 24112 30010 24168
rect 30066 24112 39486 24168
rect 39542 24112 39547 24168
rect 30005 24110 39547 24112
rect 30005 24107 30071 24110
rect 39481 24107 39547 24110
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 17861 23898 17927 23901
rect 20437 23898 20503 23901
rect 17861 23896 20503 23898
rect 17861 23840 17866 23896
rect 17922 23840 20442 23896
rect 20498 23840 20503 23896
rect 17861 23838 20503 23840
rect 17861 23835 17927 23838
rect 20437 23835 20503 23838
rect 40217 23898 40283 23901
rect 42813 23898 43613 23928
rect 40217 23896 43613 23898
rect 40217 23840 40222 23896
rect 40278 23840 43613 23896
rect 40217 23838 43613 23840
rect 40217 23835 40283 23838
rect 42813 23808 43613 23838
rect 17125 23762 17191 23765
rect 31293 23762 31359 23765
rect 17125 23760 31359 23762
rect 17125 23704 17130 23760
rect 17186 23704 31298 23760
rect 31354 23704 31359 23760
rect 17125 23702 31359 23704
rect 17125 23699 17191 23702
rect 31293 23699 31359 23702
rect 40033 23762 40099 23765
rect 41137 23762 41203 23765
rect 40033 23760 41203 23762
rect 40033 23704 40038 23760
rect 40094 23704 41142 23760
rect 41198 23704 41203 23760
rect 40033 23702 41203 23704
rect 40033 23699 40099 23702
rect 41137 23699 41203 23702
rect 17585 23490 17651 23493
rect 17718 23490 17724 23492
rect 17585 23488 17724 23490
rect 17585 23432 17590 23488
rect 17646 23432 17724 23488
rect 17585 23430 17724 23432
rect 17585 23427 17651 23430
rect 17718 23428 17724 23430
rect 17788 23428 17794 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23218 800 23248
rect 1577 23218 1643 23221
rect 0 23216 1643 23218
rect 0 23160 1582 23216
rect 1638 23160 1643 23216
rect 0 23158 1643 23160
rect 0 23128 800 23158
rect 1577 23155 1643 23158
rect 35525 23218 35591 23221
rect 36445 23218 36511 23221
rect 35525 23216 36511 23218
rect 35525 23160 35530 23216
rect 35586 23160 36450 23216
rect 36506 23160 36511 23216
rect 35525 23158 36511 23160
rect 35525 23155 35591 23158
rect 36445 23155 36511 23158
rect 39389 23218 39455 23221
rect 40125 23218 40191 23221
rect 41597 23218 41663 23221
rect 39389 23216 41663 23218
rect 39389 23160 39394 23216
rect 39450 23160 40130 23216
rect 40186 23160 41602 23216
rect 41658 23160 41663 23216
rect 39389 23158 41663 23160
rect 39389 23155 39455 23158
rect 40125 23155 40191 23158
rect 41597 23155 41663 23158
rect 42149 23218 42215 23221
rect 42813 23218 43613 23248
rect 42149 23216 43613 23218
rect 42149 23160 42154 23216
rect 42210 23160 43613 23216
rect 42149 23158 43613 23160
rect 42149 23155 42215 23158
rect 42813 23128 43613 23158
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 0 22538 800 22568
rect 1301 22538 1367 22541
rect 0 22536 1367 22538
rect 0 22480 1306 22536
rect 1362 22480 1367 22536
rect 0 22478 1367 22480
rect 0 22448 800 22478
rect 1301 22475 1367 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 5993 21994 6059 21997
rect 7465 21994 7531 21997
rect 5993 21992 7531 21994
rect 5993 21936 5998 21992
rect 6054 21936 7470 21992
rect 7526 21936 7531 21992
rect 5993 21934 7531 21936
rect 5993 21931 6059 21934
rect 7465 21931 7531 21934
rect 33501 21860 33567 21861
rect 33501 21858 33548 21860
rect 33456 21856 33548 21858
rect 33456 21800 33506 21856
rect 33456 21798 33548 21800
rect 33501 21796 33548 21798
rect 33612 21796 33618 21860
rect 33501 21795 33567 21796
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 33777 21316 33843 21317
rect 33726 21252 33732 21316
rect 33796 21314 33843 21316
rect 33796 21312 33888 21314
rect 33838 21256 33888 21312
rect 33796 21254 33888 21256
rect 33796 21252 33843 21254
rect 33777 21251 33843 21252
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 16021 21042 16087 21045
rect 17534 21042 17540 21044
rect 16021 21040 17540 21042
rect 16021 20984 16026 21040
rect 16082 20984 17540 21040
rect 16021 20982 17540 20984
rect 16021 20979 16087 20982
rect 17534 20980 17540 20982
rect 17604 20980 17610 21044
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19558 18532 19564 18596
rect 19628 18594 19634 18596
rect 19701 18594 19767 18597
rect 19628 18592 19767 18594
rect 19628 18536 19706 18592
rect 19762 18536 19767 18592
rect 19628 18534 19767 18536
rect 19628 18532 19634 18534
rect 19701 18531 19767 18534
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 841 17234 907 17237
rect 798 17232 907 17234
rect 798 17176 846 17232
rect 902 17176 907 17232
rect 798 17171 907 17176
rect 4889 17234 4955 17237
rect 5533 17234 5599 17237
rect 4889 17232 5599 17234
rect 4889 17176 4894 17232
rect 4950 17176 5538 17232
rect 5594 17176 5599 17232
rect 4889 17174 5599 17176
rect 4889 17171 4955 17174
rect 5533 17171 5599 17174
rect 798 17128 858 17171
rect 0 17038 858 17128
rect 5349 17098 5415 17101
rect 6729 17098 6795 17101
rect 31937 17100 32003 17101
rect 5349 17096 6795 17098
rect 5349 17040 5354 17096
rect 5410 17040 6734 17096
rect 6790 17040 6795 17096
rect 5349 17038 6795 17040
rect 0 17008 800 17038
rect 5349 17035 5415 17038
rect 6729 17035 6795 17038
rect 31886 17036 31892 17100
rect 31956 17098 32003 17100
rect 31956 17096 32048 17098
rect 31998 17040 32048 17096
rect 31956 17038 32048 17040
rect 31956 17036 32003 17038
rect 31937 17035 32003 17036
rect 4981 16962 5047 16965
rect 6453 16962 6519 16965
rect 4981 16960 6519 16962
rect 4981 16904 4986 16960
rect 5042 16904 6458 16960
rect 6514 16904 6519 16960
rect 4981 16902 6519 16904
rect 4981 16899 5047 16902
rect 6453 16899 6519 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 17125 16148 17191 16149
rect 17125 16146 17172 16148
rect 17080 16144 17172 16146
rect 17080 16088 17130 16144
rect 17080 16086 17172 16088
rect 17125 16084 17172 16086
rect 17236 16084 17242 16148
rect 17125 16083 17191 16084
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 0 15648 800 15678
rect 21817 15602 21883 15605
rect 22461 15602 22527 15605
rect 21817 15600 22527 15602
rect 21817 15544 21822 15600
rect 21878 15544 22466 15600
rect 22522 15544 22527 15600
rect 21817 15542 22527 15544
rect 21817 15539 21883 15542
rect 22461 15539 22527 15542
rect 27245 15332 27311 15333
rect 27245 15328 27292 15332
rect 27356 15330 27362 15332
rect 27245 15272 27250 15328
rect 27245 15268 27292 15272
rect 27356 15270 27402 15330
rect 27356 15268 27362 15270
rect 27245 15267 27311 15268
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 18045 15194 18111 15197
rect 19558 15194 19564 15196
rect 18045 15192 19564 15194
rect 18045 15136 18050 15192
rect 18106 15136 19564 15192
rect 18045 15134 19564 15136
rect 18045 15131 18111 15134
rect 19558 15132 19564 15134
rect 19628 15132 19634 15196
rect 25589 15194 25655 15197
rect 26233 15194 26299 15197
rect 25589 15192 26299 15194
rect 25589 15136 25594 15192
rect 25650 15136 26238 15192
rect 26294 15136 26299 15192
rect 25589 15134 26299 15136
rect 25589 15131 25655 15134
rect 26233 15131 26299 15134
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 0 13018 800 13048
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 1485 13018 1551 13021
rect 0 13016 1551 13018
rect 0 12960 1490 13016
rect 1546 12960 1551 13016
rect 0 12958 1551 12960
rect 0 12928 800 12958
rect 1485 12955 1551 12958
rect 28073 12882 28139 12885
rect 29545 12882 29611 12885
rect 28073 12880 29611 12882
rect 28073 12824 28078 12880
rect 28134 12824 29550 12880
rect 29606 12824 29611 12880
rect 28073 12822 29611 12824
rect 28073 12819 28139 12822
rect 29545 12819 29611 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 1209 12338 1275 12341
rect 33685 12340 33751 12341
rect 33685 12338 33732 12340
rect 0 12336 1275 12338
rect 0 12280 1214 12336
rect 1270 12280 1275 12336
rect 0 12278 1275 12280
rect 33640 12336 33732 12338
rect 33640 12280 33690 12336
rect 33640 12278 33732 12280
rect 0 12248 800 12278
rect 1209 12275 1275 12278
rect 33685 12276 33732 12278
rect 33796 12276 33802 12340
rect 33685 12275 33751 12276
rect 5901 12202 5967 12205
rect 6637 12202 6703 12205
rect 5901 12200 6703 12202
rect 5901 12144 5906 12200
rect 5962 12144 6642 12200
rect 6698 12144 6703 12200
rect 5901 12142 6703 12144
rect 5901 12139 5967 12142
rect 6637 12139 6703 12142
rect 32949 12202 33015 12205
rect 33542 12202 33548 12204
rect 32949 12200 33548 12202
rect 32949 12144 32954 12200
rect 33010 12144 33548 12200
rect 32949 12142 33548 12144
rect 32949 12139 33015 12142
rect 33542 12140 33548 12142
rect 33612 12140 33618 12204
rect 35709 12202 35775 12205
rect 33734 12200 35775 12202
rect 33734 12144 35714 12200
rect 35770 12144 35775 12200
rect 33734 12142 35775 12144
rect 32489 12066 32555 12069
rect 33734 12066 33794 12142
rect 35709 12139 35775 12142
rect 38929 12202 38995 12205
rect 39757 12202 39823 12205
rect 38929 12200 39823 12202
rect 38929 12144 38934 12200
rect 38990 12144 39762 12200
rect 39818 12144 39823 12200
rect 38929 12142 39823 12144
rect 38929 12139 38995 12142
rect 39757 12139 39823 12142
rect 32489 12064 33794 12066
rect 32489 12008 32494 12064
rect 32550 12008 33794 12064
rect 32489 12006 33794 12008
rect 32489 12003 32555 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 31845 11932 31911 11933
rect 31845 11930 31892 11932
rect 31800 11928 31892 11930
rect 31800 11872 31850 11928
rect 31800 11870 31892 11872
rect 31845 11868 31892 11870
rect 31956 11868 31962 11932
rect 31845 11867 31911 11868
rect 0 11658 800 11688
rect 3325 11658 3391 11661
rect 0 11656 3391 11658
rect 0 11600 3330 11656
rect 3386 11600 3391 11656
rect 0 11598 3391 11600
rect 0 11568 800 11598
rect 3325 11595 3391 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 27337 10980 27403 10981
rect 27286 10978 27292 10980
rect 27246 10918 27292 10978
rect 27356 10976 27403 10980
rect 27398 10920 27403 10976
rect 27286 10916 27292 10918
rect 27356 10916 27403 10920
rect 27337 10915 27403 10916
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 30281 6354 30347 6357
rect 32581 6354 32647 6357
rect 30281 6352 32647 6354
rect 30281 6296 30286 6352
rect 30342 6296 32586 6352
rect 32642 6296 32647 6352
rect 30281 6294 32647 6296
rect 30281 6291 30347 6294
rect 32581 6291 32647 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 42057 5538 42123 5541
rect 42813 5538 43613 5568
rect 42057 5536 43613 5538
rect 42057 5480 42062 5536
rect 42118 5480 43613 5536
rect 42057 5478 43613 5480
rect 42057 5475 42123 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 42813 5448 43613 5478
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 35596 43548 35660 43552
rect 35596 43492 35600 43548
rect 35600 43492 35656 43548
rect 35656 43492 35660 43548
rect 35596 43488 35660 43492
rect 35676 43548 35740 43552
rect 35676 43492 35680 43548
rect 35680 43492 35736 43548
rect 35736 43492 35740 43548
rect 35676 43488 35740 43492
rect 35756 43548 35820 43552
rect 35756 43492 35760 43548
rect 35760 43492 35816 43548
rect 35816 43492 35820 43548
rect 35756 43488 35820 43492
rect 35836 43548 35900 43552
rect 35836 43492 35840 43548
rect 35840 43492 35896 43548
rect 35896 43492 35900 43548
rect 35836 43488 35900 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 35596 42460 35660 42464
rect 35596 42404 35600 42460
rect 35600 42404 35656 42460
rect 35656 42404 35660 42460
rect 35596 42400 35660 42404
rect 35676 42460 35740 42464
rect 35676 42404 35680 42460
rect 35680 42404 35736 42460
rect 35736 42404 35740 42460
rect 35676 42400 35740 42404
rect 35756 42460 35820 42464
rect 35756 42404 35760 42460
rect 35760 42404 35816 42460
rect 35816 42404 35820 42460
rect 35756 42400 35820 42404
rect 35836 42460 35900 42464
rect 35836 42404 35840 42460
rect 35840 42404 35896 42460
rect 35896 42404 35900 42460
rect 35836 42400 35900 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 35596 41372 35660 41376
rect 35596 41316 35600 41372
rect 35600 41316 35656 41372
rect 35656 41316 35660 41372
rect 35596 41312 35660 41316
rect 35676 41372 35740 41376
rect 35676 41316 35680 41372
rect 35680 41316 35736 41372
rect 35736 41316 35740 41372
rect 35676 41312 35740 41316
rect 35756 41372 35820 41376
rect 35756 41316 35760 41372
rect 35760 41316 35816 41372
rect 35816 41316 35820 41372
rect 35756 41312 35820 41316
rect 35836 41372 35900 41376
rect 35836 41316 35840 41372
rect 35840 41316 35896 41372
rect 35896 41316 35900 41372
rect 35836 41312 35900 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 35596 40284 35660 40288
rect 35596 40228 35600 40284
rect 35600 40228 35656 40284
rect 35656 40228 35660 40284
rect 35596 40224 35660 40228
rect 35676 40284 35740 40288
rect 35676 40228 35680 40284
rect 35680 40228 35736 40284
rect 35736 40228 35740 40284
rect 35676 40224 35740 40228
rect 35756 40284 35820 40288
rect 35756 40228 35760 40284
rect 35760 40228 35816 40284
rect 35816 40228 35820 40284
rect 35756 40224 35820 40228
rect 35836 40284 35900 40288
rect 35836 40228 35840 40284
rect 35840 40228 35896 40284
rect 35896 40228 35900 40284
rect 35836 40224 35900 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 34652 38796 34716 38860
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 33916 38584 33980 38588
rect 33916 38528 33930 38584
rect 33930 38528 33980 38584
rect 33916 38524 33980 38528
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 22140 34232 22204 34236
rect 22140 34176 22154 34232
rect 22154 34176 22204 34232
rect 22140 34172 22204 34176
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 40172 33220 40236 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 17724 32404 17788 32468
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 24900 31180 24964 31244
rect 17540 31044 17604 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 36124 30636 36188 30700
rect 22324 30560 22388 30564
rect 22324 30504 22374 30560
rect 22374 30504 22388 30560
rect 22324 30500 22388 30504
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 34468 30364 34532 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 17172 29412 17236 29476
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 36124 29004 36188 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 22140 28460 22204 28524
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 22324 27704 22388 27708
rect 22324 27648 22374 27704
rect 22374 27648 22388 27704
rect 22324 27644 22388 27648
rect 24900 27644 24964 27708
rect 38700 27644 38764 27708
rect 23060 27568 23124 27572
rect 23060 27512 23074 27568
rect 23074 27512 23124 27568
rect 23060 27508 23124 27512
rect 33916 27508 33980 27572
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 34468 27100 34532 27164
rect 40172 27100 40236 27164
rect 34652 26964 34716 27028
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 17724 23428 17788 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 33548 21856 33612 21860
rect 33548 21800 33562 21856
rect 33562 21800 33612 21856
rect 33548 21796 33612 21800
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 33732 21312 33796 21316
rect 33732 21256 33782 21312
rect 33782 21256 33796 21312
rect 33732 21252 33796 21256
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 17540 20980 17604 21044
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19564 18532 19628 18596
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 31892 17096 31956 17100
rect 31892 17040 31942 17096
rect 31942 17040 31956 17096
rect 31892 17036 31956 17040
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 17172 16144 17236 16148
rect 17172 16088 17186 16144
rect 17186 16088 17236 16144
rect 17172 16084 17236 16088
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 27292 15328 27356 15332
rect 27292 15272 27306 15328
rect 27306 15272 27356 15328
rect 27292 15268 27356 15272
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 19564 15132 19628 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 33732 12336 33796 12340
rect 33732 12280 33746 12336
rect 33746 12280 33796 12336
rect 33732 12276 33796 12280
rect 33548 12140 33612 12204
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 31892 11928 31956 11932
rect 31892 11872 31906 11928
rect 31906 11872 31956 11928
rect 31892 11868 31956 11872
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 27292 10976 27356 10980
rect 27292 10920 27342 10976
rect 27342 10920 27356 10976
rect 27292 10916 27356 10920
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 43008 4528 43568
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 43552 5188 43568
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 34928 43008 35248 43568
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34651 38860 34717 38861
rect 34651 38796 34652 38860
rect 34716 38796 34717 38860
rect 34651 38795 34717 38796
rect 33915 38588 33981 38589
rect 33915 38524 33916 38588
rect 33980 38524 33981 38588
rect 33915 38523 33981 38524
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 22139 34236 22205 34237
rect 22139 34172 22140 34236
rect 22204 34172 22205 34236
rect 22139 34171 22205 34172
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 17723 32468 17789 32469
rect 17723 32404 17724 32468
rect 17788 32404 17789 32468
rect 17723 32403 17789 32404
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 17539 31108 17605 31109
rect 17539 31044 17540 31108
rect 17604 31044 17605 31108
rect 17539 31043 17605 31044
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 17171 29476 17237 29477
rect 17171 29412 17172 29476
rect 17236 29412 17237 29476
rect 17171 29411 17237 29412
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 17174 16149 17234 29411
rect 17542 21045 17602 31043
rect 17726 23493 17786 32403
rect 22142 28525 22202 34171
rect 24899 31244 24965 31245
rect 24899 31180 24900 31244
rect 24964 31180 24965 31244
rect 24899 31179 24965 31180
rect 22323 30564 22389 30565
rect 22323 30500 22324 30564
rect 22388 30500 22389 30564
rect 22323 30499 22389 30500
rect 22139 28524 22205 28525
rect 22139 28460 22140 28524
rect 22204 28460 22205 28524
rect 22139 28459 22205 28460
rect 22326 27709 22386 30499
rect 24902 27709 24962 31179
rect 22323 27708 22389 27709
rect 22323 27644 22324 27708
rect 22388 27644 22389 27708
rect 24899 27708 24965 27709
rect 22323 27643 22389 27644
rect 24899 27644 24900 27708
rect 24964 27644 24965 27708
rect 24899 27643 24965 27644
rect 33918 27573 33978 38523
rect 34467 30428 34533 30429
rect 34467 30364 34468 30428
rect 34532 30364 34533 30428
rect 34467 30363 34533 30364
rect 33915 27572 33981 27573
rect 33915 27508 33916 27572
rect 33980 27508 33981 27572
rect 33915 27507 33981 27508
rect 34470 27165 34530 30363
rect 34467 27164 34533 27165
rect 34467 27100 34468 27164
rect 34532 27100 34533 27164
rect 34467 27099 34533 27100
rect 34654 27029 34714 38795
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34651 27028 34717 27029
rect 34651 26964 34652 27028
rect 34716 26964 34717 27028
rect 34651 26963 34717 26964
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 17723 23492 17789 23493
rect 17723 23428 17724 23492
rect 17788 23428 17789 23492
rect 17723 23427 17789 23428
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 33547 21860 33613 21861
rect 33547 21796 33548 21860
rect 33612 21796 33613 21860
rect 33547 21795 33613 21796
rect 17539 21044 17605 21045
rect 17539 20980 17540 21044
rect 17604 20980 17605 21044
rect 17539 20979 17605 20980
rect 19563 18596 19629 18597
rect 19563 18532 19564 18596
rect 19628 18532 19629 18596
rect 19563 18531 19629 18532
rect 17171 16148 17237 16149
rect 17171 16084 17172 16148
rect 17236 16084 17237 16148
rect 17171 16083 17237 16084
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 19566 15197 19626 18531
rect 31891 17100 31957 17101
rect 31891 17036 31892 17100
rect 31956 17036 31957 17100
rect 31891 17035 31957 17036
rect 27291 15332 27357 15333
rect 27291 15268 27292 15332
rect 27356 15268 27357 15332
rect 27291 15267 27357 15268
rect 19563 15196 19629 15197
rect 19563 15132 19564 15196
rect 19628 15132 19629 15196
rect 19563 15131 19629 15132
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 27294 10981 27354 15267
rect 31894 11933 31954 17035
rect 33550 12205 33610 21795
rect 33731 21316 33797 21317
rect 33731 21252 33732 21316
rect 33796 21252 33797 21316
rect 33731 21251 33797 21252
rect 33734 12341 33794 21251
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 33731 12340 33797 12341
rect 33731 12276 33732 12340
rect 33796 12276 33797 12340
rect 33731 12275 33797 12276
rect 33547 12204 33613 12205
rect 33547 12140 33548 12204
rect 33612 12140 33613 12204
rect 33547 12139 33613 12140
rect 31891 11932 31957 11933
rect 31891 11868 31892 11932
rect 31956 11868 31957 11932
rect 31891 11867 31957 11868
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 27291 10980 27357 10981
rect 27291 10916 27292 10980
rect 27356 10916 27357 10980
rect 27291 10915 27357 10916
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 43552 35908 43568
rect 35588 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35908 43552
rect 35588 42464 35908 43488
rect 35588 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35908 42464
rect 35588 41376 35908 42400
rect 35588 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35908 41376
rect 35588 40288 35908 41312
rect 35588 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35908 40288
rect 35588 39200 35908 40224
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 40171 33284 40237 33285
rect 40171 33220 40172 33284
rect 40236 33220 40237 33284
rect 40171 33219 40237 33220
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 36123 30700 36189 30701
rect 36123 30636 36124 30700
rect 36188 30636 36189 30700
rect 36123 30635 36189 30636
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 36126 29069 36186 30635
rect 36123 29068 36189 29069
rect 36123 29004 36124 29068
rect 36188 29004 36189 29068
rect 36123 29003 36189 29004
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 38699 27708 38765 27709
rect 38699 27658 38700 27708
rect 38764 27658 38765 27708
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 40174 27165 40234 33219
rect 40171 27164 40237 27165
rect 40171 27100 40172 27164
rect 40236 27100 40237 27164
rect 40171 27099 40237 27100
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 22974 27572 23210 27658
rect 22974 27508 23060 27572
rect 23060 27508 23124 27572
rect 23124 27508 23210 27572
rect 22974 27422 23210 27508
rect 34970 36024 35206 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 38614 27644 38700 27658
rect 38700 27644 38764 27658
rect 38764 27644 38850 27658
rect 38614 27422 38850 27644
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 42552 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 42552 36920
rect 1056 36642 42552 36684
rect 1056 36260 42552 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 42552 36260
rect 1056 35982 42552 36024
rect 22932 27658 38892 27700
rect 22932 27422 22974 27658
rect 23210 27422 38614 27658
rect 38850 27422 38892 27658
rect 22932 27380 38892 27422
rect 1056 6284 42552 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 42552 6284
rect 1056 6006 42552 6048
rect 1056 5624 42552 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 42552 5624
rect 1056 5346 42552 5388
use sky130_fd_sc_hd__or4b_4  _1216_
timestamp 28801
transform -1 0 20424 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _1217_
timestamp 28801
transform 1 0 18124 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1218_
timestamp 28801
transform 1 0 18768 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1219_
timestamp 28801
transform -1 0 20148 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1220_
timestamp 28801
transform -1 0 23828 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1221_
timestamp 28801
transform 1 0 17756 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _1222_
timestamp 28801
transform 1 0 17480 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1223_
timestamp 28801
transform -1 0 17664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1224_
timestamp 28801
transform 1 0 17388 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1225_
timestamp 28801
transform -1 0 18952 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1226_
timestamp 28801
transform 1 0 17020 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1227_
timestamp 28801
transform 1 0 18400 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1228_
timestamp 28801
transform 1 0 20700 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 28801
transform -1 0 19688 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1230_
timestamp 28801
transform 1 0 19596 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1231_
timestamp 28801
transform 1 0 18492 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1232_
timestamp 28801
transform -1 0 20332 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1233_
timestamp 28801
transform 1 0 20056 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1234_
timestamp 28801
transform 1 0 19228 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1235_
timestamp 28801
transform 1 0 20976 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1236_
timestamp 28801
transform 1 0 22448 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1237_
timestamp 28801
transform 1 0 21896 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1238_
timestamp 28801
transform -1 0 21712 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 28801
transform -1 0 22540 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1240_
timestamp 28801
transform -1 0 21896 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1241_
timestamp 28801
transform -1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1242_
timestamp 28801
transform 1 0 21068 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1243_
timestamp 28801
transform 1 0 24104 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 28801
transform 1 0 22724 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 28801
transform -1 0 24196 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1246_
timestamp 28801
transform -1 0 23736 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1247_
timestamp 28801
transform -1 0 23460 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1248_
timestamp 28801
transform 1 0 23460 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1249_
timestamp 28801
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1250_
timestamp 28801
transform -1 0 25024 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1251_
timestamp 28801
transform 1 0 25576 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1252_
timestamp 28801
transform 1 0 26496 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1253_
timestamp 28801
transform 1 0 25668 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1254_
timestamp 28801
transform 1 0 25024 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1255_
timestamp 28801
transform -1 0 25852 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1256_
timestamp 28801
transform 1 0 24564 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1257_
timestamp 28801
transform -1 0 27416 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1258_
timestamp 28801
transform -1 0 27692 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1259_
timestamp 28801
transform 1 0 26128 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1260_
timestamp 28801
transform 1 0 26220 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1261_
timestamp 28801
transform -1 0 26496 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1262_
timestamp 28801
transform -1 0 27324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1263_
timestamp 28801
transform 1 0 27048 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1264_
timestamp 28801
transform 1 0 27692 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1265_
timestamp 28801
transform 1 0 28612 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1266_
timestamp 28801
transform 1 0 30084 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1267_
timestamp 28801
transform 1 0 30176 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 28801
transform 1 0 30544 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1269_
timestamp 28801
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1270_
timestamp 28801
transform 1 0 29532 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1271_
timestamp 28801
transform 1 0 30820 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 28801
transform -1 0 31096 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1273_
timestamp 28801
transform 1 0 30268 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1274_
timestamp 28801
transform 1 0 22632 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1275_
timestamp 28801
transform 1 0 30452 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1276_
timestamp 28801
transform 1 0 30084 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1277_
timestamp 28801
transform 1 0 30820 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1278_
timestamp 28801
transform -1 0 32108 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1279_
timestamp 28801
transform -1 0 31832 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1280_
timestamp 28801
transform -1 0 34224 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1281_
timestamp 28801
transform 1 0 32108 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1282_
timestamp 28801
transform -1 0 35788 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1283_
timestamp 28801
transform -1 0 36156 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1284_
timestamp 28801
transform 1 0 35696 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1285_
timestamp 28801
transform -1 0 36432 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1286_
timestamp 28801
transform -1 0 34960 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1287_
timestamp 28801
transform 1 0 34960 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1288_
timestamp 28801
transform 1 0 34776 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1289_
timestamp 28801
transform 1 0 35972 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1290_
timestamp 28801
transform -1 0 35972 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1291_
timestamp 28801
transform 1 0 34040 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1292_
timestamp 28801
transform 1 0 34684 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1293_
timestamp 28801
transform -1 0 35236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1294_
timestamp 28801
transform -1 0 36248 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1295_
timestamp 28801
transform 1 0 35236 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1296_
timestamp 28801
transform 1 0 34224 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1297_
timestamp 28801
transform 1 0 34224 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1298_
timestamp 28801
transform -1 0 35972 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1299_
timestamp 28801
transform 1 0 34684 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1300_
timestamp 28801
transform -1 0 34224 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1301_
timestamp 28801
transform -1 0 34684 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1302_
timestamp 28801
transform -1 0 34224 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1303_
timestamp 28801
transform -1 0 34316 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1304_
timestamp 28801
transform -1 0 33672 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1305_
timestamp 28801
transform 1 0 32476 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1306_
timestamp 28801
transform -1 0 21344 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _1307_
timestamp 28801
transform 1 0 18124 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1308_
timestamp 28801
transform 1 0 18032 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1309_
timestamp 28801
transform 1 0 18032 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 28801
transform -1 0 19504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1311_
timestamp 28801
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1312_
timestamp 28801
transform -1 0 18860 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1313_
timestamp 28801
transform 1 0 17756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1314_
timestamp 28801
transform 1 0 19412 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1315_
timestamp 28801
transform -1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1316_
timestamp 28801
transform -1 0 20700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1317_
timestamp 28801
transform -1 0 20332 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1318_
timestamp 28801
transform 1 0 19504 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1319_
timestamp 28801
transform 1 0 19228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _1320_
timestamp 28801
transform -1 0 20424 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1321_
timestamp 28801
transform -1 0 21712 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 28801
transform 1 0 21712 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1323_
timestamp 28801
transform -1 0 21712 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1324_
timestamp 28801
transform -1 0 23092 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1325_
timestamp 28801
transform -1 0 21988 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1326_
timestamp 28801
transform 1 0 21804 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _1327_
timestamp 28801
transform 1 0 21988 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1328_
timestamp 28801
transform 1 0 23092 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1329_
timestamp 28801
transform 1 0 23920 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1330_
timestamp 28801
transform 1 0 23828 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1331_
timestamp 28801
transform -1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1332_
timestamp 28801
transform 1 0 23000 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1333_
timestamp 28801
transform 1 0 22632 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _1334_
timestamp 28801
transform -1 0 23828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1335_
timestamp 28801
transform -1 0 25576 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1336_
timestamp 28801
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 28801
transform -1 0 26036 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1338_
timestamp 28801
transform -1 0 25576 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1339_
timestamp 28801
transform 1 0 24932 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1340_
timestamp 28801
transform -1 0 24932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1341_
timestamp 28801
transform 1 0 26312 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1342_
timestamp 28801
transform 1 0 25668 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1343_
timestamp 28801
transform 1 0 25576 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1344_
timestamp 28801
transform 1 0 24932 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1345_
timestamp 28801
transform 1 0 26128 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1346_
timestamp 28801
transform 1 0 26588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp 28801
transform 1 0 26956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1348_
timestamp 28801
transform 1 0 27140 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1349_
timestamp 28801
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1350_
timestamp 28801
transform -1 0 29900 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1351_
timestamp 28801
transform 1 0 28428 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1352_
timestamp 28801
transform 1 0 28704 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1353_
timestamp 28801
transform 1 0 28152 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1354_
timestamp 28801
transform 1 0 29716 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 28801
transform -1 0 31372 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1356_
timestamp 28801
transform -1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1357_
timestamp 28801
transform 1 0 30636 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1358_
timestamp 28801
transform 1 0 30268 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1359_
timestamp 28801
transform 1 0 32384 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1360_
timestamp 28801
transform 1 0 32660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1361_
timestamp 28801
transform -1 0 33948 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1362_
timestamp 28801
transform -1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1363_
timestamp 28801
transform 1 0 36156 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1364_
timestamp 28801
transform -1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1365_
timestamp 28801
transform -1 0 37168 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1366_
timestamp 28801
transform -1 0 35328 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1367_
timestamp 28801
transform 1 0 34868 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1368_
timestamp 28801
transform 1 0 35328 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1369_
timestamp 28801
transform -1 0 36984 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1370_
timestamp 28801
transform -1 0 35696 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1371_
timestamp 28801
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1372_
timestamp 28801
transform 1 0 36248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1373_
timestamp 28801
transform -1 0 36984 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1374_
timestamp 28801
transform 1 0 34776 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1375_
timestamp 28801
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1376_
timestamp 28801
transform 1 0 35512 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1377_
timestamp 28801
transform 1 0 34684 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1378_
timestamp 28801
transform 1 0 30912 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1379_
timestamp 28801
transform -1 0 31740 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1380_
timestamp 28801
transform 1 0 31188 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1381_
timestamp 28801
transform 1 0 30360 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1382_
timestamp 28801
transform 1 0 9016 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1383_
timestamp 28801
transform -1 0 37904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1384_
timestamp 28801
transform 1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1385_
timestamp 28801
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1386_
timestamp 28801
transform -1 0 22448 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1387_
timestamp 28801
transform 1 0 22540 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1388_
timestamp 28801
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1389_
timestamp 28801
transform 1 0 24564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1390_
timestamp 28801
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1391_
timestamp 28801
transform 1 0 28796 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1392_
timestamp 28801
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1393_
timestamp 28801
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1394_
timestamp 28801
transform 1 0 32108 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1395_
timestamp 28801
transform 1 0 34684 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1396_
timestamp 28801
transform 1 0 35696 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1397_
timestamp 28801
transform 1 0 35972 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1398_
timestamp 28801
transform 1 0 37260 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1399_
timestamp 28801
transform 1 0 14076 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1400_
timestamp 28801
transform 1 0 14720 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1401_
timestamp 28801
transform 1 0 16836 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1402_
timestamp 28801
transform 1 0 15180 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1403_
timestamp 28801
transform 1 0 15916 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1404_
timestamp 28801
transform 1 0 16652 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1405_
timestamp 28801
transform 1 0 18308 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1406_
timestamp 28801
transform 1 0 19228 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1407_
timestamp 28801
transform 1 0 20700 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1408_
timestamp 28801
transform 1 0 22448 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1409_
timestamp 28801
transform 1 0 24380 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1410_
timestamp 28801
transform 1 0 25668 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1411_
timestamp 28801
transform 1 0 27416 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1412_
timestamp 28801
transform 1 0 28428 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1413_
timestamp 28801
transform 1 0 30452 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1414_
timestamp 28801
transform 1 0 33396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1415_
timestamp 28801
transform 1 0 35788 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1416_
timestamp 28801
transform 1 0 35696 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1417_
timestamp 28801
transform 1 0 35972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1418_
timestamp 28801
transform 1 0 36156 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1419_
timestamp 28801
transform 1 0 32108 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1420_
timestamp 28801
transform 1 0 17296 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1421_
timestamp 28801
transform -1 0 19872 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1422_
timestamp 28801
transform -1 0 19872 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1423_
timestamp 28801
transform -1 0 22816 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1424_
timestamp 28801
transform 1 0 22080 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1425_
timestamp 28801
transform -1 0 25760 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1426_
timestamp 28801
transform 1 0 24656 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1427_
timestamp 28801
transform 1 0 27508 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1428_
timestamp 28801
transform -1 0 29992 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1429_
timestamp 28801
transform 1 0 30452 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1430_
timestamp 28801
transform -1 0 35236 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1431_
timestamp 28801
transform -1 0 42228 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1432_
timestamp 28801
transform 1 0 39560 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1433_
timestamp 28801
transform -1 0 40480 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 28801
transform 1 0 39100 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1435_
timestamp 28801
transform -1 0 35328 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1436_
timestamp 28801
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1437_
timestamp 28801
transform 1 0 17112 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1438_
timestamp 28801
transform 1 0 17664 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1439_
timestamp 28801
transform 1 0 17020 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1440_
timestamp 28801
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1441_
timestamp 28801
transform 1 0 22724 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1442_
timestamp 28801
transform 1 0 24380 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1443_
timestamp 28801
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1444_
timestamp 28801
transform 1 0 27140 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1445_
timestamp 28801
transform 1 0 29532 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1446_
timestamp 28801
transform 1 0 33948 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1447_
timestamp 28801
transform -1 0 38548 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1448_
timestamp 28801
transform 1 0 40204 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1449_
timestamp 28801
transform 1 0 41124 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1450_
timestamp 28801
transform 1 0 37260 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1451_
timestamp 28801
transform 1 0 40572 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1452_
timestamp 28801
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1453_
timestamp 28801
transform 1 0 19136 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1454_
timestamp 28801
transform 1 0 18308 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1455_
timestamp 28801
transform 1 0 22172 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1456_
timestamp 28801
transform 1 0 22540 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1457_
timestamp 28801
transform 1 0 24472 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1458_
timestamp 28801
transform 1 0 25484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1459_
timestamp 28801
transform 1 0 26956 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1460_
timestamp 28801
transform -1 0 29256 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1461_
timestamp 28801
transform 1 0 29992 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1462_
timestamp 28801
transform 1 0 32936 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1463_
timestamp 28801
transform 1 0 32108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1464_
timestamp 28801
transform 1 0 34684 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1465_
timestamp 28801
transform 1 0 36340 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1466_
timestamp 28801
transform 1 0 34868 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 28801
transform 1 0 33212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1468_
timestamp 28801
transform 1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1469_
timestamp 28801
transform 1 0 18676 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1470_
timestamp 28801
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1471_
timestamp 28801
transform 1 0 18584 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1472_
timestamp 28801
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1473_
timestamp 28801
transform 1 0 19872 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1474_
timestamp 28801
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1475_
timestamp 28801
transform 1 0 19688 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1476_
timestamp 28801
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1477_
timestamp 28801
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1478_
timestamp 28801
transform -1 0 21712 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _1479_
timestamp 28801
transform 1 0 19964 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1480_
timestamp 28801
transform 1 0 20332 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1481_
timestamp 28801
transform 1 0 20516 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1482_
timestamp 28801
transform -1 0 21436 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1483_
timestamp 28801
transform -1 0 23184 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1484_
timestamp 28801
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1485_
timestamp 28801
transform -1 0 22080 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1486_
timestamp 28801
transform -1 0 22448 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1487_
timestamp 28801
transform 1 0 20792 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1488_
timestamp 28801
transform -1 0 21712 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1489_
timestamp 28801
transform 1 0 25760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1490_
timestamp 28801
transform -1 0 26312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1491_
timestamp 28801
transform -1 0 24748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1492_
timestamp 28801
transform 1 0 20792 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 28801
transform 1 0 23736 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1494_
timestamp 28801
transform -1 0 24288 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1495_
timestamp 28801
transform -1 0 24104 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1496_
timestamp 28801
transform -1 0 26588 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1497_
timestamp 28801
transform 1 0 26772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1498_
timestamp 28801
transform -1 0 26036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1499_
timestamp 28801
transform 1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1500_
timestamp 28801
transform -1 0 25300 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1501_
timestamp 28801
transform -1 0 26496 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1502_
timestamp 28801
transform -1 0 26772 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1503_
timestamp 28801
transform 1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1504_
timestamp 28801
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1505_
timestamp 28801
transform 1 0 26772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1506_
timestamp 28801
transform -1 0 29348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1507_
timestamp 28801
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 28801
transform 1 0 27416 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1509_
timestamp 28801
transform 1 0 28428 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1510_
timestamp 28801
transform 1 0 29072 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1511_
timestamp 28801
transform -1 0 30820 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1512_
timestamp 28801
transform 1 0 30176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1513_
timestamp 28801
transform -1 0 29440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1514_
timestamp 28801
transform -1 0 29716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1515_
timestamp 28801
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1516_
timestamp 28801
transform 1 0 28888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1517_
timestamp 28801
transform 1 0 27876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1518_
timestamp 28801
transform 1 0 33580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1519_
timestamp 28801
transform -1 0 33672 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1520_
timestamp 28801
transform -1 0 33396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1521_
timestamp 28801
transform -1 0 29348 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1522_
timestamp 28801
transform 1 0 31740 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1523_
timestamp 28801
transform -1 0 32844 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1524_
timestamp 28801
transform -1 0 31832 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1525_
timestamp 28801
transform -1 0 35604 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1526_
timestamp 28801
transform -1 0 35604 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1527_
timestamp 28801
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1528_
timestamp 28801
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1529_
timestamp 28801
transform -1 0 36064 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1530_
timestamp 28801
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1531_
timestamp 28801
transform -1 0 40296 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1532_
timestamp 28801
transform 1 0 41032 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1533_
timestamp 28801
transform -1 0 42228 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1534_
timestamp 28801
transform 1 0 32476 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1535_
timestamp 28801
transform 1 0 36064 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1536_
timestamp 28801
transform 1 0 37260 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1537_
timestamp 28801
transform -1 0 38548 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1538_
timestamp 28801
transform -1 0 42136 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1539_
timestamp 28801
transform -1 0 41860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1540_
timestamp 28801
transform -1 0 40204 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1541_
timestamp 28801
transform 1 0 41032 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1542_
timestamp 28801
transform -1 0 40848 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 28801
transform -1 0 39192 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1544_
timestamp 28801
transform 1 0 39836 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1545_
timestamp 28801
transform 1 0 39468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1546_
timestamp 28801
transform -1 0 40204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1547_
timestamp 28801
transform -1 0 40204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1548_
timestamp 28801
transform 1 0 38916 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1549_
timestamp 28801
transform 1 0 37996 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1550_
timestamp 28801
transform -1 0 41584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1551_
timestamp 28801
transform -1 0 41308 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1552_
timestamp 28801
transform -1 0 39652 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1553_
timestamp 28801
transform 1 0 39192 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1554_
timestamp 28801
transform 1 0 38640 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1555_
timestamp 28801
transform -1 0 40572 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1556_
timestamp 28801
transform -1 0 34960 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1557_
timestamp 28801
transform 1 0 38456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1558_
timestamp 28801
transform 1 0 33948 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1559_
timestamp 28801
transform 1 0 34960 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1560_
timestamp 28801
transform 1 0 15732 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1561_
timestamp 28801
transform 1 0 16836 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1562_
timestamp 28801
transform -1 0 18216 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1563_
timestamp 28801
transform 1 0 16560 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1564_
timestamp 28801
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1565_
timestamp 28801
transform 1 0 18308 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1566_
timestamp 28801
transform 1 0 17940 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1567_
timestamp 28801
transform 1 0 30268 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1568_
timestamp 28801
transform -1 0 29440 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1569_
timestamp 28801
transform -1 0 31556 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1570_
timestamp 28801
transform 1 0 33304 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1571_
timestamp 28801
transform -1 0 33304 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1572_
timestamp 28801
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1573_
timestamp 28801
transform -1 0 34776 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1574_
timestamp 28801
transform -1 0 38640 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1575_
timestamp 28801
transform -1 0 39560 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1576_
timestamp 28801
transform 1 0 37812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1577_
timestamp 28801
transform -1 0 39376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1578_
timestamp 28801
transform -1 0 40388 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1579_
timestamp 28801
transform -1 0 39744 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1580_
timestamp 28801
transform -1 0 40112 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1581_
timestamp 28801
transform 1 0 40112 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1582_
timestamp 28801
transform -1 0 40296 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1583_
timestamp 28801
transform -1 0 40204 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1584_
timestamp 28801
transform 1 0 39376 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1585_
timestamp 28801
transform -1 0 39744 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1586_
timestamp 28801
transform 1 0 40020 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1587_
timestamp 28801
transform 1 0 38088 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1588_
timestamp 28801
transform 1 0 36800 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1589_
timestamp 28801
transform -1 0 37812 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1590_
timestamp 28801
transform 1 0 33672 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1591_
timestamp 28801
transform -1 0 33120 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1592_
timestamp 28801
transform -1 0 34500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1593_
timestamp 28801
transform -1 0 34316 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1594_
timestamp 28801
transform -1 0 31188 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1595_
timestamp 28801
transform -1 0 31832 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1596_
timestamp 28801
transform 1 0 31188 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1597_
timestamp 28801
transform -1 0 31924 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1598_
timestamp 28801
transform 1 0 28980 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1599_
timestamp 28801
transform 1 0 27784 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1600_
timestamp 28801
transform -1 0 28520 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1601_
timestamp 28801
transform 1 0 28520 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1602_
timestamp 28801
transform -1 0 27048 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1603_
timestamp 28801
transform -1 0 27232 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1604_
timestamp 28801
transform -1 0 26496 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1605_
timestamp 28801
transform 1 0 25760 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1606_
timestamp 28801
transform 1 0 25668 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1607_
timestamp 28801
transform -1 0 25024 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1608_
timestamp 28801
transform -1 0 25484 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1609_
timestamp 28801
transform 1 0 24748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1610_
timestamp 28801
transform -1 0 23920 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1611_
timestamp 28801
transform 1 0 23920 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1612_
timestamp 28801
transform -1 0 24748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1613_
timestamp 28801
transform 1 0 22264 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1614_
timestamp 28801
transform 1 0 21252 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1615_
timestamp 28801
transform 1 0 21068 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1616_
timestamp 28801
transform 1 0 21252 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1617_
timestamp 28801
transform -1 0 22172 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1618_
timestamp 28801
transform 1 0 15916 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1619_
timestamp 28801
transform -1 0 19504 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1620_
timestamp 28801
transform -1 0 17572 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1621_
timestamp 28801
transform 1 0 18584 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1622_
timestamp 28801
transform -1 0 20792 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1623_
timestamp 28801
transform -1 0 20792 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1624_
timestamp 28801
transform -1 0 21528 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1625_
timestamp 28801
transform -1 0 24840 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1626_
timestamp 28801
transform -1 0 25576 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1627_
timestamp 28801
transform 1 0 24932 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1628_
timestamp 28801
transform -1 0 27692 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1629_
timestamp 28801
transform 1 0 28796 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1630_
timestamp 28801
transform 1 0 28060 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1631_
timestamp 28801
transform -1 0 32016 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1632_
timestamp 28801
transform 1 0 32752 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1633_
timestamp 28801
transform -1 0 33856 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1634_
timestamp 28801
transform -1 0 37536 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1635_
timestamp 28801
transform 1 0 37904 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1636_
timestamp 28801
transform 1 0 37904 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1637_
timestamp 28801
transform -1 0 37628 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1638_
timestamp 28801
transform 1 0 37168 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1639_
timestamp 28801
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1640_
timestamp 28801
transform -1 0 31556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1641_
timestamp 28801
transform -1 0 31188 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1642_
timestamp 28801
transform -1 0 30728 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1643_
timestamp 28801
transform -1 0 31372 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1644_
timestamp 28801
transform 1 0 18308 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1645_
timestamp 28801
transform 1 0 18492 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1646_
timestamp 28801
transform 1 0 20608 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1647_
timestamp 28801
transform -1 0 20516 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1648_
timestamp 28801
transform 1 0 20240 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1649_
timestamp 28801
transform 1 0 19320 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1650_
timestamp 28801
transform 1 0 19596 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1651_
timestamp 28801
transform -1 0 21252 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1652_
timestamp 28801
transform 1 0 20516 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1653_
timestamp 28801
transform 1 0 21988 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1654_
timestamp 28801
transform 1 0 21344 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1655_
timestamp 28801
transform 1 0 20976 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1656_
timestamp 28801
transform 1 0 21252 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1657_
timestamp 28801
transform -1 0 23000 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1658_
timestamp 28801
transform 1 0 21804 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1659_
timestamp 28801
transform -1 0 22172 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1660_
timestamp 28801
transform 1 0 22448 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1661_
timestamp 28801
transform 1 0 22448 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1662_
timestamp 28801
transform 1 0 22908 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1663_
timestamp 28801
transform 1 0 24380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1664_
timestamp 28801
transform 1 0 25208 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1665_
timestamp 28801
transform 1 0 24564 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1666_
timestamp 28801
transform 1 0 25024 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 28801
transform 1 0 25484 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1668_
timestamp 28801
transform 1 0 25576 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1669_
timestamp 28801
transform -1 0 26496 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1670_
timestamp 28801
transform 1 0 25668 0 -1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1671_
timestamp 28801
transform -1 0 27048 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1672_
timestamp 28801
transform 1 0 27048 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1673_
timestamp 28801
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1674_
timestamp 28801
transform -1 0 28612 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _1675_
timestamp 28801
transform -1 0 28152 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1676_
timestamp 28801
transform 1 0 27784 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1677_
timestamp 28801
transform 1 0 27876 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 28801
transform 1 0 27968 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _1679_
timestamp 28801
transform 1 0 28060 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1680_
timestamp 28801
transform -1 0 31556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1681_
timestamp 28801
transform 1 0 28152 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1682_
timestamp 28801
transform 1 0 28520 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 28801
transform 1 0 29072 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1684_
timestamp 28801
transform 1 0 28612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1685_
timestamp 28801
transform 1 0 30084 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1686_
timestamp 28801
transform -1 0 33488 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1687_
timestamp 28801
transform 1 0 32108 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1688_
timestamp 28801
transform -1 0 31004 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 28801
transform -1 0 23644 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1690_
timestamp 28801
transform 1 0 31740 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1691_
timestamp 28801
transform -1 0 36984 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1692_
timestamp 28801
transform -1 0 33028 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1693_
timestamp 28801
transform -1 0 32476 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1694_
timestamp 28801
transform 1 0 32200 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1695_
timestamp 28801
transform 1 0 32108 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1696_
timestamp 28801
transform 1 0 32844 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1697_
timestamp 28801
transform -1 0 36708 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1698_
timestamp 28801
transform -1 0 39008 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1699_
timestamp 28801
transform -1 0 37904 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1700_
timestamp 28801
transform -1 0 36432 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1701_
timestamp 28801
transform 1 0 35604 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1702_
timestamp 28801
transform -1 0 34592 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1703_
timestamp 28801
transform -1 0 38640 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1704_
timestamp 28801
transform -1 0 38088 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1705_
timestamp 28801
transform -1 0 34592 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1706_
timestamp 28801
transform -1 0 35328 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1707_
timestamp 28801
transform 1 0 34684 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1708_
timestamp 28801
transform -1 0 35880 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1709_
timestamp 28801
transform 1 0 35052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1710_
timestamp 28801
transform 1 0 37996 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1711_
timestamp 28801
transform -1 0 37168 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1712_
timestamp 28801
transform -1 0 36616 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 28801
transform 1 0 35512 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1714_
timestamp 28801
transform 1 0 35052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1715_
timestamp 28801
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1716_
timestamp 28801
transform 1 0 34684 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1717_
timestamp 28801
transform -1 0 35972 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1718_
timestamp 28801
transform -1 0 36340 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1719_
timestamp 28801
transform 1 0 34868 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1720_
timestamp 28801
transform 1 0 35328 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1721_
timestamp 28801
transform 1 0 30820 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1722_
timestamp 28801
transform 1 0 31372 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1723_
timestamp 28801
transform 1 0 31924 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1724_
timestamp 28801
transform 1 0 32200 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1725_
timestamp 28801
transform -1 0 19228 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1726_
timestamp 28801
transform 1 0 19228 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1727_
timestamp 28801
transform 1 0 15640 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1728_
timestamp 28801
transform -1 0 17112 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1729_
timestamp 28801
transform 1 0 16652 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1730_
timestamp 28801
transform 1 0 17480 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1731_
timestamp 28801
transform 1 0 16652 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1732_
timestamp 28801
transform 1 0 20332 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 28801
transform 1 0 19228 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1734_
timestamp 28801
transform -1 0 22908 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1735_
timestamp 28801
transform 1 0 22448 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 28801
transform 1 0 24840 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1737_
timestamp 28801
transform 1 0 24380 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1738_
timestamp 28801
transform 1 0 25852 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1739_
timestamp 28801
transform 1 0 25208 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1740_
timestamp 28801
transform 1 0 27876 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1741_
timestamp 28801
transform 1 0 27508 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1742_
timestamp 28801
transform 1 0 29992 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1743_
timestamp 28801
transform 1 0 29900 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1744_
timestamp 28801
transform 1 0 34316 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1745_
timestamp 28801
transform 1 0 33120 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 28801
transform 1 0 39284 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1747_
timestamp 28801
transform 1 0 39192 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 28801
transform 1 0 41124 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1749_
timestamp 28801
transform 1 0 41032 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 28801
transform 1 0 40940 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1751_
timestamp 28801
transform 1 0 40112 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 28801
transform 1 0 38732 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1753_
timestamp 28801
transform 1 0 38548 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 28801
transform 1 0 34316 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1755_
timestamp 28801
transform 1 0 33948 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 28801
transform 1 0 30176 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1757_
timestamp 28801
transform 1 0 29808 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1758_
timestamp 28801
transform -1 0 16284 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 28801
transform 1 0 15640 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1760_
timestamp 28801
transform 1 0 17756 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 28801
transform 1 0 17480 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1762_
timestamp 28801
transform 1 0 20516 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 28801
transform 1 0 20056 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1764_
timestamp 28801
transform 1 0 22908 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1765_
timestamp 28801
transform 1 0 22632 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1766_
timestamp 28801
transform 1 0 25668 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 28801
transform 1 0 24840 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1768_
timestamp 28801
transform 1 0 26956 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 28801
transform 1 0 26036 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1770_
timestamp 28801
transform 1 0 27876 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1771_
timestamp 28801
transform 1 0 27600 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1772_
timestamp 28801
transform 1 0 30820 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 28801
transform 1 0 30084 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1774_
timestamp 28801
transform 1 0 35144 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 28801
transform 1 0 34684 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 28801
transform 1 0 38364 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1777_
timestamp 28801
transform 1 0 37260 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 28801
transform 1 0 40296 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1779_
timestamp 28801
transform 1 0 39836 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1780_
timestamp 28801
transform 1 0 40848 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1781_
timestamp 28801
transform 1 0 40664 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 28801
transform 1 0 37904 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1783_
timestamp 28801
transform 1 0 37628 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1784_
timestamp 28801
transform 1 0 33488 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1785_
timestamp 28801
transform 1 0 32844 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1786_
timestamp 28801
transform 1 0 31096 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 28801
transform 1 0 30268 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1788_
timestamp 28801
transform -1 0 13432 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 28801
transform 1 0 14076 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1790_
timestamp 28801
transform 1 0 22632 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1791_
timestamp 28801
transform 1 0 14904 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1792_
timestamp 28801
transform -1 0 14996 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1793_
timestamp 28801
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1794_
timestamp 28801
transform -1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1795_
timestamp 28801
transform 1 0 14812 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1796_
timestamp 28801
transform 1 0 16192 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1797_
timestamp 28801
transform -1 0 16192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1798_
timestamp 28801
transform -1 0 15640 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1799_
timestamp 28801
transform -1 0 17848 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1800_
timestamp 28801
transform 1 0 16652 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 28801
transform -1 0 20056 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 28801
transform 1 0 16652 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1803_
timestamp 28801
transform -1 0 22632 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 28801
transform 1 0 21804 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1805_
timestamp 28801
transform 1 0 23460 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1806_
timestamp 28801
transform 1 0 23092 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1807_
timestamp 28801
transform -1 0 26036 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1808_
timestamp 28801
transform 1 0 24196 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1809_
timestamp 28801
transform -1 0 27048 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1810_
timestamp 28801
transform 1 0 25944 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1811_
timestamp 28801
transform -1 0 28704 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1812_
timestamp 28801
transform 1 0 27508 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1813_
timestamp 28801
transform -1 0 30176 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1814_
timestamp 28801
transform 1 0 29532 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1815_
timestamp 28801
transform -1 0 32936 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1816_
timestamp 28801
transform 1 0 32476 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 28801
transform -1 0 38916 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1818_
timestamp 28801
transform 1 0 38732 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 28801
transform -1 0 40204 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1820_
timestamp 28801
transform 1 0 40296 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1821_
timestamp 28801
transform -1 0 40572 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1822_
timestamp 28801
transform 1 0 40664 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1823_
timestamp 28801
transform -1 0 38272 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1824_
timestamp 28801
transform 1 0 38180 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1825_
timestamp 28801
transform -1 0 35512 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1826_
timestamp 28801
transform 1 0 39836 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1827_
timestamp 28801
transform 1 0 32108 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1828_
timestamp 28801
transform 1 0 31004 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1829_
timestamp 28801
transform -1 0 17480 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1830_
timestamp 28801
transform 1 0 15548 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_2  _1831_
timestamp 28801
transform 1 0 13432 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1832_
timestamp 28801
transform -1 0 13892 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1833_
timestamp 28801
transform 1 0 13616 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1834_
timestamp 28801
transform 1 0 13432 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1835_
timestamp 28801
transform 1 0 11684 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1836_
timestamp 28801
transform 1 0 12236 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1837_
timestamp 28801
transform 1 0 12052 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1838_
timestamp 28801
transform 1 0 14076 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1839_
timestamp 28801
transform -1 0 12236 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1840_
timestamp 28801
transform 1 0 16376 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1841_
timestamp 28801
transform 1 0 18676 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1842_
timestamp 28801
transform 1 0 20516 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1843_
timestamp 28801
transform 1 0 23736 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1844_
timestamp 28801
transform 1 0 24748 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1845_
timestamp 28801
transform 1 0 25760 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1846_
timestamp 28801
transform 1 0 27692 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1847_
timestamp 28801
transform 1 0 29900 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1848_
timestamp 28801
transform 1 0 32108 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1849_
timestamp 28801
transform 1 0 40112 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1850_
timestamp 28801
transform 1 0 39836 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1851_
timestamp 28801
transform 1 0 41400 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1852_
timestamp 28801
transform 1 0 38088 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1853_
timestamp 28801
transform 1 0 33672 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1854_
timestamp 28801
transform 1 0 30360 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1855_
timestamp 28801
transform 1 0 14444 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1856_
timestamp 28801
transform -1 0 17296 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1857_
timestamp 28801
transform -1 0 17756 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1858_
timestamp 28801
transform 1 0 21436 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1859_
timestamp 28801
transform 1 0 22816 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1860_
timestamp 28801
transform 1 0 24840 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1861_
timestamp 28801
transform 1 0 26036 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1862_
timestamp 28801
transform 1 0 27600 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1863_
timestamp 28801
transform 1 0 29532 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1864_
timestamp 28801
transform 1 0 34960 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1865_
timestamp 28801
transform 1 0 38180 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1866_
timestamp 28801
transform 1 0 40940 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1867_
timestamp 28801
transform 1 0 40112 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1868_
timestamp 28801
transform 1 0 37260 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1869_
timestamp 28801
transform 1 0 33304 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1870_
timestamp 28801
transform 1 0 31188 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1871_
timestamp 28801
transform 1 0 15548 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1872_
timestamp 28801
transform 1 0 13432 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1873_
timestamp 28801
transform 1 0 12604 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1874_
timestamp 28801
transform -1 0 12788 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1875_
timestamp 28801
transform -1 0 13800 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1876_
timestamp 28801
transform 1 0 10488 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1877_
timestamp 28801
transform 1 0 11500 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1878_
timestamp 28801
transform 1 0 11500 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1879_
timestamp 28801
transform 1 0 11500 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1880_
timestamp 28801
transform -1 0 17020 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1881_
timestamp 28801
transform -1 0 15548 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1882_
timestamp 28801
transform -1 0 13524 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1883_
timestamp 28801
transform -1 0 14996 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1884_
timestamp 28801
transform -1 0 14536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1885_
timestamp 28801
transform -1 0 17296 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1886_
timestamp 28801
transform 1 0 18308 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1887_
timestamp 28801
transform 1 0 18032 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1888_
timestamp 28801
transform -1 0 17388 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1889_
timestamp 28801
transform 1 0 16284 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1890_
timestamp 28801
transform 1 0 16928 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1891_
timestamp 28801
transform -1 0 19688 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1892_
timestamp 28801
transform -1 0 21804 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1893_
timestamp 28801
transform -1 0 22080 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1894_
timestamp 28801
transform 1 0 19136 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1895_
timestamp 28801
transform 1 0 19780 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1896_
timestamp 28801
transform 1 0 19872 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1897_
timestamp 28801
transform -1 0 20976 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1898_
timestamp 28801
transform 1 0 20976 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1899_
timestamp 28801
transform 1 0 21528 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1900_
timestamp 28801
transform -1 0 22540 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1901_
timestamp 28801
transform 1 0 21896 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1902_
timestamp 28801
transform 1 0 23276 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1903_
timestamp 28801
transform 1 0 23460 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1904_
timestamp 28801
transform 1 0 24380 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1905_
timestamp 28801
transform 1 0 26128 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1906_
timestamp 28801
transform -1 0 41308 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1907_
timestamp 28801
transform 1 0 40480 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1908_
timestamp 28801
transform 1 0 27600 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1909_
timestamp 28801
transform -1 0 38916 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1910_
timestamp 28801
transform -1 0 37904 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1911_
timestamp 28801
transform 1 0 28704 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1912_
timestamp 28801
transform -1 0 39744 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1913_
timestamp 28801
transform 1 0 39284 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1914_
timestamp 28801
transform 1 0 30176 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1915_
timestamp 28801
transform -1 0 39744 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1916_
timestamp 28801
transform 1 0 40204 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1917_
timestamp 28801
transform 1 0 31280 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1918_
timestamp 28801
transform 1 0 35604 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1919_
timestamp 28801
transform -1 0 37996 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1920_
timestamp 28801
transform 1 0 33580 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1921_
timestamp 28801
transform -1 0 41124 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1922_
timestamp 28801
transform 1 0 40572 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1923_
timestamp 28801
transform 1 0 36248 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1924_
timestamp 28801
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1925_
timestamp 28801
transform -1 0 40388 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1926_
timestamp 28801
transform 1 0 36064 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1927_
timestamp 28801
transform -1 0 41952 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1928_
timestamp 28801
transform -1 0 40388 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1929_
timestamp 28801
transform 1 0 35052 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1930_
timestamp 28801
transform 1 0 36616 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1931_
timestamp 28801
transform -1 0 40388 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1932_
timestamp 28801
transform 1 0 36708 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1933_
timestamp 28801
transform -1 0 40480 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1934_
timestamp 28801
transform -1 0 39560 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1935_
timestamp 28801
transform 1 0 31464 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1936_
timestamp 28801
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1937_
timestamp 28801
transform 1 0 40940 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1938_
timestamp 28801
transform -1 0 18400 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1939_
timestamp 28801
transform -1 0 19044 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1940_
timestamp 28801
transform 1 0 17756 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1941_
timestamp 28801
transform 1 0 19228 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1942_
timestamp 28801
transform -1 0 21068 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1943_
timestamp 28801
transform -1 0 21712 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1944_
timestamp 28801
transform 1 0 25024 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1945_
timestamp 28801
transform 1 0 25576 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1946_
timestamp 28801
transform 1 0 25576 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1947_
timestamp 28801
transform 1 0 28428 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1948_
timestamp 28801
transform -1 0 31740 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1949_
timestamp 28801
transform -1 0 33028 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1950_
timestamp 28801
transform -1 0 35328 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1951_
timestamp 28801
transform -1 0 36800 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1952_
timestamp 28801
transform 1 0 34500 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1953_
timestamp 28801
transform 1 0 32660 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1954_
timestamp 28801
transform -1 0 34500 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1955_
timestamp 28801
transform -1 0 15640 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1956_
timestamp 28801
transform 1 0 15272 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1957_
timestamp 28801
transform -1 0 36064 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1958_
timestamp 28801
transform 1 0 30176 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1959_
timestamp 28801
transform -1 0 13524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1960_
timestamp 28801
transform -1 0 7544 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1961_
timestamp 28801
transform 1 0 5336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1962_
timestamp 28801
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1963_
timestamp 28801
transform -1 0 20148 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1964_
timestamp 28801
transform -1 0 20700 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1965_
timestamp 28801
transform -1 0 20424 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1966_
timestamp 28801
transform -1 0 15272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1967_
timestamp 28801
transform 1 0 34776 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1968_
timestamp 28801
transform -1 0 20332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1969_
timestamp 28801
transform 1 0 20240 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1970_
timestamp 28801
transform 1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1971_
timestamp 28801
transform -1 0 6900 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1972_
timestamp 28801
transform -1 0 10488 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1973_
timestamp 28801
transform -1 0 20332 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1974_
timestamp 28801
transform 1 0 2944 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1975_
timestamp 28801
transform 1 0 5060 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1976_
timestamp 28801
transform 1 0 8280 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1977_
timestamp 28801
transform 1 0 5152 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1978_
timestamp 28801
transform 1 0 5704 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _1979_
timestamp 28801
transform -1 0 6164 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1980_
timestamp 28801
transform 1 0 4048 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_4  _1981_
timestamp 28801
transform -1 0 3864 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_2  _1982_
timestamp 28801
transform -1 0 4968 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _1983_
timestamp 28801
transform 1 0 4876 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1984_
timestamp 28801
transform 1 0 5612 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1985_
timestamp 28801
transform -1 0 4600 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1986_
timestamp 28801
transform 1 0 4600 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1987_
timestamp 28801
transform -1 0 4048 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1988_
timestamp 28801
transform 1 0 5704 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1989_
timestamp 28801
transform 1 0 4508 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1990_
timestamp 28801
transform 1 0 3588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1991_
timestamp 28801
transform -1 0 5888 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1992_
timestamp 28801
transform 1 0 3864 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1993_
timestamp 28801
transform -1 0 4416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1994_
timestamp 28801
transform 1 0 5060 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1995_
timestamp 28801
transform 1 0 4416 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1996_
timestamp 28801
transform 1 0 4876 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1997_
timestamp 28801
transform 1 0 4140 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1998_
timestamp 28801
transform 1 0 2116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1999_
timestamp 28801
transform -1 0 5612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _2000_
timestamp 28801
transform 1 0 40480 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2001_
timestamp 28801
transform -1 0 27508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2002_
timestamp 28801
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2003_
timestamp 28801
transform 1 0 32660 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2004_
timestamp 28801
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2005_
timestamp 28801
transform 1 0 26404 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2006_
timestamp 28801
transform 1 0 28612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2007_
timestamp 28801
transform 1 0 22356 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2008_
timestamp 28801
transform 1 0 22080 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2009_
timestamp 28801
transform 1 0 25208 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2010_
timestamp 28801
transform 1 0 27692 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2011_
timestamp 28801
transform -1 0 31004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2012_
timestamp 28801
transform 1 0 31004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2013_
timestamp 28801
transform 1 0 34224 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2014_
timestamp 28801
transform 1 0 38272 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2015_
timestamp 28801
transform 1 0 38640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2016_
timestamp 28801
transform 1 0 37536 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2017_
timestamp 28801
transform 1 0 38180 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2018_
timestamp 28801
transform -1 0 34224 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2019_
timestamp 28801
transform 1 0 35420 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2020_
timestamp 28801
transform -1 0 35880 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2021_
timestamp 28801
transform 1 0 22724 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2022_
timestamp 28801
transform -1 0 21804 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2023_
timestamp 28801
transform 1 0 23276 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2024_
timestamp 28801
transform -1 0 22356 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2025_
timestamp 28801
transform -1 0 20608 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2026_
timestamp 28801
transform -1 0 20608 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2027_
timestamp 28801
transform -1 0 20148 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2028_
timestamp 28801
transform -1 0 21712 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2029_
timestamp 28801
transform 1 0 22448 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2030_
timestamp 28801
transform 1 0 24380 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2031_
timestamp 28801
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2032_
timestamp 28801
transform -1 0 27048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2033_
timestamp 28801
transform 1 0 26956 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2034_
timestamp 28801
transform 1 0 24932 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2035_
timestamp 28801
transform -1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2036_
timestamp 28801
transform 1 0 28152 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2037_
timestamp 28801
transform -1 0 27600 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2038_
timestamp 28801
transform -1 0 30820 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2039_
timestamp 28801
transform -1 0 29348 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2040_
timestamp 28801
transform 1 0 28060 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2041_
timestamp 28801
transform 1 0 28796 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2042_
timestamp 28801
transform 1 0 30268 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2043_
timestamp 28801
transform -1 0 31648 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2044_
timestamp 28801
transform 1 0 32108 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2045_
timestamp 28801
transform -1 0 31280 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2046_
timestamp 28801
transform 1 0 30912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2047_
timestamp 28801
transform 1 0 31464 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _2048_
timestamp 28801
transform 1 0 33212 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _2049_
timestamp 28801
transform -1 0 32844 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2050_
timestamp 28801
transform 1 0 35972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2051_
timestamp 28801
transform 1 0 35972 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2052_
timestamp 28801
transform -1 0 36892 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2053_
timestamp 28801
transform 1 0 34224 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2054_
timestamp 28801
transform 1 0 36708 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2055_
timestamp 28801
transform 1 0 38456 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2056_
timestamp 28801
transform -1 0 36340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _2057_
timestamp 28801
transform 1 0 36156 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2058_
timestamp 28801
transform -1 0 36064 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2059_
timestamp 28801
transform 1 0 35328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2060_
timestamp 28801
transform -1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _2061_
timestamp 28801
transform 1 0 27416 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2062_
timestamp 28801
transform 1 0 13432 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2063_
timestamp 28801
transform -1 0 6992 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2064_
timestamp 28801
transform 1 0 6072 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2065_
timestamp 28801
transform 1 0 6348 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2066_
timestamp 28801
transform 1 0 5888 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2067_
timestamp 28801
transform -1 0 5612 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _2068_
timestamp 28801
transform -1 0 5888 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2069_
timestamp 28801
transform -1 0 5520 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2070_
timestamp 28801
transform -1 0 6164 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2071_
timestamp 28801
transform 1 0 7728 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2072_
timestamp 28801
transform -1 0 8556 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2073_
timestamp 28801
transform 1 0 7360 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _2074_
timestamp 28801
transform -1 0 8832 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2075_
timestamp 28801
transform 1 0 9568 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2076_
timestamp 28801
transform 1 0 8832 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _2077_
timestamp 28801
transform 1 0 8648 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2078_
timestamp 28801
transform -1 0 10212 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2079_
timestamp 28801
transform 1 0 10028 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2080_
timestamp 28801
transform 1 0 9292 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2081_
timestamp 28801
transform -1 0 10948 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2082_
timestamp 28801
transform -1 0 10672 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2083_
timestamp 28801
transform 1 0 9476 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2084_
timestamp 28801
transform -1 0 11776 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2085_
timestamp 28801
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2086_
timestamp 28801
transform -1 0 10580 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2087_
timestamp 28801
transform -1 0 10304 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2088_
timestamp 28801
transform 1 0 8924 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2089_
timestamp 28801
transform -1 0 9016 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _2090_
timestamp 28801
transform 1 0 7544 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2091_
timestamp 28801
transform -1 0 11224 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2092_
timestamp 28801
transform -1 0 7544 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2093_
timestamp 28801
transform 1 0 8372 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2094_
timestamp 28801
transform -1 0 8464 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2095_
timestamp 28801
transform 1 0 10580 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2096_
timestamp 28801
transform -1 0 8740 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2097_
timestamp 28801
transform -1 0 10580 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2098_
timestamp 28801
transform 1 0 6348 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2099_
timestamp 28801
transform -1 0 6256 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _2100_
timestamp 28801
transform -1 0 3772 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2101_
timestamp 28801
transform 1 0 4876 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2102_
timestamp 28801
transform 1 0 5336 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2103_
timestamp 28801
transform 1 0 3956 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2104_
timestamp 28801
transform 1 0 4508 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2105_
timestamp 28801
transform -1 0 4508 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2106_
timestamp 28801
transform -1 0 4968 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2107_
timestamp 28801
transform 1 0 3864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2108_
timestamp 28801
transform 1 0 4508 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2109_
timestamp 28801
transform 1 0 3128 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2110_
timestamp 28801
transform -1 0 5060 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2111_
timestamp 28801
transform 1 0 4968 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2112_
timestamp 28801
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _2113_
timestamp 28801
transform -1 0 4784 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2114_
timestamp 28801
transform 1 0 5612 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2115_
timestamp 28801
transform 1 0 5244 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _2116_
timestamp 28801
transform 1 0 4968 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2117_
timestamp 28801
transform 1 0 5428 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2118_
timestamp 28801
transform 1 0 4232 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2119_
timestamp 28801
transform 1 0 4692 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2120_
timestamp 28801
transform -1 0 4692 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2121_
timestamp 28801
transform 1 0 6164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2122_
timestamp 28801
transform 1 0 4784 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2123_
timestamp 28801
transform -1 0 4784 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2124_
timestamp 28801
transform -1 0 5428 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _2125_
timestamp 28801
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2126_
timestamp 28801
transform -1 0 4416 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2127_
timestamp 28801
transform 1 0 2392 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2128_
timestamp 28801
transform -1 0 2392 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2129_
timestamp 28801
transform 1 0 2208 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2130_
timestamp 28801
transform 1 0 2392 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2131_
timestamp 28801
transform 1 0 1564 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2132_
timestamp 28801
transform 1 0 3220 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2133_
timestamp 28801
transform 1 0 2852 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2134_
timestamp 28801
transform 1 0 2024 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2135_
timestamp 28801
transform -1 0 2852 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2136_
timestamp 28801
transform 1 0 1748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2137_
timestamp 28801
transform 1 0 3772 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2138_
timestamp 28801
transform 1 0 2024 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2139_
timestamp 28801
transform -1 0 4416 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2140_
timestamp 28801
transform -1 0 3496 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2141_
timestamp 28801
transform 1 0 5612 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2142_
timestamp 28801
transform 1 0 5888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2143_
timestamp 28801
transform 1 0 5244 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2144_
timestamp 28801
transform 1 0 6256 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2145_
timestamp 28801
transform -1 0 5428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2146_
timestamp 28801
transform -1 0 6808 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2147_
timestamp 28801
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2148_
timestamp 28801
transform -1 0 6256 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2149_
timestamp 28801
transform -1 0 6900 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2150_
timestamp 28801
transform -1 0 5152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2151_
timestamp 28801
transform 1 0 5152 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2152_
timestamp 28801
transform -1 0 5244 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2153_
timestamp 28801
transform 1 0 5060 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2154_
timestamp 28801
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2155_
timestamp 28801
transform -1 0 6164 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _2156_
timestamp 28801
transform 1 0 4600 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2157_
timestamp 28801
transform -1 0 6440 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2158_
timestamp 28801
transform -1 0 7268 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2159_
timestamp 28801
transform -1 0 5796 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2160_
timestamp 28801
transform 1 0 5704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2161_
timestamp 28801
transform 1 0 4416 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2162_
timestamp 28801
transform 1 0 6624 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2163_
timestamp 28801
transform 1 0 6900 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2164_
timestamp 28801
transform -1 0 7912 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2165_
timestamp 28801
transform 1 0 6900 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _2166_
timestamp 28801
transform 1 0 19228 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2167_
timestamp 28801
transform 1 0 14628 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2168_
timestamp 28801
transform 1 0 14260 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _2169_
timestamp 28801
transform 1 0 20056 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _2170_
timestamp 28801
transform 1 0 20792 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _2171_
timestamp 28801
transform -1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2172_
timestamp 28801
transform -1 0 16100 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2173_
timestamp 28801
transform 1 0 18400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2174_
timestamp 28801
transform -1 0 18400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2175_
timestamp 28801
transform -1 0 18584 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2176_
timestamp 28801
transform -1 0 18584 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2177_
timestamp 28801
transform -1 0 17756 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2178_
timestamp 28801
transform -1 0 16192 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2179_
timestamp 28801
transform -1 0 16836 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2180_
timestamp 28801
transform 1 0 12512 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2181_
timestamp 28801
transform -1 0 12696 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2182_
timestamp 28801
transform -1 0 13340 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2183_
timestamp 28801
transform 1 0 13524 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _2184_
timestamp 28801
transform 1 0 19596 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _2185_
timestamp 28801
transform -1 0 19596 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2186_
timestamp 28801
transform 1 0 14352 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2187_
timestamp 28801
transform 1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2188_
timestamp 28801
transform 1 0 14996 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2189_
timestamp 28801
transform -1 0 13984 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2190_
timestamp 28801
transform -1 0 14996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _2191_
timestamp 28801
transform 1 0 14352 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2192_
timestamp 28801
transform 1 0 14628 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2193_
timestamp 28801
transform -1 0 15364 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2194_
timestamp 28801
transform 1 0 15824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2195_
timestamp 28801
transform 1 0 15088 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2196_
timestamp 28801
transform -1 0 15732 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2197_
timestamp 28801
transform 1 0 14628 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _2198_
timestamp 28801
transform -1 0 5980 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2199_
timestamp 28801
transform 1 0 6624 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2200_
timestamp 28801
transform 1 0 3956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2201_
timestamp 28801
transform 1 0 6624 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2202_
timestamp 28801
transform 1 0 4508 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2203_
timestamp 28801
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2204_
timestamp 28801
transform -1 0 6532 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2205_
timestamp 28801
transform -1 0 6624 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2206_
timestamp 28801
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2207_
timestamp 28801
transform -1 0 11408 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2208_
timestamp 28801
transform 1 0 9016 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _2209_
timestamp 28801
transform -1 0 6992 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2210_
timestamp 28801
transform 1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2211_
timestamp 28801
transform -1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2212_
timestamp 28801
transform 1 0 6440 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2213_
timestamp 28801
transform 1 0 8372 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2214_
timestamp 28801
transform -1 0 12144 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2215_
timestamp 28801
transform -1 0 8648 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2216_
timestamp 28801
transform -1 0 7360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2217_
timestamp 28801
transform -1 0 7820 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2218_
timestamp 28801
transform 1 0 12328 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2219_
timestamp 28801
transform -1 0 12880 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2220_
timestamp 28801
transform -1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2221_
timestamp 28801
transform 1 0 4140 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2222_
timestamp 28801
transform 1 0 5520 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _2223_
timestamp 28801
transform 1 0 3772 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2224_
timestamp 28801
transform -1 0 6256 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _2225_
timestamp 28801
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2226_
timestamp 28801
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _2227_
timestamp 28801
transform 1 0 6440 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2228_
timestamp 28801
transform 1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _2229_
timestamp 28801
transform -1 0 12328 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2230_
timestamp 28801
transform -1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _2231_
timestamp 28801
transform -1 0 12052 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2232_
timestamp 28801
transform -1 0 9752 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2233_
timestamp 28801
transform 1 0 8188 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2234_
timestamp 28801
transform 1 0 7360 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2235_
timestamp 28801
transform -1 0 7452 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2236_
timestamp 28801
transform -1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _2237_
timestamp 28801
transform -1 0 5336 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2238_
timestamp 28801
transform -1 0 5428 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2239_
timestamp 28801
transform -1 0 6164 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2240_
timestamp 28801
transform -1 0 14444 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2241_
timestamp 28801
transform 1 0 12236 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2242_
timestamp 28801
transform 1 0 30268 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2243_
timestamp 28801
transform 1 0 16100 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2244_
timestamp 28801
transform 1 0 16192 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2245_
timestamp 28801
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _2246_
timestamp 28801
transform 1 0 9292 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _2247_
timestamp 28801
transform -1 0 12696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2248_
timestamp 28801
transform 1 0 9844 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2249_
timestamp 28801
transform 1 0 6348 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2250_
timestamp 28801
transform -1 0 6256 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _2251_
timestamp 28801
transform -1 0 11960 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2252_
timestamp 28801
transform -1 0 11040 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2253_
timestamp 28801
transform 1 0 10580 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2254_
timestamp 28801
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2255_
timestamp 28801
transform -1 0 7820 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2256_
timestamp 28801
transform 1 0 10488 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _2257_
timestamp 28801
transform -1 0 12880 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2258_
timestamp 28801
transform -1 0 11040 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _2259_
timestamp 28801
transform -1 0 11408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _2260_
timestamp 28801
transform 1 0 9016 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2261_
timestamp 28801
transform -1 0 10396 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2262_
timestamp 28801
transform -1 0 7268 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2263_
timestamp 28801
transform 1 0 8096 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2264_
timestamp 28801
transform -1 0 9108 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2265_
timestamp 28801
transform 1 0 8372 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2266_
timestamp 28801
transform 1 0 9200 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2267_
timestamp 28801
transform 1 0 9568 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2268_
timestamp 28801
transform -1 0 9752 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2269_
timestamp 28801
transform -1 0 10948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2270_
timestamp 28801
transform 1 0 11316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2271_
timestamp 28801
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2272_
timestamp 28801
transform 1 0 11684 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2273_
timestamp 28801
transform 1 0 12328 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2274_
timestamp 28801
transform 1 0 12972 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2275_
timestamp 28801
transform -1 0 12328 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2276_
timestamp 28801
transform -1 0 13892 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2277_
timestamp 28801
transform 1 0 13340 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2278_
timestamp 28801
transform -1 0 12972 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2279_
timestamp 28801
transform 1 0 12420 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2280_
timestamp 28801
transform 1 0 12144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2281_
timestamp 28801
transform 1 0 12880 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2282_
timestamp 28801
transform -1 0 13064 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2283_
timestamp 28801
transform 1 0 13064 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2284_
timestamp 28801
transform 1 0 12420 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2285_
timestamp 28801
transform -1 0 12788 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2286_
timestamp 28801
transform 1 0 11500 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2287_
timestamp 28801
transform 1 0 10304 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2288_
timestamp 28801
transform -1 0 8832 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2289_
timestamp 28801
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2290_
timestamp 28801
transform -1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2291_
timestamp 28801
transform 1 0 8004 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2292_
timestamp 28801
transform 1 0 8924 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2293_
timestamp 28801
transform -1 0 9016 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2294_
timestamp 28801
transform 1 0 8464 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2295_
timestamp 28801
transform -1 0 8464 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2296_
timestamp 28801
transform -1 0 8096 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2297_
timestamp 28801
transform -1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2298_
timestamp 28801
transform -1 0 7636 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2299_
timestamp 28801
transform 1 0 3588 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2300_
timestamp 28801
transform 1 0 4324 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2301_
timestamp 28801
transform 1 0 4508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2302_
timestamp 28801
transform -1 0 5244 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2303_
timestamp 28801
transform -1 0 3496 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2304_
timestamp 28801
transform -1 0 4232 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2305_
timestamp 28801
transform -1 0 2208 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2306_
timestamp 28801
transform -1 0 3680 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2307_
timestamp 28801
transform 1 0 7176 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _2308_
timestamp 28801
transform -1 0 7820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2309_
timestamp 28801
transform -1 0 7820 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _2310_
timestamp 28801
transform -1 0 8096 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2311_
timestamp 28801
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2312_
timestamp 28801
transform 1 0 9660 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2313_
timestamp 28801
transform 1 0 9292 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2314_
timestamp 28801
transform -1 0 9292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2315_
timestamp 28801
transform 1 0 9292 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a311oi_4  _2316_
timestamp 28801
transform 1 0 6164 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _2317_
timestamp 28801
transform 1 0 6532 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2318_
timestamp 28801
transform 1 0 7176 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2319_
timestamp 28801
transform 1 0 6808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2320_
timestamp 28801
transform 1 0 7084 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2321_
timestamp 28801
transform 1 0 7084 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2322_
timestamp 28801
transform 1 0 7544 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2323_
timestamp 28801
transform 1 0 7636 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2324_
timestamp 28801
transform 1 0 7636 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2325_
timestamp 28801
transform 1 0 7728 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2326_
timestamp 28801
transform 1 0 8188 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2327_
timestamp 28801
transform 1 0 8832 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2328_
timestamp 28801
transform 1 0 8372 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2329_
timestamp 28801
transform 1 0 8924 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2330_
timestamp 28801
transform 1 0 8188 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2331_
timestamp 28801
transform 1 0 8924 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2332_
timestamp 28801
transform -1 0 8464 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2333_
timestamp 28801
transform 1 0 19964 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2334_
timestamp 28801
transform 1 0 18492 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2335_
timestamp 28801
transform -1 0 24380 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2336_
timestamp 28801
transform -1 0 22540 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2337_
timestamp 28801
transform 1 0 24104 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2338_
timestamp 28801
transform 1 0 25116 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2339_
timestamp 28801
transform -1 0 30176 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2340_
timestamp 28801
transform -1 0 31188 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2341_
timestamp 28801
transform 1 0 29348 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2342_
timestamp 28801
transform -1 0 32016 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2343_
timestamp 28801
transform 1 0 32844 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2344_
timestamp 28801
transform -1 0 35328 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2345_
timestamp 28801
transform 1 0 36432 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2346_
timestamp 28801
transform 1 0 37076 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2347_
timestamp 28801
transform -1 0 39284 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2348_
timestamp 28801
transform 1 0 5060 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2349_
timestamp 28801
transform -1 0 5060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2350_
timestamp 28801
transform 1 0 5244 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2351_
timestamp 28801
transform -1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2352_
timestamp 28801
transform 1 0 6072 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2353_
timestamp 28801
transform 1 0 5796 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2354_
timestamp 28801
transform -1 0 8004 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2355_
timestamp 28801
transform -1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2356_
timestamp 28801
transform 1 0 6532 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2357_
timestamp 28801
transform -1 0 6072 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2358_
timestamp 28801
transform -1 0 5704 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2359_
timestamp 28801
transform -1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2360_
timestamp 28801
transform 1 0 4600 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2361_
timestamp 28801
transform -1 0 4968 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2362_
timestamp 28801
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2363_
timestamp 28801
transform 1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2364_
timestamp 28801
transform -1 0 4232 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2365_
timestamp 28801
transform 1 0 2392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2366_
timestamp 28801
transform -1 0 2208 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2367_
timestamp 28801
transform -1 0 3128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2368_
timestamp 28801
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2369_
timestamp 28801
transform 1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2370_
timestamp 28801
transform -1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2371_
timestamp 28801
transform 1 0 2944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2372_
timestamp 28801
transform -1 0 3680 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2373_
timestamp 28801
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2374_
timestamp 28801
transform 1 0 1564 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2375_
timestamp 28801
transform -1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2376_
timestamp 28801
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2377_
timestamp 28801
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2378_
timestamp 28801
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2379_
timestamp 28801
transform -1 0 3588 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2380_
timestamp 28801
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2381_
timestamp 28801
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2382_
timestamp 28801
transform -1 0 3772 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2383_
timestamp 28801
transform 1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2384_
timestamp 28801
transform -1 0 4416 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2385_
timestamp 28801
transform -1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _2386_
timestamp 28801
transform -1 0 5888 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2387_
timestamp 28801
transform -1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2388_
timestamp 28801
transform -1 0 7360 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2389_
timestamp 28801
transform 1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2390_
timestamp 28801
transform 1 0 6348 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2391_
timestamp 28801
transform -1 0 7728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2392_
timestamp 28801
transform -1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2393_
timestamp 28801
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2394_
timestamp 28801
transform -1 0 8648 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2395_
timestamp 28801
transform 1 0 8648 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2396_
timestamp 28801
transform -1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2397_
timestamp 28801
transform 1 0 8372 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2398_
timestamp 28801
transform -1 0 9568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2399_
timestamp 28801
transform 1 0 9752 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2400_
timestamp 28801
transform -1 0 9108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2401_
timestamp 28801
transform -1 0 9936 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2402_
timestamp 28801
transform -1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2403_
timestamp 28801
transform 1 0 9936 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2404_
timestamp 28801
transform 1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2405_
timestamp 28801
transform 1 0 10396 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2406_
timestamp 28801
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2407_
timestamp 28801
transform -1 0 13340 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2408_
timestamp 28801
transform 1 0 12788 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2409_
timestamp 28801
transform -1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2410_
timestamp 28801
transform -1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2411_
timestamp 28801
transform -1 0 12788 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2412_
timestamp 28801
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _2413_
timestamp 28801
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2414_
timestamp 28801
transform -1 0 11960 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _2415_
timestamp 28801
transform 1 0 10580 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2416_
timestamp 28801
transform -1 0 8372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _2417_
timestamp 28801
transform -1 0 9108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2418_
timestamp 28801
transform -1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2419_
timestamp 28801
transform 1 0 8372 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2420_
timestamp 28801
transform -1 0 13984 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2421_
timestamp 28801
transform 1 0 13340 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2422_
timestamp 28801
transform -1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2423_
timestamp 28801
transform 1 0 13064 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2424_
timestamp 28801
transform 1 0 13524 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2425_
timestamp 28801
transform 1 0 14076 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2426_
timestamp 28801
transform -1 0 12972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2427_
timestamp 28801
transform -1 0 13340 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2428_
timestamp 28801
transform -1 0 12696 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2429_
timestamp 28801
transform -1 0 12328 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2430_
timestamp 28801
transform 1 0 13340 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _2431_
timestamp 28801
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2432_
timestamp 28801
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2433_
timestamp 28801
transform -1 0 13524 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2434_
timestamp 28801
transform -1 0 12972 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2435_
timestamp 28801
transform 1 0 12328 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2436_
timestamp 28801
transform -1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2437_
timestamp 28801
transform 1 0 11868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _2438_
timestamp 28801
transform -1 0 11684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2439_
timestamp 28801
transform -1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2440_
timestamp 28801
transform -1 0 11684 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _2441_
timestamp 28801
transform 1 0 10028 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2442_
timestamp 28801
transform 1 0 10488 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _2443_
timestamp 28801
transform 1 0 20424 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2444_
timestamp 28801
transform 1 0 6624 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2445_
timestamp 28801
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2446_
timestamp 28801
transform 1 0 9476 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2447_
timestamp 28801
transform 1 0 9752 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2448_
timestamp 28801
transform 1 0 11960 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2449_
timestamp 28801
transform 1 0 11868 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2450_
timestamp 28801
transform -1 0 14536 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2451_
timestamp 28801
transform -1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2452_
timestamp 28801
transform -1 0 14444 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2453_
timestamp 28801
transform -1 0 14536 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2454_
timestamp 28801
transform -1 0 14996 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2455_
timestamp 28801
transform 1 0 10856 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2456_
timestamp 28801
transform 1 0 8924 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2457_
timestamp 28801
transform 1 0 8648 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2458_
timestamp 28801
transform 1 0 7820 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2459_
timestamp 28801
transform 1 0 7084 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2460_
timestamp 28801
transform -1 0 5704 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2461_
timestamp 28801
transform 1 0 2208 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2462_
timestamp 28801
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2463_
timestamp 28801
transform 1 0 1748 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _2464_
timestamp 28801
transform 1 0 4324 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2465_
timestamp 28801
transform 1 0 6348 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2466_
timestamp 28801
transform 1 0 3864 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _2467_
timestamp 28801
transform 1 0 3404 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2468_
timestamp 28801
transform 1 0 6624 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2469_
timestamp 28801
transform 1 0 6716 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2470_
timestamp 28801
transform 1 0 8924 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2471_
timestamp 28801
transform 1 0 9108 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2472_
timestamp 28801
transform 1 0 9200 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2473_
timestamp 28801
transform 1 0 9568 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2474_
timestamp 28801
transform 1 0 6716 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2475_
timestamp 28801
transform -1 0 8740 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2476_
timestamp 28801
transform -1 0 10764 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2477_
timestamp 28801
transform 1 0 5244 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2478_
timestamp 28801
transform 1 0 3772 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2479_
timestamp 28801
transform 1 0 2668 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2480_
timestamp 28801
transform -1 0 4968 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2481_
timestamp 28801
transform -1 0 7544 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2482_
timestamp 28801
transform 1 0 3956 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2483_
timestamp 28801
transform -1 0 3220 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2484_
timestamp 28801
transform 1 0 1380 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2485_
timestamp 28801
transform 1 0 1380 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2486_
timestamp 28801
transform 1 0 1932 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2487_
timestamp 28801
transform 1 0 8096 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2488_
timestamp 28801
transform 1 0 9936 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2489_
timestamp 28801
transform 1 0 10120 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2490_
timestamp 28801
transform 1 0 9936 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2491_
timestamp 28801
transform -1 0 9016 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2492_
timestamp 28801
transform -1 0 10856 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2493_
timestamp 28801
transform -1 0 10856 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2494_
timestamp 28801
transform -1 0 10488 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _2495_
timestamp 28801
transform -1 0 21436 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2496_
timestamp 28801
transform 1 0 19320 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2497_
timestamp 28801
transform -1 0 23644 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2498_
timestamp 28801
transform 1 0 21436 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2499_
timestamp 28801
transform -1 0 26220 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2500_
timestamp 28801
transform -1 0 27140 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2501_
timestamp 28801
transform -1 0 28796 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2502_
timestamp 28801
transform 1 0 29532 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2503_
timestamp 28801
transform -1 0 31372 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2504_
timestamp 28801
transform 1 0 31188 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2505_
timestamp 28801
transform 1 0 33948 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2506_
timestamp 28801
transform -1 0 35052 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2507_
timestamp 28801
transform -1 0 37720 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2508_
timestamp 28801
transform -1 0 39192 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2509_
timestamp 28801
transform 1 0 38640 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2510_
timestamp 28801
transform 1 0 1380 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2511_
timestamp 28801
transform 1 0 1380 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2512_
timestamp 28801
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2513_
timestamp 28801
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2514_
timestamp 28801
transform -1 0 7544 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2515_
timestamp 28801
transform 1 0 3036 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2516_
timestamp 28801
transform -1 0 8372 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2517_
timestamp 28801
transform 1 0 4784 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2518_
timestamp 28801
transform 1 0 3772 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2519_
timestamp 28801
transform 1 0 1472 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2520_
timestamp 28801
transform 1 0 1472 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2521_
timestamp 28801
transform 1 0 1564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2522_
timestamp 28801
transform 1 0 1380 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2523_
timestamp 28801
transform 1 0 2944 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2524_
timestamp 28801
transform 1 0 1380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2525_
timestamp 28801
transform 1 0 1380 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2526_
timestamp 28801
transform 1 0 1748 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2527_
timestamp 28801
transform 1 0 3772 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2528_
timestamp 28801
transform 1 0 4140 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2529_
timestamp 28801
transform 1 0 5888 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2530_
timestamp 28801
transform 1 0 6808 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2531_
timestamp 28801
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2532_
timestamp 28801
transform -1 0 11132 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2533_
timestamp 28801
transform -1 0 9292 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2534_
timestamp 28801
transform 1 0 9476 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2535_
timestamp 28801
transform -1 0 15364 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2536_
timestamp 28801
transform -1 0 13892 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2537_
timestamp 28801
transform 1 0 10120 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2538_
timestamp 28801
transform 1 0 8924 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2539_
timestamp 28801
transform -1 0 15916 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2540_
timestamp 28801
transform -1 0 15824 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2541_
timestamp 28801
transform 1 0 11500 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2542_
timestamp 28801
transform -1 0 15364 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2543_
timestamp 28801
transform 1 0 11868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2544_
timestamp 28801
transform 1 0 9568 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2545_
timestamp 28801
transform 1 0 9384 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2546_
timestamp 28801
transform -1 0 3220 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2547_
timestamp 28801
transform -1 0 3220 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2548_
timestamp 28801
transform -1 0 3220 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2549_
timestamp 28801
transform 1 0 6348 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2550_
timestamp 28801
transform 1 0 1748 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2551_
timestamp 28801
transform 1 0 2668 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2552_
timestamp 28801
transform 1 0 2576 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2553_
timestamp 28801
transform 1 0 2668 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2554_
timestamp 28801
transform 1 0 16376 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2555_
timestamp 28801
transform -1 0 19596 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2556_
timestamp 28801
transform 1 0 20884 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2557_
timestamp 28801
transform -1 0 25024 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2558_
timestamp 28801
transform 1 0 24380 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2559_
timestamp 28801
transform 1 0 25760 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2560_
timestamp 28801
transform -1 0 28612 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2561_
timestamp 28801
transform 1 0 28244 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2562_
timestamp 28801
transform 1 0 29900 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2563_
timestamp 28801
transform 1 0 31648 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2564_
timestamp 28801
transform 1 0 37260 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2565_
timestamp 28801
transform 1 0 35972 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2566_
timestamp 28801
transform 1 0 35052 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2567_
timestamp 28801
transform -1 0 34960 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2568_
timestamp 28801
transform 1 0 32016 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2569_
timestamp 28801
transform 1 0 17204 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2570_
timestamp 28801
transform 1 0 18492 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2571_
timestamp 28801
transform -1 0 22172 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2572_
timestamp 28801
transform 1 0 22172 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2573_
timestamp 28801
transform 1 0 24472 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2574_
timestamp 28801
transform 1 0 24288 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2575_
timestamp 28801
transform 1 0 26864 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2576_
timestamp 28801
transform 1 0 27600 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2577_
timestamp 28801
transform 1 0 30084 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2578_
timestamp 28801
transform -1 0 34592 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2579_
timestamp 28801
transform 1 0 36984 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2580_
timestamp 28801
transform 1 0 37260 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2581_
timestamp 28801
transform 1 0 36248 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2582_
timestamp 28801
transform -1 0 35236 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2583_
timestamp 28801
transform 1 0 29992 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2584_
timestamp 28801
transform 1 0 11500 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2585_
timestamp 28801
transform 1 0 13340 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2586_
timestamp 28801
transform 1 0 12052 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2587_
timestamp 28801
transform 1 0 11960 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2588_
timestamp 28801
transform 1 0 9108 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2589_
timestamp 28801
transform 1 0 18400 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2590_
timestamp 28801
transform 1 0 17296 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2591_
timestamp 28801
transform 1 0 20424 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2592_
timestamp 28801
transform -1 0 23644 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2593_
timestamp 28801
transform 1 0 23184 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2594_
timestamp 28801
transform 1 0 23828 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2595_
timestamp 28801
transform 1 0 26220 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2596_
timestamp 28801
transform 1 0 28152 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2597_
timestamp 28801
transform -1 0 30084 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2598_
timestamp 28801
transform 1 0 31372 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2599_
timestamp 28801
transform 1 0 32108 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2600_
timestamp 28801
transform 1 0 32752 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2601_
timestamp 28801
transform 1 0 35144 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2602_
timestamp 28801
transform 1 0 35604 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2603_
timestamp 28801
transform 1 0 37904 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2604_
timestamp 28801
transform 1 0 14444 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2605_
timestamp 28801
transform 1 0 15456 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2606_
timestamp 28801
transform 1 0 17664 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2607_
timestamp 28801
transform 1 0 18124 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2608_
timestamp 28801
transform 1 0 19872 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2609_
timestamp 28801
transform 1 0 22080 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2610_
timestamp 28801
transform 1 0 23828 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2611_
timestamp 28801
transform 1 0 25300 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2612_
timestamp 28801
transform 1 0 26588 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2613_
timestamp 28801
transform 1 0 27968 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2614_
timestamp 28801
transform 1 0 29808 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2615_
timestamp 28801
transform 1 0 32568 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2616_
timestamp 28801
transform 1 0 35052 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2617_
timestamp 28801
transform 1 0 34960 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2618_
timestamp 28801
transform 1 0 35236 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2619_
timestamp 28801
transform 1 0 35512 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2620_
timestamp 28801
transform 1 0 30176 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2621_
timestamp 28801
transform 1 0 16652 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2622_
timestamp 28801
transform 1 0 18492 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2623_
timestamp 28801
transform 1 0 16836 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2624_
timestamp 28801
transform 1 0 20608 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2625_
timestamp 28801
transform -1 0 23736 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2626_
timestamp 28801
transform 1 0 24104 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2627_
timestamp 28801
transform 1 0 24932 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2628_
timestamp 28801
transform -1 0 28980 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2629_
timestamp 28801
transform 1 0 28704 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2630_
timestamp 28801
transform 1 0 30820 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2631_
timestamp 28801
transform 1 0 35236 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2632_
timestamp 28801
transform 1 0 39836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2633_
timestamp 28801
transform 1 0 40204 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2634_
timestamp 28801
transform 1 0 40112 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2635_
timestamp 28801
transform 1 0 38916 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2636_
timestamp 28801
transform -1 0 34316 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2637_
timestamp 28801
transform -1 0 17112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2638_
timestamp 28801
transform 1 0 15916 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2639_
timestamp 28801
transform 1 0 15640 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2640_
timestamp 28801
transform -1 0 22356 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2641_
timestamp 28801
transform 1 0 21988 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2642_
timestamp 28801
transform 1 0 23092 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2643_
timestamp 28801
transform 1 0 25208 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2644_
timestamp 28801
transform 1 0 26956 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2645_
timestamp 28801
transform 1 0 28336 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2646_
timestamp 28801
transform -1 0 33948 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2647_
timestamp 28801
transform -1 0 38916 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2648_
timestamp 28801
transform 1 0 39928 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2649_
timestamp 28801
transform 1 0 40388 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2650_
timestamp 28801
transform 1 0 37168 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2651_
timestamp 28801
transform 1 0 40388 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2652_
timestamp 28801
transform 1 0 31924 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2653_
timestamp 28801
transform 1 0 19228 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2654_
timestamp 28801
transform 1 0 18308 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2655_
timestamp 28801
transform -1 0 22172 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2656_
timestamp 28801
transform 1 0 22356 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2657_
timestamp 28801
transform 1 0 24196 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2658_
timestamp 28801
transform 1 0 24932 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2659_
timestamp 28801
transform 1 0 26220 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2660_
timestamp 28801
transform -1 0 29808 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2661_
timestamp 28801
transform 1 0 29532 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2662_
timestamp 28801
transform -1 0 32660 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2663_
timestamp 28801
transform 1 0 31372 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2664_
timestamp 28801
transform 1 0 33580 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2665_
timestamp 28801
transform 1 0 35788 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2666_
timestamp 28801
transform 1 0 34500 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2667_
timestamp 28801
transform 1 0 32660 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2668_
timestamp 28801
transform 1 0 16652 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2669_
timestamp 28801
transform 1 0 17848 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2670_
timestamp 28801
transform 1 0 19872 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2671_
timestamp 28801
transform 1 0 20240 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2672_
timestamp 28801
transform 1 0 22448 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2673_
timestamp 28801
transform 1 0 23828 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2674_
timestamp 28801
transform 1 0 29532 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2675_
timestamp 28801
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2676_
timestamp 28801
transform -1 0 31740 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2677_
timestamp 28801
transform 1 0 33488 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2678_
timestamp 28801
transform 1 0 37536 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2679_
timestamp 28801
transform 1 0 37628 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2680_
timestamp 28801
transform 1 0 37444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2681_
timestamp 28801
transform -1 0 39192 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2682_
timestamp 28801
transform -1 0 36800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 28801
transform 1 0 14996 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2684_
timestamp 28801
transform 1 0 15732 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2685_
timestamp 28801
transform 1 0 27876 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 28801
transform 1 0 27324 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 28801
transform 1 0 16652 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 28801
transform -1 0 31464 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2689_
timestamp 28801
transform 1 0 15640 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 28801
transform 1 0 17296 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2691_
timestamp 28801
transform 1 0 18768 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2692_
timestamp 28801
transform 1 0 20608 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 28801
transform 1 0 22172 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 28801
transform 1 0 25024 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 28801
transform 1 0 26220 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 28801
transform 1 0 27232 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2697_
timestamp 28801
transform 1 0 28520 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2698_
timestamp 28801
transform -1 0 23736 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2699_
timestamp 28801
transform 1 0 32108 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2700_
timestamp 28801
transform 1 0 35328 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 28801
transform 1 0 33948 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 28801
transform 1 0 34960 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2703_
timestamp 28801
transform 1 0 34776 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2704_
timestamp 28801
transform 1 0 32108 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2705_
timestamp 28801
transform 1 0 17296 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2706_
timestamp 28801
transform 1 0 14720 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2707_
timestamp 28801
transform 1 0 15364 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2708_
timestamp 28801
transform 1 0 19228 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2709_
timestamp 28801
transform 1 0 21712 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2710_
timestamp 28801
transform 1 0 23276 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2711_
timestamp 28801
transform 1 0 24288 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2712_
timestamp 28801
transform 1 0 26864 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2713_
timestamp 28801
transform 1 0 29532 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2714_
timestamp 28801
transform 1 0 32108 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2715_
timestamp 28801
transform -1 0 39744 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2716_
timestamp 28801
transform 1 0 40388 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2717_
timestamp 28801
transform 1 0 39560 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2718_
timestamp 28801
transform 1 0 37260 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2719_
timestamp 28801
transform 1 0 32016 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2720_
timestamp 28801
transform 1 0 29532 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2721_
timestamp 28801
transform 1 0 14812 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2722_
timestamp 28801
transform 1 0 16836 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2723_
timestamp 28801
transform 1 0 19412 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2724_
timestamp 28801
transform 1 0 22172 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2725_
timestamp 28801
transform 1 0 24380 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2726_
timestamp 28801
transform 1 0 24748 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2727_
timestamp 28801
transform 1 0 27048 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2728_
timestamp 28801
transform 1 0 29716 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2729_
timestamp 28801
transform -1 0 35788 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2730_
timestamp 28801
transform 1 0 35972 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2731_
timestamp 28801
transform 1 0 39192 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2732_
timestamp 28801
transform 1 0 40388 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2733_
timestamp 28801
transform 1 0 37260 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2734_
timestamp 28801
transform 1 0 32108 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2735_
timestamp 28801
transform 1 0 29716 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2736_
timestamp 28801
transform 1 0 12880 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2737_
timestamp 28801
transform 1 0 15364 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2738_
timestamp 28801
transform 1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2739_
timestamp 28801
transform 1 0 20884 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2740_
timestamp 28801
transform 1 0 22540 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2741_
timestamp 28801
transform 1 0 23460 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2742_
timestamp 28801
transform 1 0 25300 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2743_
timestamp 28801
transform 1 0 26956 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2744_
timestamp 28801
transform 1 0 28428 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2745_
timestamp 28801
transform 1 0 31004 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2746_
timestamp 28801
transform 1 0 37260 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2747_
timestamp 28801
transform 1 0 38824 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2748_
timestamp 28801
transform 1 0 39928 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2749_
timestamp 28801
transform 1 0 37260 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2750_
timestamp 28801
transform 1 0 39836 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2751_
timestamp 28801
transform 1 0 30452 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2752_
timestamp 28801
transform 1 0 14444 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2753_
timestamp 28801
transform -1 0 13892 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2754_
timestamp 28801
transform 1 0 11960 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2755_
timestamp 28801
transform 1 0 11592 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2756_
timestamp 28801
transform 1 0 11776 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2757_
timestamp 28801
transform 1 0 10948 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2758_
timestamp 28801
transform -1 0 16560 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2759_
timestamp 28801
transform -1 0 18676 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2760_
timestamp 28801
transform 1 0 19872 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2761_
timestamp 28801
transform -1 0 23644 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2762_
timestamp 28801
transform 1 0 24380 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2763_
timestamp 28801
transform 1 0 25300 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2764_
timestamp 28801
transform 1 0 27324 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2765_
timestamp 28801
transform 1 0 28428 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2766_
timestamp 28801
transform 1 0 31096 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2767_
timestamp 28801
transform -1 0 39376 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2768_
timestamp 28801
transform 1 0 39652 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2769_
timestamp 28801
transform 1 0 40296 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2770_
timestamp 28801
transform 1 0 37076 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2771_
timestamp 28801
transform 1 0 33028 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2772_
timestamp 28801
transform 1 0 29716 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2773_
timestamp 28801
transform 1 0 14076 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2774_
timestamp 28801
transform -1 0 18124 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2775_
timestamp 28801
transform 1 0 17112 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2776_
timestamp 28801
transform 1 0 19964 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2777_
timestamp 28801
transform -1 0 23736 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2778_
timestamp 28801
transform 1 0 24380 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2779_
timestamp 28801
transform 1 0 25852 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2780_
timestamp 28801
transform 1 0 27140 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2781_
timestamp 28801
transform 1 0 28796 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2782_
timestamp 28801
transform 1 0 34500 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2783_
timestamp 28801
transform 1 0 37812 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2784_
timestamp 28801
transform 1 0 39652 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2785_
timestamp 28801
transform 1 0 39928 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2786_
timestamp 28801
transform 1 0 37260 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2787_
timestamp 28801
transform 1 0 32752 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2788_
timestamp 28801
transform -1 0 32660 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2789_
timestamp 28801
transform -1 0 16192 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2790_
timestamp 28801
transform 1 0 12512 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2791_
timestamp 28801
transform 1 0 11592 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2792_
timestamp 28801
transform 1 0 11224 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2793_
timestamp 28801
transform 1 0 11592 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2794_
timestamp 28801
transform 1 0 9476 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2795_
timestamp 28801
transform 1 0 10304 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2796_
timestamp 28801
transform 1 0 10856 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2797_
timestamp 28801
transform 1 0 9200 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2798_
timestamp 28801
transform 1 0 14260 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2799_
timestamp 28801
transform 1 0 14720 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2800_
timestamp 28801
transform -1 0 13984 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2801_
timestamp 28801
transform 1 0 19228 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2802_
timestamp 28801
transform 1 0 19320 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2803_
timestamp 28801
transform 1 0 21160 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2804_
timestamp 28801
transform -1 0 24380 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2805_
timestamp 28801
transform 1 0 40388 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2806_
timestamp 28801
transform 1 0 37904 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2807_
timestamp 28801
transform 1 0 39468 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2808_
timestamp 28801
transform 1 0 40112 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2809_
timestamp 28801
transform 1 0 37260 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2810_
timestamp 28801
transform 1 0 40388 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2811_
timestamp 28801
transform 1 0 40388 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2812_
timestamp 28801
transform 1 0 40388 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2813_
timestamp 28801
transform 1 0 40388 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2814_
timestamp 28801
transform 1 0 38824 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2815_
timestamp 28801
transform 1 0 40388 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2816_
timestamp 28801
transform 1 0 17848 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2817_
timestamp 28801
transform 1 0 12696 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2818_
timestamp 28801
transform 1 0 15364 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2819_
timestamp 28801
transform 1 0 15548 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2820_
timestamp 28801
transform 1 0 14904 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _2821_
timestamp 28801
transform 1 0 18676 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2822_
timestamp 28801
transform 1 0 18860 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2823_
timestamp 28801
transform 1 0 19964 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2824_
timestamp 28801
transform 1 0 21436 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2825_
timestamp 28801
transform 1 0 25116 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2826_
timestamp 28801
transform 1 0 26588 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2827_
timestamp 28801
transform 1 0 26220 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2828_
timestamp 28801
transform -1 0 29072 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2829_
timestamp 28801
transform 1 0 30452 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2830_
timestamp 28801
transform 1 0 32108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2831_
timestamp 28801
transform -1 0 33580 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2832_
timestamp 28801
transform -1 0 35512 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2833_
timestamp 28801
transform -1 0 36616 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2834_
timestamp 28801
transform 1 0 34684 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2835_
timestamp 28801
transform 1 0 32200 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2836_
timestamp 28801
transform 1 0 14076 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _2837_
timestamp 28801
transform -1 0 3588 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2838_
timestamp 28801
transform 1 0 1564 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2839_
timestamp 28801
transform 1 0 4968 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2840_
timestamp 28801
transform 1 0 15088 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 28801
transform 1 0 40296 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 28801
transform 1 0 37720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 28801
transform 1 0 20608 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 28801
transform -1 0 10948 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 28801
transform 1 0 12052 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 28801
transform 1 0 31096 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 28801
transform 1 0 32108 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_0_clk
timestamp 28801
transform -1 0 3220 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_1_clk
timestamp 28801
transform 1 0 6808 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_2_clk
timestamp 28801
transform 1 0 2484 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_3_clk
timestamp 28801
transform -1 0 9200 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_4_clk
timestamp 28801
transform 1 0 14076 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_5_clk
timestamp 28801
transform -1 0 17664 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_6_clk
timestamp 28801
transform 1 0 11500 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_7_clk
timestamp 28801
transform 1 0 5244 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_8_clk
timestamp 28801
transform -1 0 5428 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_9_clk
timestamp 28801
transform 1 0 7636 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_10_clk
timestamp 28801
transform -1 0 8188 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_11_clk
timestamp 28801
transform 1 0 14076 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_12_clk
timestamp 28801
transform 1 0 19504 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_13_clk
timestamp 28801
transform 1 0 17756 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_14_clk
timestamp 28801
transform 1 0 16836 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_15_clk
timestamp 28801
transform -1 0 24196 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_16_clk
timestamp 28801
transform 1 0 26680 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_17_clk
timestamp 28801
transform 1 0 23368 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_18_clk
timestamp 28801
transform -1 0 31004 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_19_clk
timestamp 28801
transform 1 0 32844 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_20_clk
timestamp 28801
transform 1 0 38272 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_21_clk
timestamp 28801
transform 1 0 39100 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_22_clk
timestamp 28801
transform 1 0 39100 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_23_clk
timestamp 28801
transform -1 0 38272 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_24_clk
timestamp 28801
transform 1 0 31096 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_25_clk
timestamp 28801
transform -1 0 29072 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_26_clk
timestamp 28801
transform 1 0 32108 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_27_clk
timestamp 28801
transform 1 0 38180 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_28_clk
timestamp 28801
transform 1 0 38088 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_29_clk
timestamp 28801
transform 1 0 37352 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_30_clk
timestamp 28801
transform -1 0 38272 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_31_clk
timestamp 28801
transform 1 0 32108 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_32_clk
timestamp 28801
transform 1 0 25668 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_33_clk
timestamp 28801
transform 1 0 25208 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_34_clk
timestamp 28801
transform 1 0 27416 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_35_clk
timestamp 28801
transform -1 0 23368 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_36_clk
timestamp 28801
transform 1 0 16652 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_37_clk
timestamp 28801
transform 1 0 18124 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_38_clk
timestamp 28801
transform 1 0 10396 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_39_clk
timestamp 28801
transform -1 0 5428 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinvlp_4  clkload0
timestamp 28801
transform 1 0 9108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload1
timestamp 28801
transform 1 0 12052 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp 28801
transform 1 0 31004 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_8  clkload3
timestamp 28801
transform 1 0 3312 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload4
timestamp 28801
transform 1 0 6808 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload5
timestamp 28801
transform 1 0 1564 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload6
timestamp 28801
transform 1 0 8188 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload7
timestamp 28801
transform 1 0 13248 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload8
timestamp 28801
transform 1 0 18124 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  clkload9
timestamp 28801
transform 1 0 11500 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload10
timestamp 28801
transform 1 0 4416 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  clkload11
timestamp 28801
transform 1 0 17572 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload12
timestamp 28801
transform 1 0 5428 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload13
timestamp 28801
transform 1 0 4416 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload14
timestamp 28801
transform 1 0 7636 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  clkload15
timestamp 28801
transform 1 0 7176 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload16
timestamp 28801
transform 1 0 13156 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload17
timestamp 28801
transform 1 0 19504 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  clkload18
timestamp 28801
transform 1 0 18676 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__inv_6  clkload19
timestamp 28801
transform 1 0 17296 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload20
timestamp 28801
transform 1 0 27784 0 -1 22848
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload21
timestamp 28801
transform 1 0 32108 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__bufinv_16  clkload22
timestamp 28801
transform 1 0 37720 0 -1 21760
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_8  clkload23
timestamp 28801
transform 1 0 38088 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload24
timestamp 28801
transform 1 0 37352 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  clkload25
timestamp 28801
transform 1 0 37444 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  clkload26
timestamp 28801
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_6  clkload27
timestamp 28801
transform 1 0 26220 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload28
timestamp 28801
transform 1 0 26220 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  clkload29
timestamp 28801
transform 1 0 27416 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload30
timestamp 28801
transform 1 0 23092 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload31
timestamp 28801
transform 1 0 23092 0 1 39168
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload32
timestamp 28801
transform 1 0 28796 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload33
timestamp 28801
transform 1 0 32844 0 -1 38080
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload34
timestamp 28801
transform 1 0 38272 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  clkload35
timestamp 28801
transform 1 0 37352 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_4  clkload36
timestamp 28801
transform 1 0 39192 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  clkload37
timestamp 28801
transform 1 0 36892 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  clkload38
timestamp 28801
transform 1 0 30820 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 28801
transform -1 0 31096 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 28801
transform -1 0 31372 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 28801
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout34
timestamp 28801
transform 1 0 17204 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 28801
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 28801
transform -1 0 4140 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 28801
transform -1 0 3588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 28801
transform 1 0 7820 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 28801
transform -1 0 38364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 28801
transform 1 0 23000 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 28801
transform 1 0 17112 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 28801
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 28801
transform -1 0 18308 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 28801
transform -1 0 16560 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 28801
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 28801
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 28801
transform -1 0 21712 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 28801
transform 1 0 32936 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 28801
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 28801
transform 1 0 25760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 28801
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 28801
transform -1 0 22632 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp 28801
transform 1 0 38916 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 28801
transform -1 0 17296 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp 28801
transform 1 0 27876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 28801
transform -1 0 26588 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout57
timestamp 28801
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 28801
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 28801
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 28801
transform -1 0 22724 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout61
timestamp 28801
transform 1 0 32108 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 28801
transform -1 0 17940 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 28801
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout64
timestamp 28801
transform -1 0 42044 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp 28801
transform 1 0 17480 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 28801
transform -1 0 22356 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp 28801
transform 1 0 29900 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout68
timestamp 28801
transform -1 0 19136 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 28801
transform 1 0 32844 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout70
timestamp 28801
transform 1 0 28796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout71
timestamp 28801
transform -1 0 19596 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout72
timestamp 28801
transform -1 0 20700 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 28801
transform -1 0 22540 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp 28801
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout76
timestamp 28801
transform -1 0 18400 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp 28801
transform 1 0 28428 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout78
timestamp 28801
transform -1 0 26864 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout79
timestamp 28801
transform -1 0 27416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout80
timestamp 28801
transform 1 0 40572 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout81
timestamp 28801
transform 1 0 39192 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 28801
transform 1 0 4968 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout83
timestamp 28801
transform -1 0 6716 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp 28801
transform -1 0 20884 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout86
timestamp 28801
transform -1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout87
timestamp 28801
transform 1 0 28704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp 28801
transform -1 0 26772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout89
timestamp 28801
transform -1 0 37720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout90
timestamp 28801
transform 1 0 38088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp 28801
transform 1 0 37996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 28801
transform -1 0 5244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 28801
transform -1 0 15456 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout94
timestamp 28801
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout95
timestamp 28801
transform -1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout96
timestamp 28801
transform -1 0 31832 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 28801
transform 1 0 33948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout98
timestamp 28801
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout99
timestamp 28801
transform -1 0 20056 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout100
timestamp 28801
transform -1 0 31924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout101
timestamp 28801
transform 1 0 35696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout102
timestamp 28801
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout103
timestamp 28801
transform -1 0 30268 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout104
timestamp 28801
transform -1 0 28704 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout105
timestamp 28801
transform 1 0 31372 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp 28801
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp 28801
transform -1 0 31924 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 28801
transform 1 0 39376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout109
timestamp 28801
transform 1 0 17388 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout110
timestamp 28801
transform -1 0 13984 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout111
timestamp 28801
transform -1 0 25576 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout112
timestamp 28801
transform -1 0 29256 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 28801
transform 1 0 38640 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout114
timestamp 28801
transform -1 0 18952 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout115
timestamp 28801
transform 1 0 33856 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout116
timestamp 28801
transform 1 0 6532 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout117
timestamp 28801
transform -1 0 6256 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout118
timestamp 28801
transform 1 0 13616 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout119
timestamp 28801
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout120
timestamp 28801
transform -1 0 7636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout121
timestamp 28801
transform 1 0 10396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout122
timestamp 28801
transform -1 0 11316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout123
timestamp 28801
transform -1 0 8096 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout124
timestamp 28801
transform 1 0 6992 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout125
timestamp 28801
transform 1 0 6440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout126
timestamp 28801
transform 1 0 20700 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout127
timestamp 28801
transform -1 0 21436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout128
timestamp 28801
transform -1 0 19872 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout129
timestamp 28801
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout130
timestamp 28801
transform -1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout131
timestamp 28801
transform -1 0 6900 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout132
timestamp 28801
transform 1 0 12696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout133
timestamp 28801
transform -1 0 13064 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout134
timestamp 28801
transform -1 0 18032 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout135
timestamp 28801
transform -1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout136
timestamp 28801
transform -1 0 17204 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout137
timestamp 28801
transform -1 0 22172 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout138
timestamp 28801
transform -1 0 23000 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout139
timestamp 28801
transform -1 0 25668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout140
timestamp 28801
transform -1 0 27876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout141
timestamp 28801
transform -1 0 30820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout142
timestamp 28801
transform -1 0 32016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout143
timestamp 28801
transform -1 0 28244 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout144
timestamp 28801
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout145
timestamp 28801
transform -1 0 31188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout146
timestamp 28801
transform -1 0 38456 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout147
timestamp 28801
transform -1 0 35696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout148
timestamp 28801
transform -1 0 39008 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout149
timestamp 28801
transform -1 0 42044 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout150
timestamp 28801
transform 1 0 41400 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout151
timestamp 28801
transform 1 0 38732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout152
timestamp 28801
transform -1 0 31648 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout153
timestamp 28801
transform -1 0 28244 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout154
timestamp 28801
transform -1 0 31924 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout155
timestamp 28801
transform -1 0 32476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout156
timestamp 28801
transform -1 0 42228 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout157
timestamp 28801
transform 1 0 41676 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout158
timestamp 28801
transform -1 0 37168 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout159
timestamp 28801
transform 1 0 41768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout160
timestamp 28801
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636997256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636997256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 28801
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636997256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636997256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 28801
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636997256
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636997256
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 28801
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636997256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636997256
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 28801
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 28801
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 1636997256
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 28801
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 28801
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636997256
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636997256
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 28801
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636997256
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636997256
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 28801
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636997256
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636997256
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 28801
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636997256
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636997256
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 28801
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636997256
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636997256
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 28801
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636997256
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636997256
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 28801
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636997256
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636997256
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 28801
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636997256
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636997256
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 28801
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636997256
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636997256
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 28801
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1636997256
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636997256
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 28801
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1636997256
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1636997256
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_445
timestamp 28801
transform 1 0 42044 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636997256
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636997256
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636997256
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636997256
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 28801
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 28801
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636997256
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636997256
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636997256
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636997256
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 28801
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 28801
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636997256
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636997256
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636997256
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636997256
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 28801
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 28801
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636997256
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636997256
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636997256
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636997256
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 28801
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 28801
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636997256
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636997256
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636997256
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636997256
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 28801
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 28801
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636997256
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636997256
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636997256
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636997256
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 28801
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 28801
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636997256
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636997256
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636997256
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636997256
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 28801
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 28801
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636997256
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636997256
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636997256
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636997256
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 28801
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636997256
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636997256
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 28801
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636997256
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636997256
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636997256
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636997256
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 28801
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 28801
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636997256
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636997256
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636997256
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636997256
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 28801
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 28801
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636997256
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636997256
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636997256
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636997256
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 28801
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 28801
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636997256
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636997256
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636997256
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636997256
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 28801
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 28801
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636997256
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636997256
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636997256
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636997256
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 28801
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 28801
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636997256
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636997256
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636997256
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636997256
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 28801
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 28801
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636997256
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636997256
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636997256
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636997256
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 28801
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 28801
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636997256
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636997256
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_445
timestamp 28801
transform 1 0 42044 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636997256
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636997256
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636997256
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636997256
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 28801
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 28801
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636997256
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636997256
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636997256
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636997256
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 28801
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 28801
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636997256
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636997256
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636997256
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636997256
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 28801
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 28801
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636997256
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636997256
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636997256
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636997256
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 28801
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 28801
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636997256
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636997256
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636997256
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636997256
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 28801
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 28801
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636997256
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636997256
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636997256
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636997256
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 28801
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 28801
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636997256
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636997256
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636997256
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636997256
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 28801
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 28801
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636997256
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636997256
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636997256
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636997256
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 28801
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636997256
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636997256
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 28801
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636997256
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_56
timestamp 28801
transform 1 0 6256 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 28801
transform 1 0 6992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_71
timestamp 28801
transform 1 0 7636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 28801
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636997256
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636997256
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636997256
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636997256
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 28801
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 28801
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636997256
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636997256
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636997256
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636997256
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 28801
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 28801
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636997256
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636997256
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636997256
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636997256
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 28801
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 28801
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636997256
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636997256
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636997256
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636997256
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 28801
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 28801
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636997256
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_321
timestamp 28801
transform 1 0 30636 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_347
timestamp 1636997256
transform 1 0 33028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_359
timestamp 28801
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 28801
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636997256
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636997256
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636997256
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636997256
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 28801
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 28801
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636997256
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636997256
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_445
timestamp 28801
transform 1 0 42044 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636997256
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_15
timestamp 28801
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_21
timestamp 28801
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_25
timestamp 28801
transform 1 0 3404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 28801
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 28801
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636997256
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 28801
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 28801
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636997256
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636997256
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636997256
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636997256
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 28801
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 28801
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636997256
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636997256
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636997256
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636997256
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 28801
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 28801
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_225
timestamp 28801
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_233
timestamp 1636997256
transform 1 0 22540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_245
timestamp 1636997256
transform 1 0 23644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_257
timestamp 1636997256
transform 1 0 24748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 28801
transform 1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 28801
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636997256
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_293
timestamp 28801
transform 1 0 28060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_314
timestamp 28801
transform 1 0 29992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_327
timestamp 28801
transform 1 0 31188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 28801
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_345
timestamp 1636997256
transform 1 0 32844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_357
timestamp 28801
transform 1 0 33948 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_372
timestamp 1636997256
transform 1 0 35328 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_384
timestamp 28801
transform 1 0 36432 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636997256
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636997256
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636997256
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636997256
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 28801
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 28801
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 28801
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_51
timestamp 28801
transform 1 0 5796 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 28801
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_88
timestamp 28801
transform 1 0 9200 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636997256
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636997256
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 28801
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 28801
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636997256
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636997256
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636997256
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636997256
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 28801
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 28801
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636997256
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636997256
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_221
timestamp 28801
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp 28801
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 28801
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636997256
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636997256
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636997256
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636997256
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 28801
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 28801
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 28801
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 28801
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_373
timestamp 28801
transform 1 0 35420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_377
timestamp 28801
transform 1 0 35788 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_398
timestamp 1636997256
transform 1 0 37720 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_410
timestamp 28801
transform 1 0 38824 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 28801
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636997256
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_433
timestamp 28801
transform 1 0 40940 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_441
timestamp 28801
transform 1 0 41676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_23
timestamp 28801
transform 1 0 3220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_29
timestamp 28801
transform 1 0 3772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 28801
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_97
timestamp 28801
transform 1 0 10028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 28801
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636997256
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636997256
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636997256
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636997256
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 28801
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 28801
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636997256
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_181
timestamp 28801
transform 1 0 17756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_187
timestamp 28801
transform 1 0 18308 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 28801
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_212
timestamp 28801
transform 1 0 20608 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 28801
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 28801
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 28801
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 28801
transform 1 0 22724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_239
timestamp 28801
transform 1 0 23092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_260
timestamp 28801
transform 1 0 25024 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_267
timestamp 1636997256
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 28801
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_309
timestamp 28801
transform 1 0 29532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_327
timestamp 28801
transform 1 0 31188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_345
timestamp 28801
transform 1 0 32844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_369
timestamp 28801
transform 1 0 35052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 28801
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_397
timestamp 1636997256
transform 1 0 37628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_409
timestamp 1636997256
transform 1 0 38732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_421
timestamp 1636997256
transform 1 0 39836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_433
timestamp 1636997256
transform 1 0 40940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_445
timestamp 28801
transform 1 0 42044 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636997256
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_15
timestamp 28801
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 28801
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 28801
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_78
timestamp 28801
transform 1 0 8280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_91
timestamp 28801
transform 1 0 9476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 28801
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1636997256
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 28801
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 28801
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636997256
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636997256
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636997256
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636997256
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 28801
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 28801
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 28801
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_241
timestamp 28801
transform 1 0 23276 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_293
timestamp 28801
transform 1 0 28060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 28801
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 28801
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_323
timestamp 28801
transform 1 0 30820 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_332
timestamp 1636997256
transform 1 0 31648 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 28801
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_375
timestamp 28801
transform 1 0 35604 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_412
timestamp 28801
transform 1 0 39008 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636997256
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636997256
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_445
timestamp 28801
transform 1 0 42044 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 28801
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_13
timestamp 1636997256
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_25
timestamp 1636997256
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1636997256
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 28801
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 28801
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636997256
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636997256
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636997256
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636997256
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 28801
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 28801
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 28801
transform 1 0 11960 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_133
timestamp 1636997256
transform 1 0 13340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_145
timestamp 1636997256
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp 28801
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 28801
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636997256
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636997256
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 28801
transform 1 0 18860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_203
timestamp 28801
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_214
timestamp 28801
transform 1 0 20792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 28801
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 28801
transform 1 0 23644 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 28801
transform 1 0 24012 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 28801
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_342
timestamp 1636997256
transform 1 0 32568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_354
timestamp 28801
transform 1 0 33672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_378
timestamp 28801
transform 1 0 35880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 28801
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_413
timestamp 1636997256
transform 1 0 39100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_425
timestamp 1636997256
transform 1 0 40204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_437
timestamp 28801
transform 1 0 41308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_445
timestamp 28801
transform 1 0 42044 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_34
timestamp 1636997256
transform 1 0 4232 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_46
timestamp 1636997256
transform 1 0 5336 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_58
timestamp 1636997256
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_70
timestamp 28801
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_78
timestamp 28801
transform 1 0 8280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_92
timestamp 28801
transform 1 0 9568 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_117
timestamp 28801
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 28801
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636997256
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636997256
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636997256
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636997256
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_216
timestamp 1636997256
transform 1 0 20976 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_228
timestamp 1636997256
transform 1 0 22080 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_240
timestamp 1636997256
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_260
timestamp 28801
transform 1 0 25024 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_285
timestamp 1636997256
transform 1 0 27324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_297
timestamp 28801
transform 1 0 28428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_329
timestamp 28801
transform 1 0 31372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_345
timestamp 28801
transform 1 0 32844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_349
timestamp 28801
transform 1 0 33212 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_358
timestamp 28801
transform 1 0 34040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_365
timestamp 28801
transform 1 0 34684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_373
timestamp 28801
transform 1 0 35420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_411
timestamp 28801
transform 1 0 38916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 28801
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1636997256
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1636997256
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_445
timestamp 28801
transform 1 0 42044 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 28801
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_40
timestamp 28801
transform 1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_48
timestamp 28801
transform 1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_64
timestamp 28801
transform 1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_68
timestamp 28801
transform 1 0 7360 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_155
timestamp 1636997256
transform 1 0 15364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 28801
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636997256
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_181
timestamp 28801
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 28801
transform 1 0 19136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 28801
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 28801
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_242
timestamp 1636997256
transform 1 0 23368 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_254
timestamp 28801
transform 1 0 24472 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_260
timestamp 28801
transform 1 0 25024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 28801
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_286
timestamp 28801
transform 1 0 27416 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_294
timestamp 28801
transform 1 0 28152 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_323
timestamp 1636997256
transform 1 0 30820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 28801
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_377
timestamp 28801
transform 1 0 35788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_382
timestamp 28801
transform 1 0 36248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_386
timestamp 28801
transform 1 0 36616 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_393
timestamp 28801
transform 1 0 37260 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_422
timestamp 1636997256
transform 1 0 39928 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_434
timestamp 1636997256
transform 1 0 41032 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_446
timestamp 28801
transform 1 0 42136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_43
timestamp 28801
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_59
timestamp 28801
transform 1 0 6532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_68
timestamp 28801
transform 1 0 7360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 28801
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_89
timestamp 28801
transform 1 0 9292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_122
timestamp 28801
transform 1 0 12328 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 28801
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 28801
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636997256
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636997256
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_165
timestamp 28801
transform 1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_173
timestamp 28801
transform 1 0 17020 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_212
timestamp 28801
transform 1 0 20608 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_220
timestamp 28801
transform 1 0 21344 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_236
timestamp 1636997256
transform 1 0 22816 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 28801
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 28801
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_283
timestamp 1636997256
transform 1 0 27140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_295
timestamp 1636997256
transform 1 0 28244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 28801
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_317
timestamp 1636997256
transform 1 0 30268 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_329
timestamp 28801
transform 1 0 31372 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_352
timestamp 1636997256
transform 1 0 33488 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1636997256
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_377
timestamp 28801
transform 1 0 35788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_387
timestamp 28801
transform 1 0 36708 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_409
timestamp 28801
transform 1 0 38732 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_417
timestamp 28801
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1636997256
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1636997256
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_445
timestamp 28801
transform 1 0 42044 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636997256
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_18
timestamp 28801
transform 1 0 2760 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1636997256
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_35
timestamp 28801
transform 1 0 4324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_43
timestamp 28801
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 28801
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp 28801
transform 1 0 7820 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_82
timestamp 1636997256
transform 1 0 8648 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_94
timestamp 28801
transform 1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_126
timestamp 1636997256
transform 1 0 12696 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_138
timestamp 1636997256
transform 1 0 13800 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_150
timestamp 1636997256
transform 1 0 14904 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 28801
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636997256
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 28801
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_192
timestamp 28801
transform 1 0 18768 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_198
timestamp 28801
transform 1 0 19320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_212
timestamp 28801
transform 1 0 20608 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_218
timestamp 28801
transform 1 0 21160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 28801
transform 1 0 23644 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 28801
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_288
timestamp 28801
transform 1 0 27600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_312
timestamp 28801
transform 1 0 29808 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_320
timestamp 28801
transform 1 0 30544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_328
timestamp 28801
transform 1 0 31280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_348
timestamp 28801
transform 1 0 33120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_352
timestamp 28801
transform 1 0 33488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_378
timestamp 28801
transform 1 0 35880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_387
timestamp 28801
transform 1 0 36708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 28801
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_393
timestamp 28801
transform 1 0 37260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_406
timestamp 28801
transform 1 0 38456 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_428
timestamp 1636997256
transform 1 0 40480 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_440
timestamp 28801
transform 1 0 41584 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_446
timestamp 28801
transform 1 0 42136 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636997256
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_15
timestamp 28801
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_21
timestamp 28801
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 28801
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636997256
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 28801
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 28801
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_68
timestamp 1636997256
transform 1 0 7360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 28801
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636997256
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636997256
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 28801
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 28801
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_122
timestamp 28801
transform 1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_161
timestamp 1636997256
transform 1 0 15916 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_173
timestamp 1636997256
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_185
timestamp 28801
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 28801
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1636997256
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_209
timestamp 28801
transform 1 0 20332 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_230
timestamp 28801
transform 1 0 22264 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 28801
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_268
timestamp 28801
transform 1 0 25760 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_272
timestamp 28801
transform 1 0 26128 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 28801
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_328
timestamp 28801
transform 1 0 31280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_355
timestamp 28801
transform 1 0 33764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_389
timestamp 28801
transform 1 0 36892 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_415
timestamp 28801
transform 1 0 39284 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 28801
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_435
timestamp 1636997256
transform 1 0 41124 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_7
timestamp 28801
transform 1 0 1748 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_13
timestamp 28801
transform 1 0 2300 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_17
timestamp 28801
transform 1 0 2668 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_22
timestamp 28801
transform 1 0 3128 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_42
timestamp 28801
transform 1 0 4968 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 28801
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_60
timestamp 28801
transform 1 0 6624 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_94
timestamp 1636997256
transform 1 0 9752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 28801
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 28801
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636997256
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 28801
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 28801
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 28801
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 28801
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_229
timestamp 28801
transform 1 0 22172 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_253
timestamp 1636997256
transform 1 0 24380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_290
timestamp 28801
transform 1 0 27784 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_296
timestamp 28801
transform 1 0 28336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_306
timestamp 28801
transform 1 0 29256 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_315
timestamp 1636997256
transform 1 0 30084 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_327
timestamp 28801
transform 1 0 31188 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 28801
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_354
timestamp 28801
transform 1 0 33672 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_364
timestamp 28801
transform 1 0 34592 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_383
timestamp 28801
transform 1 0 36340 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 28801
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_393
timestamp 28801
transform 1 0 37260 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_433
timestamp 1636997256
transform 1 0 40940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_445
timestamp 28801
transform 1 0 42044 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 28801
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_49
timestamp 28801
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_57
timestamp 28801
transform 1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_62
timestamp 1636997256
transform 1 0 6808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_74
timestamp 28801
transform 1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_105
timestamp 28801
transform 1 0 10764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_113
timestamp 28801
transform 1 0 11500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_129
timestamp 28801
transform 1 0 12972 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 28801
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_151
timestamp 28801
transform 1 0 14996 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_180
timestamp 28801
transform 1 0 17664 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_186
timestamp 28801
transform 1 0 18216 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_217
timestamp 28801
transform 1 0 21068 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_232
timestamp 28801
transform 1 0 22448 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_242
timestamp 28801
transform 1 0 23368 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 28801
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_287
timestamp 28801
transform 1 0 27508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_297
timestamp 28801
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 28801
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_343
timestamp 1636997256
transform 1 0 32660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_355
timestamp 28801
transform 1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 28801
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_365
timestamp 28801
transform 1 0 34684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_369
timestamp 28801
transform 1 0 35052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_376
timestamp 28801
transform 1 0 35696 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_400
timestamp 28801
transform 1 0 37904 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_405
timestamp 1636997256
transform 1 0 38364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_417
timestamp 28801
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1636997256
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1636997256
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_445
timestamp 28801
transform 1 0 42044 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 28801
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_42
timestamp 28801
transform 1 0 4968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 28801
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 28801
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_75
timestamp 28801
transform 1 0 8004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_102
timestamp 28801
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 28801
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 28801
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 28801
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp 28801
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 28801
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636997256
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 28801
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_189
timestamp 28801
transform 1 0 18492 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_195
timestamp 28801
transform 1 0 19044 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 28801
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 28801
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 28801
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_271
timestamp 28801
transform 1 0 26036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_311
timestamp 28801
transform 1 0 29716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_323
timestamp 28801
transform 1 0 30820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_337
timestamp 28801
transform 1 0 32108 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1636997256
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_405
timestamp 28801
transform 1 0 38364 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1636997256
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 28801
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 28801
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 28801
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 28801
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 28801
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 28801
transform 1 0 5336 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_66
timestamp 28801
transform 1 0 7176 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 28801
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 28801
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 28801
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 28801
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 28801
transform 1 0 12880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 28801
transform 1 0 13248 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_149
timestamp 1636997256
transform 1 0 14812 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_161
timestamp 28801
transform 1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_183
timestamp 1636997256
transform 1 0 17940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 28801
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 28801
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_253
timestamp 28801
transform 1 0 24380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_263
timestamp 28801
transform 1 0 25300 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 28801
transform 1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_284
timestamp 28801
transform 1 0 27232 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 28801
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_322
timestamp 28801
transform 1 0 30728 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 28801
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_376
timestamp 28801
transform 1 0 35696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_393
timestamp 28801
transform 1 0 37260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_440
timestamp 28801
transform 1 0 41584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_446
timestamp 28801
transform 1 0 42136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 28801
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 28801
transform 1 0 4324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_39
timestamp 28801
transform 1 0 4692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 28801
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 28801
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 28801
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_64
timestamp 1636997256
transform 1 0 6992 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_76
timestamp 28801
transform 1 0 8096 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 28801
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 28801
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 28801
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_155
timestamp 1636997256
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 28801
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636997256
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 28801
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 28801
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_197
timestamp 28801
transform 1 0 19228 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_206
timestamp 1636997256
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 28801
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 28801
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_231
timestamp 28801
transform 1 0 22356 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_241
timestamp 1636997256
transform 1 0 23276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_253
timestamp 28801
transform 1 0 24380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_261
timestamp 28801
transform 1 0 25116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 28801
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 28801
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 28801
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 28801
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_305
timestamp 28801
transform 1 0 29164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_330
timestamp 28801
transform 1 0 31464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_371
timestamp 28801
transform 1 0 35236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_380
timestamp 28801
transform 1 0 36064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 28801
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_393
timestamp 28801
transform 1 0 37260 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_437
timestamp 28801
transform 1 0 41308 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_445
timestamp 28801
transform 1 0 42044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 28801
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 28801
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_37
timestamp 28801
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_46
timestamp 28801
transform 1 0 5336 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_50
timestamp 28801
transform 1 0 5704 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 28801
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 28801
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 28801
transform 1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 28801
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 28801
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_153
timestamp 28801
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_183
timestamp 1636997256
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 28801
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_204
timestamp 28801
transform 1 0 19872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 28801
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_253
timestamp 28801
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_284
timestamp 28801
transform 1 0 27232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 28801
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 28801
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1636997256
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_321
timestamp 28801
transform 1 0 30636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_325
timestamp 28801
transform 1 0 31004 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 28801
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_372
timestamp 28801
transform 1 0 35328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_403
timestamp 28801
transform 1 0 38180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 28801
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_421
timestamp 28801
transform 1 0 39836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_7
timestamp 28801
transform 1 0 1748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_44
timestamp 28801
transform 1 0 5152 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 28801
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 28801
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_63
timestamp 1636997256
transform 1 0 6900 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_75
timestamp 1636997256
transform 1 0 8004 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 28801
transform 1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_91
timestamp 28801
transform 1 0 9476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 28801
transform 1 0 12420 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_129
timestamp 1636997256
transform 1 0 12972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_141
timestamp 1636997256
transform 1 0 14076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_153
timestamp 1636997256
transform 1 0 15180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 28801
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_209
timestamp 28801
transform 1 0 20332 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_215
timestamp 28801
transform 1 0 20884 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 28801
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_236
timestamp 28801
transform 1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 28801
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_305
timestamp 28801
transform 1 0 29164 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_313
timestamp 28801
transform 1 0 29900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_337
timestamp 28801
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 28801
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 28801
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_401
timestamp 28801
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_406
timestamp 28801
transform 1 0 38456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_412
timestamp 28801
transform 1 0 39008 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_420
timestamp 28801
transform 1 0 39744 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_426
timestamp 28801
transform 1 0 40296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_438
timestamp 28801
transform 1 0 41400 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 28801
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_37
timestamp 28801
transform 1 0 4508 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 28801
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1636997256
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 28801
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_101
timestamp 28801
transform 1 0 10396 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_106
timestamp 1636997256
transform 1 0 10856 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_118
timestamp 1636997256
transform 1 0 11960 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 28801
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 28801
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636997256
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 28801
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 28801
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 28801
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_224
timestamp 28801
transform 1 0 21712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 28801
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 28801
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_282
timestamp 28801
transform 1 0 27048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 28801
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 28801
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_355
timestamp 28801
transform 1 0 33764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_365
timestamp 28801
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_369
timestamp 28801
transform 1 0 35052 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_378
timestamp 1636997256
transform 1 0 35880 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_390
timestamp 28801
transform 1 0 36984 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_398
timestamp 28801
transform 1 0 37720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_409
timestamp 28801
transform 1 0 38732 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_433
timestamp 28801
transform 1 0 40940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_437
timestamp 28801
transform 1 0 41308 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_444
timestamp 28801
transform 1 0 41952 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636997256
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_15
timestamp 28801
transform 1 0 2484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_42
timestamp 28801
transform 1 0 4968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_50
timestamp 28801
transform 1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 28801
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 28801
transform 1 0 7820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_106
timestamp 28801
transform 1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 28801
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 28801
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_130
timestamp 28801
transform 1 0 13064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_134
timestamp 28801
transform 1 0 13432 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_151
timestamp 28801
transform 1 0 14996 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 28801
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 28801
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 28801
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_235
timestamp 1636997256
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_247
timestamp 28801
transform 1 0 23828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_253
timestamp 28801
transform 1 0 24380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_262
timestamp 28801
transform 1 0 25208 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 28801
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_281
timestamp 28801
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 28801
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 28801
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_348
timestamp 28801
transform 1 0 33120 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_361
timestamp 28801
transform 1 0 34316 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_367
timestamp 28801
transform 1 0 34868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_375
timestamp 28801
transform 1 0 35604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 28801
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 28801
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_423
timestamp 28801
transform 1 0 40020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_444
timestamp 28801
transform 1 0 41952 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_6
timestamp 28801
transform 1 0 1656 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636997256
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 28801
transform 1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 28801
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 28801
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 28801
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636997256
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_153
timestamp 28801
transform 1 0 15180 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_191
timestamp 28801
transform 1 0 18676 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 28801
transform 1 0 20516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_222
timestamp 28801
transform 1 0 21528 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_232
timestamp 28801
transform 1 0 22448 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_236
timestamp 28801
transform 1 0 22816 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_240
timestamp 1636997256
transform 1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_261
timestamp 28801
transform 1 0 25116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_271
timestamp 28801
transform 1 0 26036 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_277
timestamp 28801
transform 1 0 26588 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 28801
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_312
timestamp 1636997256
transform 1 0 29808 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_324
timestamp 28801
transform 1 0 30912 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_342
timestamp 1636997256
transform 1 0 32568 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 28801
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 28801
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_365
timestamp 28801
transform 1 0 34684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_391
timestamp 28801
transform 1 0 37076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_412
timestamp 28801
transform 1 0 39008 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 28801
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_428
timestamp 28801
transform 1 0 40480 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_445
timestamp 28801
transform 1 0 42044 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_6
timestamp 28801
transform 1 0 1656 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 28801
transform 1 0 2392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_37
timestamp 28801
transform 1 0 4508 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_45
timestamp 28801
transform 1 0 5244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_49
timestamp 28801
transform 1 0 5612 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 28801
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636997256
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636997256
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_86
timestamp 1636997256
transform 1 0 9016 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_98
timestamp 1636997256
transform 1 0 10120 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 28801
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 28801
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_150
timestamp 28801
transform 1 0 14904 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_210
timestamp 28801
transform 1 0 20424 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_228
timestamp 1636997256
transform 1 0 22080 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_240
timestamp 28801
transform 1 0 23184 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_263
timestamp 1636997256
transform 1 0 25300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 28801
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 28801
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_311
timestamp 28801
transform 1 0 29716 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 28801
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1636997256
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_349
timestamp 28801
transform 1 0 33212 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_375
timestamp 1636997256
transform 1 0 35604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_387
timestamp 28801
transform 1 0 36708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 28801
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_419
timestamp 28801
transform 1 0 39652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_432
timestamp 28801
transform 1 0 40848 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_443
timestamp 28801
transform 1 0 41860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 28801
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_37
timestamp 28801
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_58
timestamp 1636997256
transform 1 0 6440 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_70
timestamp 28801
transform 1 0 7544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_74
timestamp 28801
transform 1 0 7912 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 28801
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_92
timestamp 28801
transform 1 0 9568 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 28801
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_108
timestamp 28801
transform 1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 28801
transform 1 0 11960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_122
timestamp 28801
transform 1 0 12328 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636997256
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 28801
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp 28801
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_186
timestamp 28801
transform 1 0 18216 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 28801
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_204
timestamp 28801
transform 1 0 19872 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 28801
transform 1 0 20700 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_236
timestamp 28801
transform 1 0 22816 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_244
timestamp 28801
transform 1 0 23552 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_274
timestamp 28801
transform 1 0 26312 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_282
timestamp 28801
transform 1 0 27048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_292
timestamp 28801
transform 1 0 27968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_351
timestamp 28801
transform 1 0 33396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 28801
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_365
timestamp 28801
transform 1 0 34684 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_386
timestamp 1636997256
transform 1 0 36616 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_398
timestamp 28801
transform 1 0 37720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 28801
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 28801
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_445
timestamp 28801
transform 1 0 42044 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_6
timestamp 28801
transform 1 0 1656 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_14
timestamp 28801
transform 1 0 2392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_67
timestamp 28801
transform 1 0 7268 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 28801
transform 1 0 7636 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_98
timestamp 28801
transform 1 0 10120 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 28801
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 28801
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_119
timestamp 28801
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_145
timestamp 1636997256
transform 1 0 14444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp 28801
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 28801
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 28801
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_177
timestamp 28801
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_186
timestamp 1636997256
transform 1 0 18216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_198
timestamp 28801
transform 1 0 19320 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_228
timestamp 28801
transform 1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 28801
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 28801
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 28801
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_285
timestamp 28801
transform 1 0 27324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_314
timestamp 28801
transform 1 0 29992 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 28801
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_356
timestamp 28801
transform 1 0 33856 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 28801
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_414
timestamp 28801
transform 1 0 39192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_425
timestamp 28801
transform 1 0 40204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_446
timestamp 28801
transform 1 0 42136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 28801
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 28801
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_58
timestamp 28801
transform 1 0 6440 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_64
timestamp 28801
transform 1 0 6992 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 28801
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 28801
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 28801
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_108
timestamp 1636997256
transform 1 0 11040 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_128
timestamp 28801
transform 1 0 12880 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 28801
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_206
timestamp 28801
transform 1 0 20056 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_261
timestamp 28801
transform 1 0 25116 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_302
timestamp 28801
transform 1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_309
timestamp 28801
transform 1 0 29532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 28801
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 28801
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_365
timestamp 28801
transform 1 0 34684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_369
timestamp 28801
transform 1 0 35052 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_375
timestamp 28801
transform 1 0 35604 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_393
timestamp 28801
transform 1 0 37260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_417
timestamp 28801
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_429
timestamp 28801
transform 1 0 40572 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_6
timestamp 1636997256
transform 1 0 1656 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_18
timestamp 1636997256
transform 1 0 2760 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_30
timestamp 1636997256
transform 1 0 3864 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_42
timestamp 1636997256
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 28801
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636997256
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 28801
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 28801
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 28801
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 28801
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 28801
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 28801
transform 1 0 12696 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_146
timestamp 1636997256
transform 1 0 14536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 28801
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 28801
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_178
timestamp 28801
transform 1 0 17480 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 28801
transform 1 0 18032 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1636997256
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 28801
transform 1 0 21068 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 28801
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_233
timestamp 1636997256
transform 1 0 22540 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_245
timestamp 1636997256
transform 1 0 23644 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_257
timestamp 1636997256
transform 1 0 24748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 28801
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_295
timestamp 28801
transform 1 0 28244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_299
timestamp 28801
transform 1 0 28612 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_320
timestamp 28801
transform 1 0 30544 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 28801
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_348
timestamp 28801
transform 1 0 33120 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_360
timestamp 1636997256
transform 1 0 34224 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_372
timestamp 28801
transform 1 0 35328 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_376
timestamp 28801
transform 1 0 35696 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 28801
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_393
timestamp 28801
transform 1 0 37260 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_416
timestamp 28801
transform 1 0 39376 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_420
timestamp 28801
transform 1 0 39744 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636997256
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636997256
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 28801
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_40
timestamp 1636997256
transform 1 0 4784 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_52
timestamp 28801
transform 1 0 5888 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_67
timestamp 28801
transform 1 0 7268 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_73
timestamp 28801
transform 1 0 7820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 28801
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 28801
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 28801
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 28801
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_103
timestamp 28801
transform 1 0 10580 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_112
timestamp 28801
transform 1 0 11408 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_118
timestamp 28801
transform 1 0 11960 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 28801
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1636997256
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1636997256
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_165
timestamp 28801
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_173
timestamp 28801
transform 1 0 17020 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_183
timestamp 28801
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 28801
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 28801
transform 1 0 19872 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_212
timestamp 28801
transform 1 0 20608 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_222
timestamp 1636997256
transform 1 0 21528 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_234
timestamp 28801
transform 1 0 22632 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 28801
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_262
timestamp 28801
transform 1 0 25208 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_279
timestamp 1636997256
transform 1 0 26772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_291
timestamp 28801
transform 1 0 27876 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 28801
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_309
timestamp 28801
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_317
timestamp 28801
transform 1 0 30268 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_328
timestamp 28801
transform 1 0 31280 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_336
timestamp 28801
transform 1 0 32016 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_341
timestamp 28801
transform 1 0 32476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 28801
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 28801
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_388
timestamp 28801
transform 1 0 36800 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_396
timestamp 28801
transform 1 0 37536 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_405
timestamp 28801
transform 1 0 38364 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 28801
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 28801
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_434
timestamp 28801
transform 1 0 41032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_444
timestamp 28801
transform 1 0 41952 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 28801
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_12
timestamp 28801
transform 1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_26
timestamp 28801
transform 1 0 3496 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_45
timestamp 28801
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 28801
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_76
timestamp 28801
transform 1 0 8096 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 28801
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 28801
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_124
timestamp 28801
transform 1 0 12512 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_139
timestamp 1636997256
transform 1 0 13892 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_151
timestamp 1636997256
transform 1 0 14996 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 28801
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 28801
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_178
timestamp 28801
transform 1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_200
timestamp 28801
transform 1 0 19504 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 28801
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_267
timestamp 28801
transform 1 0 25668 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 28801
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_289
timestamp 28801
transform 1 0 27692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 28801
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_366
timestamp 28801
transform 1 0 34776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 28801
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_393
timestamp 28801
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_397
timestamp 28801
transform 1 0 37628 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_407
timestamp 1636997256
transform 1 0 38548 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_419
timestamp 28801
transform 1 0 39652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_437
timestamp 28801
transform 1 0 41308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 28801
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 28801
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_68
timestamp 28801
transform 1 0 7360 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 28801
transform 1 0 10948 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_134
timestamp 28801
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_152
timestamp 28801
transform 1 0 15088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 28801
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_204
timestamp 28801
transform 1 0 19872 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_210
timestamp 28801
transform 1 0 20424 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_242
timestamp 28801
transform 1 0 23368 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 28801
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636997256
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1636997256
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_297
timestamp 28801
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 28801
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1636997256
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_321
timestamp 28801
transform 1 0 30636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 28801
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_388
timestamp 28801
transform 1 0 36800 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 28801
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_421
timestamp 28801
transform 1 0 39836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_442
timestamp 28801
transform 1 0 41768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_446
timestamp 28801
transform 1 0 42136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 28801
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_28
timestamp 28801
transform 1 0 3680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 28801
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 28801
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_62
timestamp 1636997256
transform 1 0 6808 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_74
timestamp 28801
transform 1 0 7912 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_95
timestamp 1636997256
transform 1 0 9844 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 28801
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 28801
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 28801
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_133
timestamp 1636997256
transform 1 0 13340 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 28801
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_207
timestamp 28801
transform 1 0 20148 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_215
timestamp 28801
transform 1 0 20884 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_234
timestamp 28801
transform 1 0 22632 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_238
timestamp 28801
transform 1 0 23000 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_259
timestamp 28801
transform 1 0 24932 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_265
timestamp 28801
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 28801
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 28801
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 28801
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_285
timestamp 28801
transform 1 0 27324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_295
timestamp 28801
transform 1 0 28244 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_316
timestamp 1636997256
transform 1 0 30176 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 28801
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_337
timestamp 28801
transform 1 0 32108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 28801
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_409
timestamp 28801
transform 1 0 38732 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_444
timestamp 28801
transform 1 0 41952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 28801
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 28801
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_41
timestamp 28801
transform 1 0 4876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_45
timestamp 28801
transform 1 0 5244 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_56
timestamp 28801
transform 1 0 6256 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 28801
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_122
timestamp 28801
transform 1 0 12328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 28801
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_180
timestamp 28801
transform 1 0 17664 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_213
timestamp 28801
transform 1 0 20700 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_231
timestamp 1636997256
transform 1 0 22356 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_243
timestamp 28801
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 28801
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_270
timestamp 28801
transform 1 0 25944 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 28801
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_318
timestamp 28801
transform 1 0 30360 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_335
timestamp 28801
transform 1 0 31924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 28801
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 28801
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 28801
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_369
timestamp 28801
transform 1 0 35052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_386
timestamp 28801
transform 1 0 36616 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_392
timestamp 28801
transform 1 0 37168 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 28801
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_421
timestamp 28801
transform 1 0 39836 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636997256
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_15
timestamp 28801
transform 1 0 2484 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_24
timestamp 1636997256
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_50
timestamp 28801
transform 1 0 5704 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1636997256
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 28801
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 28801
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 28801
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_130
timestamp 1636997256
transform 1 0 13064 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_142
timestamp 28801
transform 1 0 14168 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_156
timestamp 28801
transform 1 0 15456 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 28801
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_179
timestamp 1636997256
transform 1 0 17572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_191
timestamp 28801
transform 1 0 18676 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 28801
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 28801
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_242
timestamp 28801
transform 1 0 23368 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_259
timestamp 28801
transform 1 0 24932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_267
timestamp 28801
transform 1 0 25668 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 28801
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_313
timestamp 28801
transform 1 0 29900 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_323
timestamp 28801
transform 1 0 30820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 28801
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_337
timestamp 28801
transform 1 0 32108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_347
timestamp 28801
transform 1 0 33028 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_370
timestamp 28801
transform 1 0 35144 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_374
timestamp 28801
transform 1 0 35512 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_383
timestamp 28801
transform 1 0 36340 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 28801
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_393
timestamp 28801
transform 1 0 37260 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_397
timestamp 28801
transform 1 0 37628 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_446
timestamp 28801
transform 1 0 42136 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_7
timestamp 1636997256
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_19
timestamp 28801
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 28801
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 28801
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_51
timestamp 28801
transform 1 0 5796 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_59
timestamp 28801
transform 1 0 6532 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 28801
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 28801
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_110
timestamp 1636997256
transform 1 0 11224 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_122
timestamp 28801
transform 1 0 12328 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 28801
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_167
timestamp 28801
transform 1 0 16468 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 28801
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_237
timestamp 28801
transform 1 0 22908 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 28801
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_333
timestamp 28801
transform 1 0 31740 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 28801
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_372
timestamp 28801
transform 1 0 35328 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_380
timestamp 28801
transform 1 0 36064 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_414
timestamp 28801
transform 1 0 39192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_445
timestamp 28801
transform 1 0 42044 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_23
timestamp 28801
transform 1 0 3220 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_46
timestamp 28801
transform 1 0 5336 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 28801
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636997256
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_69
timestamp 28801
transform 1 0 7452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_100
timestamp 28801
transform 1 0 10304 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 28801
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 28801
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_130
timestamp 28801
transform 1 0 13064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_180
timestamp 28801
transform 1 0 17664 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_187
timestamp 28801
transform 1 0 18308 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_249
timestamp 28801
transform 1 0 24012 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_281
timestamp 28801
transform 1 0 26956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 28801
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_337
timestamp 28801
transform 1 0 32108 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_376
timestamp 28801
transform 1 0 35696 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_380
timestamp 28801
transform 1 0 36064 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 28801
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 28801
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_401
timestamp 28801
transform 1 0 37996 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_412
timestamp 28801
transform 1 0 39008 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_416
timestamp 28801
transform 1 0 39376 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 28801
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 28801
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636997256
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 28801
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_50
timestamp 1636997256
transform 1 0 5704 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_62
timestamp 28801
transform 1 0 6808 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_73
timestamp 28801
transform 1 0 7820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_81
timestamp 28801
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636997256
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_97
timestamp 28801
transform 1 0 10028 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_114
timestamp 1636997256
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_126
timestamp 28801
transform 1 0 12696 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 28801
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_141
timestamp 28801
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_186
timestamp 28801
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 28801
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_206
timestamp 28801
transform 1 0 20056 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_232
timestamp 28801
transform 1 0 22448 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_241
timestamp 28801
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 28801
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636997256
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_265
timestamp 28801
transform 1 0 25484 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_273
timestamp 1636997256
transform 1 0 26220 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_285
timestamp 28801
transform 1 0 27324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 28801
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 28801
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_317
timestamp 28801
transform 1 0 30268 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_335
timestamp 28801
transform 1 0 31924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_353
timestamp 28801
transform 1 0 33580 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_359
timestamp 28801
transform 1 0 34132 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_390
timestamp 28801
transform 1 0 36984 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_398
timestamp 28801
transform 1 0 37720 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_409
timestamp 28801
transform 1 0 38732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_421
timestamp 28801
transform 1 0 39836 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 28801
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_15
timestamp 28801
transform 1 0 2484 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_23
timestamp 28801
transform 1 0 3220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_61
timestamp 28801
transform 1 0 6716 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_65
timestamp 28801
transform 1 0 7084 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_74
timestamp 28801
transform 1 0 7912 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_82
timestamp 28801
transform 1 0 8648 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_87
timestamp 28801
transform 1 0 9108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 28801
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_117
timestamp 28801
transform 1 0 11868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_151
timestamp 28801
transform 1 0 14996 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_159
timestamp 28801
transform 1 0 15732 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 28801
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_193
timestamp 28801
transform 1 0 18860 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_201
timestamp 28801
transform 1 0 19596 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 28801
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 28801
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_229
timestamp 28801
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_233
timestamp 28801
transform 1 0 22540 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_243
timestamp 28801
transform 1 0 23460 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_251
timestamp 28801
transform 1 0 24196 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 28801
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_304
timestamp 1636997256
transform 1 0 29072 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_319
timestamp 28801
transform 1 0 30452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_323
timestamp 28801
transform 1 0 30820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 28801
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1636997256
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1636997256
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_361
timestamp 28801
transform 1 0 34316 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_365
timestamp 28801
transform 1 0 34684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_371
timestamp 28801
transform 1 0 35236 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_376
timestamp 1636997256
transform 1 0 35696 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 28801
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_414
timestamp 28801
transform 1 0 39192 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_444
timestamp 28801
transform 1 0 41952 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 28801
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_76
timestamp 28801
transform 1 0 8096 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 28801
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_85
timestamp 28801
transform 1 0 8924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_112
timestamp 28801
transform 1 0 11408 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_156
timestamp 1636997256
transform 1 0 15456 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_176
timestamp 28801
transform 1 0 17296 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 28801
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 28801
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 28801
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 28801
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 28801
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 28801
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_316
timestamp 28801
transform 1 0 30176 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_329
timestamp 28801
transform 1 0 31372 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_337
timestamp 28801
transform 1 0 32108 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_347
timestamp 1636997256
transform 1 0 33028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_359
timestamp 28801
transform 1 0 34132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 28801
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_380
timestamp 28801
transform 1 0 36064 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_413
timestamp 28801
transform 1 0 39100 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 28801
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1636997256
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_19
timestamp 28801
transform 1 0 2852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_44
timestamp 28801
transform 1 0 5152 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 28801
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_90
timestamp 28801
transform 1 0 9384 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_100
timestamp 28801
transform 1 0 10304 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 28801
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp 28801
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_125
timestamp 28801
transform 1 0 12604 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_135
timestamp 28801
transform 1 0 13524 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_151
timestamp 28801
transform 1 0 14996 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_157
timestamp 28801
transform 1 0 15548 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 28801
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 28801
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_169
timestamp 28801
transform 1 0 16652 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_176
timestamp 28801
transform 1 0 17296 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_184
timestamp 28801
transform 1 0 18032 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_192
timestamp 28801
transform 1 0 18768 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_210
timestamp 1636997256
transform 1 0 20424 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 28801
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_238
timestamp 1636997256
transform 1 0 23000 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_250
timestamp 28801
transform 1 0 24104 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_256
timestamp 28801
transform 1 0 24656 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_266
timestamp 28801
transform 1 0 25576 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 28801
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 28801
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_295
timestamp 28801
transform 1 0 28244 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_313
timestamp 28801
transform 1 0 29900 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_341
timestamp 28801
transform 1 0 32476 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_357
timestamp 28801
transform 1 0 33948 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_365
timestamp 28801
transform 1 0 34684 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_381
timestamp 28801
transform 1 0 36156 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_404
timestamp 28801
transform 1 0 38272 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 28801
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 28801
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636997256
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_41
timestamp 28801
transform 1 0 4876 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1636997256
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_58
timestamp 1636997256
transform 1 0 6440 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_70
timestamp 28801
transform 1 0 7544 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_74
timestamp 28801
transform 1 0 7912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 28801
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1636997256
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1636997256
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1636997256
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_121
timestamp 28801
transform 1 0 12236 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_129
timestamp 28801
transform 1 0 12972 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 28801
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 28801
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_141
timestamp 28801
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 28801
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 28801
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636997256
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 28801
transform 1 0 20332 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_217
timestamp 28801
transform 1 0 21068 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_231
timestamp 28801
transform 1 0 22356 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_237
timestamp 28801
transform 1 0 22908 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_246
timestamp 28801
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 28801
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_271
timestamp 28801
transform 1 0 26036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_279
timestamp 28801
transform 1 0 26772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_284
timestamp 28801
transform 1 0 27232 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_292
timestamp 28801
transform 1 0 27968 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp 28801
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 28801
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_327
timestamp 1636997256
transform 1 0 31188 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_339
timestamp 28801
transform 1 0 32292 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 28801
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_380
timestamp 28801
transform 1 0 36064 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_387
timestamp 28801
transform 1 0 36708 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_402
timestamp 1636997256
transform 1 0 38088 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_414
timestamp 28801
transform 1 0 39192 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_421
timestamp 28801
transform 1 0 39836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_425
timestamp 28801
transform 1 0 40204 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_433
timestamp 28801
transform 1 0 40940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_7
timestamp 28801
transform 1 0 1748 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_13
timestamp 28801
transform 1 0 2300 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 28801
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 28801
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_86
timestamp 28801
transform 1 0 9016 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 28801
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_122
timestamp 28801
transform 1 0 12328 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_127
timestamp 1636997256
transform 1 0 12788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_139
timestamp 28801
transform 1 0 13892 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_143
timestamp 28801
transform 1 0 14260 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_159
timestamp 28801
transform 1 0 15732 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 28801
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_173
timestamp 1636997256
transform 1 0 17020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_185
timestamp 1636997256
transform 1 0 18124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_197
timestamp 28801
transform 1 0 19228 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_203
timestamp 28801
transform 1 0 19780 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_210
timestamp 28801
transform 1 0 20424 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_216
timestamp 28801
transform 1 0 20976 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 28801
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_239
timestamp 28801
transform 1 0 23092 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_252
timestamp 28801
transform 1 0 24288 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_258
timestamp 28801
transform 1 0 24840 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_265
timestamp 1636997256
transform 1 0 25484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 28801
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 28801
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_287
timestamp 28801
transform 1 0 27508 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_309
timestamp 1636997256
transform 1 0 29532 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_321
timestamp 1636997256
transform 1 0 30636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 28801
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_346
timestamp 1636997256
transform 1 0 32936 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_358
timestamp 1636997256
transform 1 0 34040 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_370
timestamp 1636997256
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 28801
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 28801
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_418
timestamp 28801
transform 1 0 39560 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_435
timestamp 28801
transform 1 0 41124 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_3
timestamp 28801
transform 1 0 1380 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 28801
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_29
timestamp 28801
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_39
timestamp 28801
transform 1 0 4692 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_76
timestamp 28801
transform 1 0 8096 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp 28801
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_149
timestamp 28801
transform 1 0 14812 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_171
timestamp 28801
transform 1 0 16836 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_190
timestamp 28801
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_233
timestamp 28801
transform 1 0 22540 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 28801
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_253
timestamp 28801
transform 1 0 24380 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_275
timestamp 1636997256
transform 1 0 26404 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_287
timestamp 1636997256
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 28801
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 28801
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_309
timestamp 28801
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_322
timestamp 28801
transform 1 0 30728 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_336
timestamp 1636997256
transform 1 0 32016 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_348
timestamp 28801
transform 1 0 33120 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_352
timestamp 28801
transform 1 0 33488 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 28801
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_374
timestamp 28801
transform 1 0 35512 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 28801
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 28801
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_421
timestamp 28801
transform 1 0 39836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_3
timestamp 28801
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_11
timestamp 28801
transform 1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1636997256
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 28801
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_63
timestamp 1636997256
transform 1 0 6900 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_75
timestamp 28801
transform 1 0 8004 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_83
timestamp 28801
transform 1 0 8740 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 28801
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_122
timestamp 1636997256
transform 1 0 12328 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_134
timestamp 1636997256
transform 1 0 13432 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_146
timestamp 28801
transform 1 0 14536 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_157
timestamp 28801
transform 1 0 15548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_161
timestamp 28801
transform 1 0 15916 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_177
timestamp 28801
transform 1 0 17388 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_190
timestamp 28801
transform 1 0 18584 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 28801
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 28801
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 28801
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_233
timestamp 28801
transform 1 0 22540 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_239
timestamp 28801
transform 1 0 23092 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_251
timestamp 28801
transform 1 0 24196 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_259
timestamp 28801
transform 1 0 24932 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_271
timestamp 28801
transform 1 0 26036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 28801
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 28801
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_289
timestamp 28801
transform 1 0 27692 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_307
timestamp 28801
transform 1 0 29348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 28801
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_347
timestamp 28801
transform 1 0 33028 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_368
timestamp 28801
transform 1 0 34960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 28801
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 28801
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 28801
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_401
timestamp 28801
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_411
timestamp 28801
transform 1 0 38916 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_419
timestamp 28801
transform 1 0 39652 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_434
timestamp 28801
transform 1 0 41032 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_442
timestamp 28801
transform 1 0 41768 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636997256
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636997256
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 28801
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_29
timestamp 28801
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_62
timestamp 28801
transform 1 0 6808 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 28801
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 28801
transform 1 0 8924 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_102
timestamp 28801
transform 1 0 10488 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_130
timestamp 28801
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 28801
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 28801
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 28801
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 28801
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 28801
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_213
timestamp 28801
transform 1 0 20700 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_221
timestamp 28801
transform 1 0 21436 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_277
timestamp 28801
transform 1 0 26588 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 28801
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 28801
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_317
timestamp 28801
transform 1 0 30268 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 28801
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_399
timestamp 1636997256
transform 1 0 37812 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_411
timestamp 28801
transform 1 0 38916 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_421
timestamp 28801
transform 1 0 39836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_444
timestamp 28801
transform 1 0 41952 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_7
timestamp 28801
transform 1 0 1748 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_29
timestamp 1636997256
transform 1 0 3772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 28801
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636997256
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_69
timestamp 28801
transform 1 0 7452 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 28801
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_122
timestamp 28801
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_146
timestamp 28801
transform 1 0 14536 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_156
timestamp 1636997256
transform 1 0 15456 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1636997256
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_181
timestamp 28801
transform 1 0 17756 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_190
timestamp 28801
transform 1 0 18584 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_195
timestamp 28801
transform 1 0 19044 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_203
timestamp 28801
transform 1 0 19780 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_207
timestamp 1636997256
transform 1 0 20148 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 28801
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 28801
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636997256
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_237
timestamp 28801
transform 1 0 22908 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_243
timestamp 28801
transform 1 0 23460 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_247
timestamp 28801
transform 1 0 23828 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_269
timestamp 28801
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_277
timestamp 28801
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 28801
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_305
timestamp 28801
transform 1 0 29164 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_326
timestamp 28801
transform 1 0 31096 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 28801
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_344
timestamp 28801
transform 1 0 32752 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_352
timestamp 28801
transform 1 0 33488 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_365
timestamp 1636997256
transform 1 0 34684 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_377
timestamp 1636997256
transform 1 0 35788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 28801
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 28801
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_415
timestamp 28801
transform 1 0 39284 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_430
timestamp 28801
transform 1 0 40664 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_438
timestamp 28801
transform 1 0 41400 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 28801
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_36
timestamp 28801
transform 1 0 4416 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_40
timestamp 28801
transform 1 0 4784 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_48
timestamp 28801
transform 1 0 5520 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_59
timestamp 28801
transform 1 0 6532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_67
timestamp 28801
transform 1 0 7268 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_78
timestamp 28801
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_48_85
timestamp 28801
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_109
timestamp 28801
transform 1 0 11132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_133
timestamp 28801
transform 1 0 13340 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 28801
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_173
timestamp 28801
transform 1 0 17020 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_181
timestamp 28801
transform 1 0 17756 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_202
timestamp 1636997256
transform 1 0 19688 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_214
timestamp 28801
transform 1 0 20792 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_231
timestamp 28801
transform 1 0 22356 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 28801
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1636997256
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_265
timestamp 28801
transform 1 0 25484 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_286
timestamp 1636997256
transform 1 0 27416 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_298
timestamp 28801
transform 1 0 28520 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_337
timestamp 1636997256
transform 1 0 32108 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_349
timestamp 28801
transform 1 0 33212 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_357
timestamp 28801
transform 1 0 33948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 28801
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_365
timestamp 28801
transform 1 0 34684 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_381
timestamp 1636997256
transform 1 0 36156 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_393
timestamp 28801
transform 1 0 37260 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_421
timestamp 28801
transform 1 0 39836 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 28801
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_39
timestamp 28801
transform 1 0 4692 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 28801
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_64
timestamp 28801
transform 1 0 6992 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_70
timestamp 1636997256
transform 1 0 7544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_82
timestamp 28801
transform 1 0 8648 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_90
timestamp 28801
transform 1 0 9384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 28801
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_138
timestamp 1636997256
transform 1 0 13800 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_150
timestamp 1636997256
transform 1 0 14904 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 28801
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_49_169
timestamp 28801
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 28801
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_208
timestamp 28801
transform 1 0 20240 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_212
timestamp 28801
transform 1 0 20608 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_216
timestamp 28801
transform 1 0 20976 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_233
timestamp 28801
transform 1 0 22540 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_255
timestamp 28801
transform 1 0 24564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_259
timestamp 28801
transform 1 0 24932 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 28801
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_285
timestamp 28801
transform 1 0 27324 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 28801
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_349
timestamp 28801
transform 1 0 33212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_365
timestamp 28801
transform 1 0 34684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_374
timestamp 28801
transform 1 0 35512 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 28801
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_421
timestamp 28801
transform 1 0 39836 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_442
timestamp 28801
transform 1 0 41768 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 28801
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_11
timestamp 28801
transform 1 0 2116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 28801
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_36
timestamp 28801
transform 1 0 4416 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_81
timestamp 28801
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_85
timestamp 28801
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_91
timestamp 28801
transform 1 0 9476 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_98
timestamp 1636997256
transform 1 0 10120 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 28801
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_156
timestamp 28801
transform 1 0 15456 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_164
timestamp 28801
transform 1 0 16192 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_188
timestamp 28801
transform 1 0 18400 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_213
timestamp 28801
transform 1 0 20700 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_235
timestamp 28801
transform 1 0 22724 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 28801
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_260
timestamp 28801
transform 1 0 25024 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_270
timestamp 28801
transform 1 0 25944 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1636997256
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_301
timestamp 28801
transform 1 0 28796 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_320
timestamp 28801
transform 1 0 30544 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_50_361
timestamp 28801
transform 1 0 34316 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_384
timestamp 28801
transform 1 0 36432 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_394
timestamp 1636997256
transform 1 0 37352 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_406
timestamp 28801
transform 1 0 38456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_410
timestamp 28801
transform 1 0 38824 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 28801
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 28801
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_11
timestamp 28801
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_27
timestamp 28801
transform 1 0 3588 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_33
timestamp 28801
transform 1 0 4140 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 28801
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_64
timestamp 1636997256
transform 1 0 6992 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_76
timestamp 28801
transform 1 0 8096 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_92
timestamp 28801
transform 1 0 9568 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_103
timestamp 28801
transform 1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 28801
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_113
timestamp 28801
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_144
timestamp 28801
transform 1 0 14352 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_184
timestamp 28801
transform 1 0 18032 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_193
timestamp 28801
transform 1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_211
timestamp 28801
transform 1 0 20516 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_233
timestamp 28801
transform 1 0 22540 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_239
timestamp 28801
transform 1 0 23092 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_260
timestamp 1636997256
transform 1 0 25024 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_272
timestamp 28801
transform 1 0 26128 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1636997256
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1636997256
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1636997256
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_317
timestamp 28801
transform 1 0 30268 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_337
timestamp 28801
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_348
timestamp 1636997256
transform 1 0 33120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_360
timestamp 28801
transform 1 0 34224 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_371
timestamp 28801
transform 1 0 35236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 28801
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_401
timestamp 28801
transform 1 0 37996 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_412
timestamp 28801
transform 1 0 39008 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_446
timestamp 28801
transform 1 0 42136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 28801
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_18
timestamp 28801
transform 1 0 2760 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 28801
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_46
timestamp 28801
transform 1 0 5336 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_58
timestamp 1636997256
transform 1 0 6440 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_70
timestamp 28801
transform 1 0 7544 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_75
timestamp 28801
transform 1 0 8004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_79
timestamp 28801
transform 1 0 8372 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_105
timestamp 1636997256
transform 1 0 10764 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_117
timestamp 28801
transform 1 0 11868 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 28801
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1636997256
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1636997256
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_165
timestamp 28801
transform 1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_180
timestamp 28801
transform 1 0 17664 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 28801
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_214
timestamp 28801
transform 1 0 20792 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_235
timestamp 28801
transform 1 0 22724 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 28801
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1636997256
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_265
timestamp 28801
transform 1 0 25484 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 28801
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_326
timestamp 28801
transform 1 0 31096 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_356
timestamp 28801
transform 1 0 33856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_365
timestamp 28801
transform 1 0 34684 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_378
timestamp 1636997256
transform 1 0 35880 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_390
timestamp 28801
transform 1 0 36984 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_398
timestamp 28801
transform 1 0 37720 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_415
timestamp 28801
transform 1 0 39284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 28801
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 28801
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 28801
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 28801
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_65
timestamp 28801
transform 1 0 7084 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_81
timestamp 28801
transform 1 0 8556 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_104
timestamp 28801
transform 1 0 10672 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_113
timestamp 28801
transform 1 0 11500 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_142
timestamp 28801
transform 1 0 14168 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_178
timestamp 28801
transform 1 0 17480 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_201
timestamp 1636997256
transform 1 0 19596 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_213
timestamp 28801
transform 1 0 20700 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 28801
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_234
timestamp 28801
transform 1 0 22632 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_242
timestamp 28801
transform 1 0 23368 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_252
timestamp 28801
transform 1 0 24288 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_267
timestamp 28801
transform 1 0 25668 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_298
timestamp 28801
transform 1 0 28520 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_317
timestamp 28801
transform 1 0 30268 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_346
timestamp 28801
transform 1 0 32936 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_367
timestamp 1636997256
transform 1 0 34868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_379
timestamp 1636997256
transform 1 0 35972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 28801
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_393
timestamp 28801
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_399
timestamp 28801
transform 1 0 37812 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_416
timestamp 28801
transform 1 0 39376 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_435
timestamp 28801
transform 1 0 41124 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_444
timestamp 28801
transform 1 0 41952 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636997256
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_15
timestamp 28801
transform 1 0 2484 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 28801
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 28801
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_37
timestamp 28801
transform 1 0 4508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_43
timestamp 28801
transform 1 0 5060 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_50
timestamp 28801
transform 1 0 5704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_58
timestamp 28801
transform 1 0 6440 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 28801
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 28801
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_115
timestamp 28801
transform 1 0 11684 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 28801
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_187
timestamp 28801
transform 1 0 18308 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 28801
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_206
timestamp 1636997256
transform 1 0 20056 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_218
timestamp 28801
transform 1 0 21160 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_231
timestamp 1636997256
transform 1 0 22356 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 28801
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 28801
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 28801
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_343
timestamp 28801
transform 1 0 32660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 28801
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_365
timestamp 28801
transform 1 0 34684 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_390
timestamp 28801
transform 1 0 36984 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_411
timestamp 28801
transform 1 0 38916 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_430
timestamp 28801
transform 1 0 40664 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_3
timestamp 28801
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_11
timestamp 28801
transform 1 0 2116 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_19
timestamp 28801
transform 1 0 2852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_29
timestamp 28801
transform 1 0 3772 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_33
timestamp 28801
transform 1 0 4140 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_46
timestamp 28801
transform 1 0 5336 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 28801
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_61
timestamp 1636997256
transform 1 0 6716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_77
timestamp 1636997256
transform 1 0 8188 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_89
timestamp 28801
transform 1 0 9292 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_95
timestamp 28801
transform 1 0 9844 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_99
timestamp 1636997256
transform 1 0 10212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 28801
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_113
timestamp 28801
transform 1 0 11500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_147
timestamp 28801
transform 1 0 14628 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 28801
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 28801
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_202
timestamp 28801
transform 1 0 19688 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_208
timestamp 28801
transform 1 0 20240 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 28801
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_225
timestamp 28801
transform 1 0 21804 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_258
timestamp 28801
transform 1 0 24840 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 28801
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_281
timestamp 28801
transform 1 0 26956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_287
timestamp 28801
transform 1 0 27508 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_322
timestamp 28801
transform 1 0 30728 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 28801
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_337
timestamp 28801
transform 1 0 32108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_343
timestamp 28801
transform 1 0 32660 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_360
timestamp 28801
transform 1 0 34224 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_387
timestamp 28801
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 28801
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_417
timestamp 28801
transform 1 0 39468 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_23
timestamp 28801
transform 1 0 3220 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_29
timestamp 28801
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_40
timestamp 28801
transform 1 0 4784 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 28801
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 28801
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 28801
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_163
timestamp 28801
transform 1 0 16100 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_183
timestamp 28801
transform 1 0 17940 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_187
timestamp 28801
transform 1 0 18308 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_197
timestamp 28801
transform 1 0 19228 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_242
timestamp 28801
transform 1 0 23368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 28801
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 28801
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_279
timestamp 28801
transform 1 0 26772 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 28801
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_309
timestamp 28801
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_56_323
timestamp 28801
transform 1 0 30820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_350
timestamp 28801
transform 1 0 33304 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 28801
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_365
timestamp 28801
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_385
timestamp 28801
transform 1 0 36524 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_415
timestamp 28801
transform 1 0 39284 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 28801
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_421
timestamp 28801
transform 1 0 39836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_425
timestamp 28801
transform 1 0 40204 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_442
timestamp 28801
transform 1 0 41768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_446
timestamp 28801
transform 1 0 42136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 28801
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_9
timestamp 28801
transform 1 0 1932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_20
timestamp 28801
transform 1 0 2944 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 28801
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636997256
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_69
timestamp 28801
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_86
timestamp 28801
transform 1 0 9016 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1636997256
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_149
timestamp 28801
transform 1 0 14812 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_157
timestamp 28801
transform 1 0 15548 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_185
timestamp 28801
transform 1 0 18124 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_195
timestamp 28801
transform 1 0 19044 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_212
timestamp 1636997256
transform 1 0 20608 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_233
timestamp 28801
transform 1 0 22540 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_239
timestamp 28801
transform 1 0 23092 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_256
timestamp 28801
transform 1 0 24656 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_266
timestamp 28801
transform 1 0 25576 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_290
timestamp 28801
transform 1 0 27784 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_300
timestamp 1636997256
transform 1 0 28704 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_312
timestamp 28801
transform 1 0 29808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_316
timestamp 28801
transform 1 0 30176 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 28801
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_343
timestamp 28801
transform 1 0 32660 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_370
timestamp 1636997256
transform 1 0 35144 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_382
timestamp 28801
transform 1 0 36248 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 28801
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_393
timestamp 28801
transform 1 0 37260 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_399
timestamp 28801
transform 1 0 37812 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_418
timestamp 28801
transform 1 0 39560 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636997256
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636997256
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 28801
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636997256
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_41
timestamp 28801
transform 1 0 4876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_49
timestamp 28801
transform 1 0 5612 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_56
timestamp 28801
transform 1 0 6256 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_60
timestamp 28801
transform 1 0 6624 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_81
timestamp 28801
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_116
timestamp 28801
transform 1 0 11776 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 28801
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_161
timestamp 28801
transform 1 0 15916 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_165
timestamp 28801
transform 1 0 16284 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_175
timestamp 1636997256
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_187
timestamp 28801
transform 1 0 18308 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 28801
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 28801
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 28801
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_289
timestamp 28801
transform 1 0 27692 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_300
timestamp 28801
transform 1 0 28704 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_58_309
timestamp 28801
transform 1 0 29532 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_315
timestamp 28801
transform 1 0 30084 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_356
timestamp 28801
transform 1 0 33856 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_365
timestamp 28801
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_388
timestamp 28801
transform 1 0 36800 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_392
timestamp 28801
transform 1 0 37168 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 28801
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 28801
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_421
timestamp 28801
transform 1 0 39836 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_442
timestamp 28801
transform 1 0 41768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_446
timestamp 28801
transform 1 0 42136 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636997256
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636997256
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_27
timestamp 28801
transform 1 0 3588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_33
timestamp 28801
transform 1 0 4140 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_41
timestamp 28801
transform 1 0 4876 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 28801
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636997256
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_69
timestamp 28801
transform 1 0 7452 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_90
timestamp 28801
transform 1 0 9384 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_121
timestamp 28801
transform 1 0 12236 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_127
timestamp 28801
transform 1 0 12788 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_148
timestamp 28801
transform 1 0 14720 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_200
timestamp 28801
transform 1 0 19504 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 28801
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 28801
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_229
timestamp 28801
transform 1 0 22172 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_255
timestamp 28801
transform 1 0 24564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 28801
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_281
timestamp 28801
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_296
timestamp 28801
transform 1 0 28336 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_306
timestamp 28801
transform 1 0 29256 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_310
timestamp 28801
transform 1 0 29624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 28801
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_445
timestamp 28801
transform 1 0 42044 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636997256
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_15
timestamp 28801
transform 1 0 2484 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_21
timestamp 28801
transform 1 0 3036 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 28801
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_42
timestamp 28801
transform 1 0 4968 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_70
timestamp 28801
transform 1 0 7544 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_74
timestamp 28801
transform 1 0 7912 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 28801
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1636997256
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1636997256
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1636997256
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_149
timestamp 28801
transform 1 0 14812 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_170
timestamp 28801
transform 1 0 16744 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_190
timestamp 28801
transform 1 0 18584 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_230
timestamp 28801
transform 1 0 22264 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 28801
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 28801
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 28801
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_257
timestamp 28801
transform 1 0 24748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_275
timestamp 28801
transform 1 0 26404 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_279
timestamp 28801
transform 1 0 26772 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 28801
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 28801
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_373
timestamp 28801
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_391
timestamp 28801
transform 1 0 37076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_416
timestamp 28801
transform 1 0 39376 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_421
timestamp 28801
transform 1 0 39836 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_441
timestamp 28801
transform 1 0 41676 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_446
timestamp 28801
transform 1 0 42136 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636997256
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_15
timestamp 28801
transform 1 0 2484 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_44
timestamp 28801
transform 1 0 5152 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 28801
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_65
timestamp 28801
transform 1 0 7084 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_87
timestamp 28801
transform 1 0 9108 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 28801
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 28801
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_169
timestamp 28801
transform 1 0 16652 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_200
timestamp 28801
transform 1 0 19504 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_225
timestamp 28801
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_246
timestamp 28801
transform 1 0 23736 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_252
timestamp 28801
transform 1 0 24288 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 28801
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 28801
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_289
timestamp 28801
transform 1 0 27692 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_301
timestamp 28801
transform 1 0 28796 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_309
timestamp 28801
transform 1 0 29532 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_321
timestamp 28801
transform 1 0 30636 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 28801
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_337
timestamp 28801
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_366
timestamp 28801
transform 1 0 34776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_383
timestamp 28801
transform 1 0 36340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 28801
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_393
timestamp 28801
transform 1 0 37260 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_406
timestamp 28801
transform 1 0 38456 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_438
timestamp 28801
transform 1 0 41400 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636997256
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636997256
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 28801
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_29
timestamp 28801
transform 1 0 3772 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_44
timestamp 28801
transform 1 0 5152 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_50
timestamp 28801
transform 1 0 5704 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_56
timestamp 28801
transform 1 0 6256 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 28801
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_105
timestamp 1636997256
transform 1 0 10764 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_117
timestamp 28801
transform 1 0 11868 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_149
timestamp 28801
transform 1 0 14812 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_205
timestamp 28801
transform 1 0 19964 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_220
timestamp 28801
transform 1 0 21344 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 28801
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_253
timestamp 28801
transform 1 0 24380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_259
timestamp 28801
transform 1 0 24932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_280
timestamp 28801
transform 1 0 26864 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_304
timestamp 28801
transform 1 0 29072 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_331
timestamp 28801
transform 1 0 31556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_337
timestamp 28801
transform 1 0 32108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_355
timestamp 28801
transform 1 0 33764 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 28801
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_373
timestamp 1636997256
transform 1 0 35420 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_421
timestamp 28801
transform 1 0 39836 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636997256
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636997256
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_27
timestamp 28801
transform 1 0 3588 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_49
timestamp 28801
transform 1 0 5612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 28801
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_57
timestamp 28801
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_65
timestamp 28801
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_77
timestamp 1636997256
transform 1 0 8188 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_89
timestamp 1636997256
transform 1 0 9292 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_101
timestamp 28801
transform 1 0 10396 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_109
timestamp 28801
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1636997256
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1636997256
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1636997256
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_149
timestamp 28801
transform 1 0 14812 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 28801
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_185
timestamp 28801
transform 1 0 18124 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_204
timestamp 28801
transform 1 0 19872 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 28801
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 28801
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_261
timestamp 28801
transform 1 0 25116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 28801
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_289
timestamp 28801
transform 1 0 27692 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_297
timestamp 28801
transform 1 0 28428 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_318
timestamp 28801
transform 1 0 30360 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_386
timestamp 28801
transform 1 0 36616 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_406
timestamp 28801
transform 1 0 38456 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_414
timestamp 28801
transform 1 0 39192 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_428
timestamp 28801
transform 1 0 40480 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636997256
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636997256
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 28801
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636997256
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1636997256
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1636997256
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1636997256
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 28801
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 28801
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1636997256
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1636997256
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1636997256
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_121
timestamp 28801
transform 1 0 12236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_129
timestamp 28801
transform 1 0 12972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_152
timestamp 28801
transform 1 0 15088 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_174
timestamp 28801
transform 1 0 17112 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_205
timestamp 28801
transform 1 0 19964 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_211
timestamp 28801
transform 1 0 20516 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_232
timestamp 28801
transform 1 0 22448 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 28801
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 28801
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_270
timestamp 28801
transform 1 0 25944 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_293
timestamp 1636997256
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 28801
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1636997256
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_321
timestamp 28801
transform 1 0 30636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_326
timestamp 28801
transform 1 0 31096 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_331
timestamp 28801
transform 1 0 31556 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_342
timestamp 28801
transform 1 0 32568 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 28801
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_365
timestamp 28801
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_372
timestamp 1636997256
transform 1 0 35328 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_384
timestamp 28801
transform 1 0 36432 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_392
timestamp 28801
transform 1 0 37168 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_397
timestamp 1636997256
transform 1 0 37628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_409
timestamp 28801
transform 1 0 38732 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 28801
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1636997256
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_433
timestamp 28801
transform 1 0 40940 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1636997256
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1636997256
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1636997256
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1636997256
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 28801
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 28801
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1636997256
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1636997256
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1636997256
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1636997256
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 28801
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 28801
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1636997256
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_125
timestamp 28801
transform 1 0 12604 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_153
timestamp 28801
transform 1 0 15180 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_157
timestamp 28801
transform 1 0 15548 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 28801
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_212
timestamp 28801
transform 1 0 20608 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 28801
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_231
timestamp 28801
transform 1 0 22356 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_240
timestamp 1636997256
transform 1 0 23184 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_252
timestamp 28801
transform 1 0 24288 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_260
timestamp 28801
transform 1 0 25024 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_266
timestamp 1636997256
transform 1 0 25576 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 28801
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_299
timestamp 28801
transform 1 0 28612 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_303
timestamp 28801
transform 1 0 28980 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_321
timestamp 1636997256
transform 1 0 30636 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_333
timestamp 28801
transform 1 0 31740 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_337
timestamp 28801
transform 1 0 32108 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_358
timestamp 1636997256
transform 1 0 34040 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_370
timestamp 28801
transform 1 0 35144 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_374
timestamp 28801
transform 1 0 35512 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_384
timestamp 28801
transform 1 0 36432 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_393
timestamp 28801
transform 1 0 37260 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_408
timestamp 1636997256
transform 1 0 38640 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_420
timestamp 28801
transform 1 0 39744 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_425
timestamp 28801
transform 1 0 40204 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_444
timestamp 28801
transform 1 0 41952 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636997256
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636997256
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 28801
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636997256
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1636997256
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1636997256
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1636997256
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 28801
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 28801
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1636997256
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1636997256
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1636997256
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1636997256
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 28801
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 28801
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_141
timestamp 28801
transform 1 0 14076 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_66_182
timestamp 28801
transform 1 0 17848 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 28801
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_197
timestamp 28801
transform 1 0 19228 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_205
timestamp 28801
transform 1 0 19964 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_217
timestamp 28801
transform 1 0 21068 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_231
timestamp 28801
transform 1 0 22356 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_240
timestamp 1636997256
transform 1 0 23184 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_256
timestamp 28801
transform 1 0 24656 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_272
timestamp 28801
transform 1 0 26128 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_289
timestamp 28801
transform 1 0 27692 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_305
timestamp 28801
transform 1 0 29164 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1636997256
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1636997256
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_333
timestamp 28801
transform 1 0 31740 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1636997256
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_357
timestamp 28801
transform 1 0 33948 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_408
timestamp 28801
transform 1 0 38640 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_426
timestamp 28801
transform 1 0 40296 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636997256
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636997256
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1636997256
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1636997256
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 28801
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 28801
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636997256
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1636997256
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1636997256
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1636997256
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 28801
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 28801
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1636997256
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1636997256
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_137
timestamp 28801
transform 1 0 13708 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_145
timestamp 28801
transform 1 0 14444 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_169
timestamp 28801
transform 1 0 16652 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_194
timestamp 28801
transform 1 0 18952 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_200
timestamp 28801
transform 1 0 19504 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_215
timestamp 28801
transform 1 0 20884 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_265
timestamp 28801
transform 1 0 25484 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_271
timestamp 28801
transform 1 0 26036 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 28801
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1636997256
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_305
timestamp 28801
transform 1 0 29164 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_313
timestamp 28801
transform 1 0 29900 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 28801
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 28801
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_387
timestamp 28801
transform 1 0 36708 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 28801
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_412
timestamp 28801
transform 1 0 39008 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_443
timestamp 28801
transform 1 0 41860 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636997256
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636997256
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 28801
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636997256
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636997256
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636997256
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1636997256
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 28801
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 28801
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1636997256
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1636997256
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1636997256
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1636997256
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 28801
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 28801
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1636997256
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1636997256
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1636997256
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1636997256
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1636997256
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1636997256
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_221
timestamp 28801
transform 1 0 21436 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_229
timestamp 28801
transform 1 0 22172 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 28801
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_267
timestamp 1636997256
transform 1 0 25668 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_279
timestamp 1636997256
transform 1 0 26772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_291
timestamp 1636997256
transform 1 0 27876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_303
timestamp 28801
transform 1 0 28980 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 28801
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_309
timestamp 28801
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_313
timestamp 28801
transform 1 0 29900 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_332
timestamp 28801
transform 1 0 31648 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_350
timestamp 28801
transform 1 0 33304 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_358
timestamp 28801
transform 1 0 34040 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_378
timestamp 1636997256
transform 1 0 35880 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_390
timestamp 28801
transform 1 0 36984 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_396
timestamp 1636997256
transform 1 0 37536 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_408
timestamp 28801
transform 1 0 38640 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_438
timestamp 28801
transform 1 0 41400 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636997256
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636997256
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636997256
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636997256
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 28801
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 28801
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636997256
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1636997256
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1636997256
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1636997256
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 28801
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 28801
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1636997256
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1636997256
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1636997256
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1636997256
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 28801
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 28801
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_194
timestamp 28801
transform 1 0 18952 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_69_209
timestamp 28801
transform 1 0 20332 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_218
timestamp 28801
transform 1 0 21160 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_232
timestamp 28801
transform 1 0 22448 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_236
timestamp 28801
transform 1 0 22816 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_253
timestamp 28801
transform 1 0 24380 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_258
timestamp 28801
transform 1 0 24840 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_266
timestamp 28801
transform 1 0 25576 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_281
timestamp 28801
transform 1 0 26956 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_289
timestamp 28801
transform 1 0 27692 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_297
timestamp 1636997256
transform 1 0 28428 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_309
timestamp 1636997256
transform 1 0 29532 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_321
timestamp 28801
transform 1 0 30636 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_326
timestamp 28801
transform 1 0 31096 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_334
timestamp 28801
transform 1 0 31832 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_341
timestamp 1636997256
transform 1 0 32476 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_353
timestamp 1636997256
transform 1 0 33580 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_365
timestamp 1636997256
transform 1 0 34684 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_377
timestamp 28801
transform 1 0 35788 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_383
timestamp 28801
transform 1 0 36340 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_390
timestamp 28801
transform 1 0 36984 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_393
timestamp 28801
transform 1 0 37260 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_401
timestamp 28801
transform 1 0 37996 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_424
timestamp 1636997256
transform 1 0 40112 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_436
timestamp 28801
transform 1 0 41216 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_444
timestamp 28801
transform 1 0 41952 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636997256
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636997256
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 28801
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636997256
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636997256
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636997256
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1636997256
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 28801
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 28801
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1636997256
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1636997256
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1636997256
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1636997256
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 28801
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 28801
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1636997256
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_153
timestamp 28801
transform 1 0 15180 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_175
timestamp 28801
transform 1 0 17204 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_194
timestamp 28801
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_222
timestamp 28801
transform 1 0 21528 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_230
timestamp 28801
transform 1 0 22264 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_238
timestamp 1636997256
transform 1 0 23000 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 28801
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_253
timestamp 28801
transform 1 0 24380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_70_267
timestamp 28801
transform 1 0 25668 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_276
timestamp 28801
transform 1 0 26496 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_284
timestamp 28801
transform 1 0 27232 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_309
timestamp 28801
transform 1 0 29532 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_324
timestamp 28801
transform 1 0 30912 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_331
timestamp 28801
transform 1 0 31556 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_339
timestamp 28801
transform 1 0 32292 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_352
timestamp 1636997256
transform 1 0 33488 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1636997256
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_377
timestamp 28801
transform 1 0 35788 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_399
timestamp 28801
transform 1 0 37812 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_403
timestamp 28801
transform 1 0 38180 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_417
timestamp 28801
transform 1 0 39468 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1636997256
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1636997256
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_445
timestamp 28801
transform 1 0 42044 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636997256
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636997256
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636997256
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636997256
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 28801
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 28801
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636997256
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1636997256
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1636997256
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1636997256
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 28801
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 28801
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1636997256
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1636997256
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1636997256
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1636997256
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_169
timestamp 28801
transform 1 0 16652 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_187
timestamp 1636997256
transform 1 0 18308 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_199
timestamp 28801
transform 1 0 19412 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 28801
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_225
timestamp 28801
transform 1 0 21804 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_231
timestamp 28801
transform 1 0 22356 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_241
timestamp 28801
transform 1 0 23276 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_251
timestamp 1636997256
transform 1 0 24196 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_263
timestamp 28801
transform 1 0 25300 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_267
timestamp 28801
transform 1 0 25668 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_276
timestamp 28801
transform 1 0 26496 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_281
timestamp 28801
transform 1 0 26956 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_289
timestamp 28801
transform 1 0 27692 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_344
timestamp 28801
transform 1 0 32752 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_356
timestamp 28801
transform 1 0 33856 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_360
timestamp 28801
transform 1 0 34224 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_379
timestamp 28801
transform 1 0 35972 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_387
timestamp 28801
transform 1 0 36708 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_428
timestamp 1636997256
transform 1 0 40480 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_440
timestamp 28801
transform 1 0 41584 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_446
timestamp 28801
transform 1 0 42136 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636997256
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636997256
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 28801
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636997256
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636997256
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636997256
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1636997256
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 28801
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 28801
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1636997256
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1636997256
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1636997256
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1636997256
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 28801
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 28801
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1636997256
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1636997256
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_165
timestamp 28801
transform 1 0 16284 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_191
timestamp 28801
transform 1 0 18676 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 28801
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_229
timestamp 28801
transform 1 0 22172 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 28801
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_282
timestamp 1636997256
transform 1 0 27048 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_302
timestamp 28801
transform 1 0 28888 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_309
timestamp 28801
transform 1 0 29532 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_335
timestamp 28801
transform 1 0 31924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_343
timestamp 28801
transform 1 0 32660 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_351
timestamp 28801
transform 1 0 33396 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 28801
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_374
timestamp 1636997256
transform 1 0 35512 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_386
timestamp 28801
transform 1 0 36616 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_394
timestamp 28801
transform 1 0 37352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_399
timestamp 28801
transform 1 0 37812 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1636997256
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1636997256
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_445
timestamp 28801
transform 1 0 42044 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636997256
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636997256
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636997256
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636997256
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 28801
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 28801
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636997256
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1636997256
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1636997256
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1636997256
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 28801
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 28801
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1636997256
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1636997256
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1636997256
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1636997256
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 28801
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 28801
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1636997256
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1636997256
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_193
timestamp 28801
transform 1 0 18860 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_225
timestamp 28801
transform 1 0 21804 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_249
timestamp 28801
transform 1 0 24012 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_284
timestamp 28801
transform 1 0 27232 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_305
timestamp 28801
transform 1 0 29164 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 28801
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_337
timestamp 28801
transform 1 0 32108 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_377
timestamp 1636997256
transform 1 0 35788 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_389
timestamp 28801
transform 1 0 36892 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_393
timestamp 28801
transform 1 0 37260 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_397
timestamp 28801
transform 1 0 37628 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_406
timestamp 28801
transform 1 0 38456 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_418
timestamp 1636997256
transform 1 0 39560 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_430
timestamp 1636997256
transform 1 0 40664 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_442
timestamp 28801
transform 1 0 41768 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_446
timestamp 28801
transform 1 0 42136 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636997256
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636997256
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 28801
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636997256
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636997256
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636997256
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1636997256
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 28801
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 28801
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1636997256
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1636997256
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1636997256
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1636997256
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 28801
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 28801
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1636997256
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1636997256
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1636997256
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1636997256
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 28801
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 28801
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_223
timestamp 28801
transform 1 0 21620 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_253
timestamp 28801
transform 1 0 24380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_261
timestamp 28801
transform 1 0 25116 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_280
timestamp 28801
transform 1 0 26864 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_302
timestamp 28801
transform 1 0 28888 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_74_361
timestamp 28801
transform 1 0 34316 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_373
timestamp 1636997256
transform 1 0 35420 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_385
timestamp 1636997256
transform 1 0 36524 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_397
timestamp 1636997256
transform 1 0 37628 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_409
timestamp 28801
transform 1 0 38732 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_417
timestamp 28801
transform 1 0 39468 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1636997256
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1636997256
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_445
timestamp 28801
transform 1 0 42044 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636997256
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636997256
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_27
timestamp 28801
transform 1 0 3588 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_29
timestamp 1636997256
transform 1 0 3772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_41
timestamp 1636997256
transform 1 0 4876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 28801
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636997256
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1636997256
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_81
timestamp 28801
transform 1 0 8556 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_85
timestamp 1636997256
transform 1 0 8924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_97
timestamp 1636997256
transform 1 0 10028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_109
timestamp 28801
transform 1 0 11132 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1636997256
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1636997256
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_137
timestamp 28801
transform 1 0 13708 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_141
timestamp 1636997256
transform 1 0 14076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_153
timestamp 1636997256
transform 1 0 15180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_165
timestamp 28801
transform 1 0 16284 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1636997256
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1636997256
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_193
timestamp 28801
transform 1 0 18860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_197
timestamp 28801
transform 1 0 19228 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_205
timestamp 28801
transform 1 0 19964 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_210
timestamp 28801
transform 1 0 20424 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_225
timestamp 28801
transform 1 0 21804 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_233
timestamp 28801
transform 1 0 22540 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_238
timestamp 28801
transform 1 0 23000 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_246
timestamp 28801
transform 1 0 23736 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_253
timestamp 1636997256
transform 1 0 24380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_265
timestamp 28801
transform 1 0 25484 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_277
timestamp 28801
transform 1 0 26588 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1636997256
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1636997256
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_305
timestamp 28801
transform 1 0 29164 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_309
timestamp 1636997256
transform 1 0 29532 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_321
timestamp 1636997256
transform 1 0 30636 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_333
timestamp 28801
transform 1 0 31740 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1636997256
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_349
timestamp 28801
transform 1 0 33212 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_363
timestamp 28801
transform 1 0 34500 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_365
timestamp 1636997256
transform 1 0 34684 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_377
timestamp 1636997256
transform 1 0 35788 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_389
timestamp 28801
transform 1 0 36892 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1636997256
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1636997256
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_417
timestamp 28801
transform 1 0 39468 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_421
timestamp 1636997256
transform 1 0 39836 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_433
timestamp 1636997256
transform 1 0 40940 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_445
timestamp 28801
transform 1 0 42044 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 28801
transform -1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 28801
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 28801
transform -1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 28801
transform -1 0 3036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 28801
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 28801
transform 1 0 31832 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 28801
transform -1 0 31096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 28801
transform -1 0 18584 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 28801
transform -1 0 42136 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 28801
transform -1 0 33948 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 28801
transform -1 0 23368 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 28801
transform -1 0 27692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 28801
transform -1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 28801
transform -1 0 3312 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 28801
transform -1 0 14996 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 28801
transform -1 0 25760 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 28801
transform 1 0 41308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 28801
transform 1 0 33304 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 28801
transform 1 0 38916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 28801
transform 1 0 17480 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 28801
transform -1 0 41952 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 28801
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 28801
transform -1 0 30820 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 28801
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 28801
transform -1 0 27692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 28801
transform -1 0 18216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 28801
transform 1 0 33304 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 28801
transform -1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 28801
transform -1 0 42228 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 28801
transform -1 0 13616 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 28801
transform -1 0 25944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 28801
transform 1 0 9016 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 28801
transform 1 0 37628 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 28801
transform -1 0 18676 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 28801
transform -1 0 41492 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 28801
transform -1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 28801
transform -1 0 17112 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 28801
transform -1 0 24196 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 28801
transform -1 0 16284 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 28801
transform -1 0 15456 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 28801
transform 1 0 3864 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 28801
transform 1 0 4600 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 28801
transform -1 0 41676 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 28801
transform -1 0 10028 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 28801
transform -1 0 42228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 28801
transform 1 0 19780 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 28801
transform -1 0 22540 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 28801
transform 1 0 17204 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 28801
transform -1 0 38732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 28801
transform -1 0 29348 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 28801
transform 1 0 41492 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 28801
transform -1 0 36708 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 28801
transform -1 0 29072 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 28801
transform -1 0 25300 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 28801
transform -1 0 14812 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 28801
transform -1 0 40480 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 28801
transform 1 0 37904 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 28801
transform -1 0 16008 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 28801
transform -1 0 42228 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 28801
transform -1 0 39652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 28801
transform -1 0 37904 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 28801
transform -1 0 29164 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 28801
transform -1 0 28428 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 28801
transform -1 0 26404 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 28801
transform -1 0 39284 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 28801
transform 1 0 40204 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 28801
transform -1 0 37168 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 28801
transform 1 0 20056 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 28801
transform -1 0 34868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 28801
transform -1 0 39468 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 28801
transform -1 0 26864 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 28801
transform 1 0 22264 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 28801
transform -1 0 39928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 28801
transform 1 0 37720 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 28801
transform 1 0 28244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 28801
transform -1 0 29348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 28801
transform -1 0 26404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 28801
transform 1 0 25760 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 28801
transform -1 0 21068 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 28801
transform -1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 28801
transform 1 0 31280 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 28801
transform 1 0 29808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 28801
transform -1 0 26220 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 28801
transform 1 0 24748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 28801
transform -1 0 4968 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 28801
transform 1 0 12236 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 28801
transform 1 0 21988 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 28801
transform -1 0 22540 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 28801
transform 1 0 15824 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 28801
transform -1 0 31740 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 28801
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 28801
transform 1 0 2300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 28801
transform -1 0 18860 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 28801
transform -1 0 30820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 28801
transform 1 0 29992 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 28801
transform 1 0 16008 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 28801
transform -1 0 27692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 28801
transform -1 0 25760 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 28801
transform -1 0 28888 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 28801
transform 1 0 23184 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 28801
transform -1 0 24656 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 28801
transform 1 0 12972 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 28801
transform -1 0 14628 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 28801
transform -1 0 33948 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 28801
transform 1 0 22540 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 28801
transform -1 0 39100 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 28801
transform -1 0 21068 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 28801
transform 1 0 19320 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 28801
transform -1 0 34040 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 28801
transform -1 0 13524 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 28801
transform 1 0 9568 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 28801
transform -1 0 19504 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 28801
transform -1 0 40848 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 28801
transform -1 0 41308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 28801
transform -1 0 11684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 28801
transform 1 0 34868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 28801
transform 1 0 14076 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 28801
transform -1 0 42228 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 28801
transform 1 0 28612 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 28801
transform -1 0 32844 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 28801
transform -1 0 19964 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 28801
transform 1 0 9752 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 28801
transform -1 0 40572 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 28801
transform -1 0 8832 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 28801
transform -1 0 39100 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 28801
transform -1 0 16560 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 28801
transform -1 0 41492 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 28801
transform 1 0 40204 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 28801
transform 1 0 25300 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 28801
transform -1 0 32108 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 28801
transform 1 0 19964 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 28801
transform -1 0 41860 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 28801
transform 1 0 23000 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 28801
transform -1 0 30360 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 28801
transform 1 0 32936 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 28801
transform -1 0 34408 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 28801
transform 1 0 34684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 28801
transform -1 0 34316 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 28801
transform 1 0 7544 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 28801
transform -1 0 35512 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 28801
transform -1 0 40020 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 28801
transform -1 0 14168 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 28801
transform -1 0 26680 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 28801
transform -1 0 25116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 28801
transform -1 0 33396 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 28801
transform -1 0 31832 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 28801
transform 1 0 33120 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 28801
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 28801
transform -1 0 17388 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 28801
transform -1 0 15732 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 28801
transform 1 0 16744 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 28801
transform -1 0 36248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 28801
transform -1 0 34592 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 28801
transform -1 0 10304 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 28801
transform -1 0 24196 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 28801
transform -1 0 21804 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 28801
transform -1 0 4048 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 28801
transform 1 0 38824 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 28801
transform -1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 28801
transform -1 0 27692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 28801
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 28801
transform -1 0 31556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 28801
transform -1 0 22816 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 28801
transform 1 0 23092 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 28801
transform -1 0 26588 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 28801
transform 1 0 22356 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 28801
transform -1 0 22540 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 28801
transform -1 0 34500 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 28801
transform 1 0 40848 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 28801
transform -1 0 41032 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 28801
transform -1 0 42228 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 28801
transform -1 0 30084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 28801
transform -1 0 30268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 28801
transform -1 0 42228 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 28801
transform -1 0 30820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 28801
transform -1 0 41860 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 28801
transform 1 0 40388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 28801
transform -1 0 21620 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 28801
transform -1 0 25944 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 28801
transform -1 0 33672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 28801
transform -1 0 32660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 28801
transform -1 0 36984 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 28801
transform -1 0 17664 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 28801
transform -1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 28801
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 28801
transform -1 0 36524 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 28801
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 28801
transform -1 0 41952 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 28801
transform -1 0 40848 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 28801
transform -1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 28801
transform -1 0 8556 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 28801
transform -1 0 35236 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 28801
transform -1 0 13984 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 28801
transform -1 0 29164 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 28801
transform -1 0 26588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 28801
transform -1 0 41400 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 28801
transform 1 0 34684 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 28801
transform -1 0 31096 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 28801
transform 1 0 35512 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 28801
transform -1 0 38456 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 28801
transform -1 0 42228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 28801
transform -1 0 34408 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 28801
transform -1 0 9844 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 28801
transform -1 0 24288 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 28801
transform -1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 28801
transform -1 0 31924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 28801
transform -1 0 31740 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 28801
transform -1 0 35420 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 28801
transform -1 0 15640 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 28801
transform 1 0 32660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 28801
transform -1 0 28428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 28801
transform 1 0 28428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 28801
transform -1 0 32108 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 28801
transform 1 0 35604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 28801
transform -1 0 11684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 28801
transform -1 0 21804 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 28801
transform 1 0 26128 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 28801
transform -1 0 23736 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 28801
transform -1 0 39284 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 28801
transform -1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 28801
transform -1 0 36524 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 28801
transform -1 0 24288 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 28801
transform -1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 28801
transform -1 0 26864 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 28801
transform 1 0 22540 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 28801
transform -1 0 39652 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 28801
transform -1 0 21712 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 28801
transform -1 0 37260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 28801
transform -1 0 9016 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 28801
transform -1 0 22172 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 28801
transform 1 0 30452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 28801
transform -1 0 27508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 28801
transform 1 0 27048 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 28801
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 28801
transform 1 0 19136 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 28801
transform -1 0 31648 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 28801
transform -1 0 25116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 28801
transform -1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 28801
transform 1 0 35144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 28801
transform -1 0 26220 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 28801
transform -1 0 11224 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 28801
transform -1 0 3956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 28801
transform -1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 28801
transform -1 0 27692 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 28801
transform -1 0 40572 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 28801
transform -1 0 37260 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 28801
transform -1 0 20700 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 28801
transform -1 0 19136 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 28801
transform -1 0 34500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 28801
transform -1 0 11316 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 28801
transform -1 0 10856 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 28801
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 28801
transform -1 0 7084 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 28801
transform -1 0 17388 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 28801
transform -1 0 39376 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 28801
transform -1 0 33304 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 28801
transform -1 0 12236 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 28801
transform -1 0 9752 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 28801
transform -1 0 11316 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 28801
transform -1 0 29440 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 28801
transform 1 0 39008 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 28801
transform -1 0 37076 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 28801
transform -1 0 13340 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 28801
transform 1 0 9200 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 28801
transform -1 0 6624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 28801
transform -1 0 3956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 28801
transform -1 0 4232 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 28801
transform 1 0 11316 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 28801
transform -1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 28801
transform -1 0 19964 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 28801
transform -1 0 3496 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 28801
transform -1 0 12236 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 28801
transform -1 0 9660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 28801
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 28801
transform 1 0 15364 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 28801
transform -1 0 23184 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 28801
transform -1 0 37076 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 28801
transform -1 0 17388 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 28801
transform -1 0 34684 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 28801
transform -1 0 30452 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 28801
transform -1 0 14812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 28801
transform -1 0 18308 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 28801
transform -1 0 30636 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 28801
transform -1 0 37904 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 28801
transform -1 0 30268 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 28801
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 28801
transform -1 0 24748 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 28801
transform -1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 28801
transform -1 0 27692 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 28801
transform -1 0 9016 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 28801
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 28801
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 28801
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 28801
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 28801
transform -1 0 42228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap75
timestamp 28801
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 28801
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 28801
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 28801
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 28801
transform -1 0 3588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 28801
transform -1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 28801
transform -1 0 21068 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 28801
transform 1 0 41768 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 28801
transform -1 0 39836 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 28801
transform 1 0 41860 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 28801
transform 1 0 41308 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 28801
transform 1 0 41860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 28801
transform 1 0 20056 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 28801
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 28801
transform -1 0 23000 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 28801
transform -1 0 24288 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 28801
transform 1 0 41308 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 28801
transform 1 0 41492 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 28801
transform 1 0 40020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 28801
transform 1 0 41860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 28801
transform 1 0 41860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 28801
transform 1 0 41860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 28801
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 28801
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 28801
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 28801
transform -1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_76
timestamp 28801
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 28801
transform -1 0 42504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_77
timestamp 28801
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 28801
transform -1 0 42504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_78
timestamp 28801
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 28801
transform -1 0 42504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_79
timestamp 28801
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 28801
transform -1 0 42504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_80
timestamp 28801
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 28801
transform -1 0 42504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_81
timestamp 28801
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 28801
transform -1 0 42504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_82
timestamp 28801
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 28801
transform -1 0 42504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_83
timestamp 28801
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 28801
transform -1 0 42504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_84
timestamp 28801
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 28801
transform -1 0 42504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_85
timestamp 28801
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 28801
transform -1 0 42504 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_86
timestamp 28801
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 28801
transform -1 0 42504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_87
timestamp 28801
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 28801
transform -1 0 42504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_88
timestamp 28801
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 28801
transform -1 0 42504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_89
timestamp 28801
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 28801
transform -1 0 42504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_90
timestamp 28801
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 28801
transform -1 0 42504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_91
timestamp 28801
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 28801
transform -1 0 42504 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_92
timestamp 28801
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 28801
transform -1 0 42504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_93
timestamp 28801
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 28801
transform -1 0 42504 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_94
timestamp 28801
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 28801
transform -1 0 42504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_95
timestamp 28801
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 28801
transform -1 0 42504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_96
timestamp 28801
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 28801
transform -1 0 42504 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_97
timestamp 28801
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 28801
transform -1 0 42504 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_98
timestamp 28801
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 28801
transform -1 0 42504 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_99
timestamp 28801
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 28801
transform -1 0 42504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_100
timestamp 28801
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 28801
transform -1 0 42504 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_101
timestamp 28801
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 28801
transform -1 0 42504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_102
timestamp 28801
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 28801
transform -1 0 42504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_103
timestamp 28801
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 28801
transform -1 0 42504 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_104
timestamp 28801
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 28801
transform -1 0 42504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_105
timestamp 28801
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 28801
transform -1 0 42504 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_106
timestamp 28801
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 28801
transform -1 0 42504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_107
timestamp 28801
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 28801
transform -1 0 42504 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_108
timestamp 28801
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 28801
transform -1 0 42504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_109
timestamp 28801
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 28801
transform -1 0 42504 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_110
timestamp 28801
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 28801
transform -1 0 42504 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_111
timestamp 28801
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 28801
transform -1 0 42504 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_112
timestamp 28801
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 28801
transform -1 0 42504 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_113
timestamp 28801
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 28801
transform -1 0 42504 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_114
timestamp 28801
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 28801
transform -1 0 42504 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_115
timestamp 28801
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 28801
transform -1 0 42504 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_116
timestamp 28801
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 28801
transform -1 0 42504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_117
timestamp 28801
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 28801
transform -1 0 42504 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_118
timestamp 28801
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 28801
transform -1 0 42504 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_119
timestamp 28801
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 28801
transform -1 0 42504 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_120
timestamp 28801
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 28801
transform -1 0 42504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_121
timestamp 28801
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 28801
transform -1 0 42504 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_122
timestamp 28801
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 28801
transform -1 0 42504 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_123
timestamp 28801
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 28801
transform -1 0 42504 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_124
timestamp 28801
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 28801
transform -1 0 42504 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_125
timestamp 28801
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 28801
transform -1 0 42504 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_126
timestamp 28801
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 28801
transform -1 0 42504 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_127
timestamp 28801
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 28801
transform -1 0 42504 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_128
timestamp 28801
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 28801
transform -1 0 42504 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_129
timestamp 28801
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 28801
transform -1 0 42504 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_130
timestamp 28801
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 28801
transform -1 0 42504 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_131
timestamp 28801
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 28801
transform -1 0 42504 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_132
timestamp 28801
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 28801
transform -1 0 42504 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_133
timestamp 28801
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 28801
transform -1 0 42504 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_134
timestamp 28801
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 28801
transform -1 0 42504 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_135
timestamp 28801
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 28801
transform -1 0 42504 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_136
timestamp 28801
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 28801
transform -1 0 42504 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_137
timestamp 28801
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 28801
transform -1 0 42504 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_138
timestamp 28801
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 28801
transform -1 0 42504 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_139
timestamp 28801
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 28801
transform -1 0 42504 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_140
timestamp 28801
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 28801
transform -1 0 42504 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_141
timestamp 28801
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 28801
transform -1 0 42504 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_142
timestamp 28801
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 28801
transform -1 0 42504 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_143
timestamp 28801
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 28801
transform -1 0 42504 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_144
timestamp 28801
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 28801
transform -1 0 42504 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_145
timestamp 28801
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 28801
transform -1 0 42504 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_146
timestamp 28801
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 28801
transform -1 0 42504 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_147
timestamp 28801
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 28801
transform -1 0 42504 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_148
timestamp 28801
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 28801
transform -1 0 42504 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_149
timestamp 28801
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 28801
transform -1 0 42504 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_150
timestamp 28801
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 28801
transform -1 0 42504 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_151
timestamp 28801
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 28801
transform -1 0 42504 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_152
timestamp 28801
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_153
timestamp 28801
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_154
timestamp 28801
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_155
timestamp 28801
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_156
timestamp 28801
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_157
timestamp 28801
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_158
timestamp 28801
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_159
timestamp 28801
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_160
timestamp 28801
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_161
timestamp 28801
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_162
timestamp 28801
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_163
timestamp 28801
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_164
timestamp 28801
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_165
timestamp 28801
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_166
timestamp 28801
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_167
timestamp 28801
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_168
timestamp 28801
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_169
timestamp 28801
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_170
timestamp 28801
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_171
timestamp 28801
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_172
timestamp 28801
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_173
timestamp 28801
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_174
timestamp 28801
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_175
timestamp 28801
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_176
timestamp 28801
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_177
timestamp 28801
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_178
timestamp 28801
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_179
timestamp 28801
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_180
timestamp 28801
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_181
timestamp 28801
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_182
timestamp 28801
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_183
timestamp 28801
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_184
timestamp 28801
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_185
timestamp 28801
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_186
timestamp 28801
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_187
timestamp 28801
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_188
timestamp 28801
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_189
timestamp 28801
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_190
timestamp 28801
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_191
timestamp 28801
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_192
timestamp 28801
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_193
timestamp 28801
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_194
timestamp 28801
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_195
timestamp 28801
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_196
timestamp 28801
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_197
timestamp 28801
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_198
timestamp 28801
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_199
timestamp 28801
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_200
timestamp 28801
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_201
timestamp 28801
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_202
timestamp 28801
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_203
timestamp 28801
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_204
timestamp 28801
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_205
timestamp 28801
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_206
timestamp 28801
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_207
timestamp 28801
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_208
timestamp 28801
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_209
timestamp 28801
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_210
timestamp 28801
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_211
timestamp 28801
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_212
timestamp 28801
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_213
timestamp 28801
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_214
timestamp 28801
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_215
timestamp 28801
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_216
timestamp 28801
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_217
timestamp 28801
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_218
timestamp 28801
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_219
timestamp 28801
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_220
timestamp 28801
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_221
timestamp 28801
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_222
timestamp 28801
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_223
timestamp 28801
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_224
timestamp 28801
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_225
timestamp 28801
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_226
timestamp 28801
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_227
timestamp 28801
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_228
timestamp 28801
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_229
timestamp 28801
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_230
timestamp 28801
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_231
timestamp 28801
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_232
timestamp 28801
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_233
timestamp 28801
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_234
timestamp 28801
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_235
timestamp 28801
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_236
timestamp 28801
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_237
timestamp 28801
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_238
timestamp 28801
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_239
timestamp 28801
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_240
timestamp 28801
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_241
timestamp 28801
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_242
timestamp 28801
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_243
timestamp 28801
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_244
timestamp 28801
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_245
timestamp 28801
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_246
timestamp 28801
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_247
timestamp 28801
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_248
timestamp 28801
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_249
timestamp 28801
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_250
timestamp 28801
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_251
timestamp 28801
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_252
timestamp 28801
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_253
timestamp 28801
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_254
timestamp 28801
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_255
timestamp 28801
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_256
timestamp 28801
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_257
timestamp 28801
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_258
timestamp 28801
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_259
timestamp 28801
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_260
timestamp 28801
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_261
timestamp 28801
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_262
timestamp 28801
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_263
timestamp 28801
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_264
timestamp 28801
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_265
timestamp 28801
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_266
timestamp 28801
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_267
timestamp 28801
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_268
timestamp 28801
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_269
timestamp 28801
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_270
timestamp 28801
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_271
timestamp 28801
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_272
timestamp 28801
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_273
timestamp 28801
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_274
timestamp 28801
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_275
timestamp 28801
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_276
timestamp 28801
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_277
timestamp 28801
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_278
timestamp 28801
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_279
timestamp 28801
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_280
timestamp 28801
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_281
timestamp 28801
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_282
timestamp 28801
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_283
timestamp 28801
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_284
timestamp 28801
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_285
timestamp 28801
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_286
timestamp 28801
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_287
timestamp 28801
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_288
timestamp 28801
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_289
timestamp 28801
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_290
timestamp 28801
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_291
timestamp 28801
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_292
timestamp 28801
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_293
timestamp 28801
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_294
timestamp 28801
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_295
timestamp 28801
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_296
timestamp 28801
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_297
timestamp 28801
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_298
timestamp 28801
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_299
timestamp 28801
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_300
timestamp 28801
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_301
timestamp 28801
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_302
timestamp 28801
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_303
timestamp 28801
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_304
timestamp 28801
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_305
timestamp 28801
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_306
timestamp 28801
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_307
timestamp 28801
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_308
timestamp 28801
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_309
timestamp 28801
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_310
timestamp 28801
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_311
timestamp 28801
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_312
timestamp 28801
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_313
timestamp 28801
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_314
timestamp 28801
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_315
timestamp 28801
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_316
timestamp 28801
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_317
timestamp 28801
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_318
timestamp 28801
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_319
timestamp 28801
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_320
timestamp 28801
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_321
timestamp 28801
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_322
timestamp 28801
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_323
timestamp 28801
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_324
timestamp 28801
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_325
timestamp 28801
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_326
timestamp 28801
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_327
timestamp 28801
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_328
timestamp 28801
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_329
timestamp 28801
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_330
timestamp 28801
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_331
timestamp 28801
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_332
timestamp 28801
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_333
timestamp 28801
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_334
timestamp 28801
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_335
timestamp 28801
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_336
timestamp 28801
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_337
timestamp 28801
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_338
timestamp 28801
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_339
timestamp 28801
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_340
timestamp 28801
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_341
timestamp 28801
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_342
timestamp 28801
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_343
timestamp 28801
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_344
timestamp 28801
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_345
timestamp 28801
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_346
timestamp 28801
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_347
timestamp 28801
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_348
timestamp 28801
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_349
timestamp 28801
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_350
timestamp 28801
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_351
timestamp 28801
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_352
timestamp 28801
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_353
timestamp 28801
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_354
timestamp 28801
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_355
timestamp 28801
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_356
timestamp 28801
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_357
timestamp 28801
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_358
timestamp 28801
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_359
timestamp 28801
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_360
timestamp 28801
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_361
timestamp 28801
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_362
timestamp 28801
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_363
timestamp 28801
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_364
timestamp 28801
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_365
timestamp 28801
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_366
timestamp 28801
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_367
timestamp 28801
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_368
timestamp 28801
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_369
timestamp 28801
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_370
timestamp 28801
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_371
timestamp 28801
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_372
timestamp 28801
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_373
timestamp 28801
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_374
timestamp 28801
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_375
timestamp 28801
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_376
timestamp 28801
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_377
timestamp 28801
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_378
timestamp 28801
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_379
timestamp 28801
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_380
timestamp 28801
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_381
timestamp 28801
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_382
timestamp 28801
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_383
timestamp 28801
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_384
timestamp 28801
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_385
timestamp 28801
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_386
timestamp 28801
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_387
timestamp 28801
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_388
timestamp 28801
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_389
timestamp 28801
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_390
timestamp 28801
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_391
timestamp 28801
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_392
timestamp 28801
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_393
timestamp 28801
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_394
timestamp 28801
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_395
timestamp 28801
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_396
timestamp 28801
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_397
timestamp 28801
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_398
timestamp 28801
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_399
timestamp 28801
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_400
timestamp 28801
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_401
timestamp 28801
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_402
timestamp 28801
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_403
timestamp 28801
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_404
timestamp 28801
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_405
timestamp 28801
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_406
timestamp 28801
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_407
timestamp 28801
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_408
timestamp 28801
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_409
timestamp 28801
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_410
timestamp 28801
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_411
timestamp 28801
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_412
timestamp 28801
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_413
timestamp 28801
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_414
timestamp 28801
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_415
timestamp 28801
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_416
timestamp 28801
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_417
timestamp 28801
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_418
timestamp 28801
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_419
timestamp 28801
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_420
timestamp 28801
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_421
timestamp 28801
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_422
timestamp 28801
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_423
timestamp 28801
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_424
timestamp 28801
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_425
timestamp 28801
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_426
timestamp 28801
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_427
timestamp 28801
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_428
timestamp 28801
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_429
timestamp 28801
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_430
timestamp 28801
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_431
timestamp 28801
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_432
timestamp 28801
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_433
timestamp 28801
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_434
timestamp 28801
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_435
timestamp 28801
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_436
timestamp 28801
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_437
timestamp 28801
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_438
timestamp 28801
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_439
timestamp 28801
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_440
timestamp 28801
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_441
timestamp 28801
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_442
timestamp 28801
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_443
timestamp 28801
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_444
timestamp 28801
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_445
timestamp 28801
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_446
timestamp 28801
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_447
timestamp 28801
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_448
timestamp 28801
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_449
timestamp 28801
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_450
timestamp 28801
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_451
timestamp 28801
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_452
timestamp 28801
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_453
timestamp 28801
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_454
timestamp 28801
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_455
timestamp 28801
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_456
timestamp 28801
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_457
timestamp 28801
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_458
timestamp 28801
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_459
timestamp 28801
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_460
timestamp 28801
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_461
timestamp 28801
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_462
timestamp 28801
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_463
timestamp 28801
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_464
timestamp 28801
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_465
timestamp 28801
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_466
timestamp 28801
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_467
timestamp 28801
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_468
timestamp 28801
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_469
timestamp 28801
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_470
timestamp 28801
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_471
timestamp 28801
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_472
timestamp 28801
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_473
timestamp 28801
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_474
timestamp 28801
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_475
timestamp 28801
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_476
timestamp 28801
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_477
timestamp 28801
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_478
timestamp 28801
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_479
timestamp 28801
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_480
timestamp 28801
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_481
timestamp 28801
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_482
timestamp 28801
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_483
timestamp 28801
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_484
timestamp 28801
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_485
timestamp 28801
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_486
timestamp 28801
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_487
timestamp 28801
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_488
timestamp 28801
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_489
timestamp 28801
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_490
timestamp 28801
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_491
timestamp 28801
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_492
timestamp 28801
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_493
timestamp 28801
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_494
timestamp 28801
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_495
timestamp 28801
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_496
timestamp 28801
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_497
timestamp 28801
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_498
timestamp 28801
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_499
timestamp 28801
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_500
timestamp 28801
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_501
timestamp 28801
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_502
timestamp 28801
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_503
timestamp 28801
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_504
timestamp 28801
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_505
timestamp 28801
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_506
timestamp 28801
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_507
timestamp 28801
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_508
timestamp 28801
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_509
timestamp 28801
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_510
timestamp 28801
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_511
timestamp 28801
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_512
timestamp 28801
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_513
timestamp 28801
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_514
timestamp 28801
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_515
timestamp 28801
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_516
timestamp 28801
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_517
timestamp 28801
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_518
timestamp 28801
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_519
timestamp 28801
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_520
timestamp 28801
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_521
timestamp 28801
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_522
timestamp 28801
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_523
timestamp 28801
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_524
timestamp 28801
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_525
timestamp 28801
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_526
timestamp 28801
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_527
timestamp 28801
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_528
timestamp 28801
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_529
timestamp 28801
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_530
timestamp 28801
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_531
timestamp 28801
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_532
timestamp 28801
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_533
timestamp 28801
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_534
timestamp 28801
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_535
timestamp 28801
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_536
timestamp 28801
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_537
timestamp 28801
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_538
timestamp 28801
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_539
timestamp 28801
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_540
timestamp 28801
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_541
timestamp 28801
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_542
timestamp 28801
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_543
timestamp 28801
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_544
timestamp 28801
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_545
timestamp 28801
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_546
timestamp 28801
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_547
timestamp 28801
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_548
timestamp 28801
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_549
timestamp 28801
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_550
timestamp 28801
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_551
timestamp 28801
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_552
timestamp 28801
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_553
timestamp 28801
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_554
timestamp 28801
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_555
timestamp 28801
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_556
timestamp 28801
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_557
timestamp 28801
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_558
timestamp 28801
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_559
timestamp 28801
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_560
timestamp 28801
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_561
timestamp 28801
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_562
timestamp 28801
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_563
timestamp 28801
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_564
timestamp 28801
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_565
timestamp 28801
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_566
timestamp 28801
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_567
timestamp 28801
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_568
timestamp 28801
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_569
timestamp 28801
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_570
timestamp 28801
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_571
timestamp 28801
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_572
timestamp 28801
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_573
timestamp 28801
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_574
timestamp 28801
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_575
timestamp 28801
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_576
timestamp 28801
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_577
timestamp 28801
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_578
timestamp 28801
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_579
timestamp 28801
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_580
timestamp 28801
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_581
timestamp 28801
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_582
timestamp 28801
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_583
timestamp 28801
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_584
timestamp 28801
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_585
timestamp 28801
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_586
timestamp 28801
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_587
timestamp 28801
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_588
timestamp 28801
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_589
timestamp 28801
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_590
timestamp 28801
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_591
timestamp 28801
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_592
timestamp 28801
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_593
timestamp 28801
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_594
timestamp 28801
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_595
timestamp 28801
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_596
timestamp 28801
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_597
timestamp 28801
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_598
timestamp 28801
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_599
timestamp 28801
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_600
timestamp 28801
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_601
timestamp 28801
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_602
timestamp 28801
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_603
timestamp 28801
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_604
timestamp 28801
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_605
timestamp 28801
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_606
timestamp 28801
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_607
timestamp 28801
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_608
timestamp 28801
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_609
timestamp 28801
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_610
timestamp 28801
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_611
timestamp 28801
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_612
timestamp 28801
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_613
timestamp 28801
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_614
timestamp 28801
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_615
timestamp 28801
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_616
timestamp 28801
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_617
timestamp 28801
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_618
timestamp 28801
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_619
timestamp 28801
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_620
timestamp 28801
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_621
timestamp 28801
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_622
timestamp 28801
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_623
timestamp 28801
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_624
timestamp 28801
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_625
timestamp 28801
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_626
timestamp 28801
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_627
timestamp 28801
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_628
timestamp 28801
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_629
timestamp 28801
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_630
timestamp 28801
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_631
timestamp 28801
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_632
timestamp 28801
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_633
timestamp 28801
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_634
timestamp 28801
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_635
timestamp 28801
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_636
timestamp 28801
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_637
timestamp 28801
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_638
timestamp 28801
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_639
timestamp 28801
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_640
timestamp 28801
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_641
timestamp 28801
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_642
timestamp 28801
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_643
timestamp 28801
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_644
timestamp 28801
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_645
timestamp 28801
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_646
timestamp 28801
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_647
timestamp 28801
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_648
timestamp 28801
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_649
timestamp 28801
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_650
timestamp 28801
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_651
timestamp 28801
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_652
timestamp 28801
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_653
timestamp 28801
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_654
timestamp 28801
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_655
timestamp 28801
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_656
timestamp 28801
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_657
timestamp 28801
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_658
timestamp 28801
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_659
timestamp 28801
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_660
timestamp 28801
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_661
timestamp 28801
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_662
timestamp 28801
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_663
timestamp 28801
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_664
timestamp 28801
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_665
timestamp 28801
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_666
timestamp 28801
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_667
timestamp 28801
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_668
timestamp 28801
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_669
timestamp 28801
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_670
timestamp 28801
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_671
timestamp 28801
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_672
timestamp 28801
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_673
timestamp 28801
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_674
timestamp 28801
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_675
timestamp 28801
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_676
timestamp 28801
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_677
timestamp 28801
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_678
timestamp 28801
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_679
timestamp 28801
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_680
timestamp 28801
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_681
timestamp 28801
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_682
timestamp 28801
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_683
timestamp 28801
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_684
timestamp 28801
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_685
timestamp 28801
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_686
timestamp 28801
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_687
timestamp 28801
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_688
timestamp 28801
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_689
timestamp 28801
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_690
timestamp 28801
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_691
timestamp 28801
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_692
timestamp 28801
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_693
timestamp 28801
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_694
timestamp 28801
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_695
timestamp 28801
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_696
timestamp 28801
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_697
timestamp 28801
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_698
timestamp 28801
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_699
timestamp 28801
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_700
timestamp 28801
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_701
timestamp 28801
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_702
timestamp 28801
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_703
timestamp 28801
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_704
timestamp 28801
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_705
timestamp 28801
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_706
timestamp 28801
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_707
timestamp 28801
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_708
timestamp 28801
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_709
timestamp 28801
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_710
timestamp 28801
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_711
timestamp 28801
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_712
timestamp 28801
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_713
timestamp 28801
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_714
timestamp 28801
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_715
timestamp 28801
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_716
timestamp 28801
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_717
timestamp 28801
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_718
timestamp 28801
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_719
timestamp 28801
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_720
timestamp 28801
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_721
timestamp 28801
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_722
timestamp 28801
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_723
timestamp 28801
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_724
timestamp 28801
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_725
timestamp 28801
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_726
timestamp 28801
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_727
timestamp 28801
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_728
timestamp 28801
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_729
timestamp 28801
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_730
timestamp 28801
transform 1 0 24288 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_731
timestamp 28801
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_732
timestamp 28801
transform 1 0 29440 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_733
timestamp 28801
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_734
timestamp 28801
transform 1 0 34592 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_735
timestamp 28801
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_736
timestamp 28801
transform 1 0 39744 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire84
timestamp 28801
transform 1 0 4048 0 -1 23936
box -38 -48 314 592
<< labels >>
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 ColOut[0]
port 0 nsew signal output
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 ColOut[1]
port 1 nsew signal output
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 ColOut[2]
port 2 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ColOut[3]
port 3 nsew signal output
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 RowIn[0]
port 4 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 RowIn[1]
port 5 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 RowIn[2]
port 6 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 RowIn[3]
port 7 nsew signal input
flabel metal4 s 4868 2128 5188 43568 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 43568 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal5 s 1056 6006 42552 6326 0 FreeSans 2560 0 0 0 VGND
port 8 nsew ground bidirectional
flabel metal5 s 1056 36642 42552 36962 0 FreeSans 2560 0 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 43568 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal4 s 34928 2128 35248 43568 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal5 s 1056 5346 42552 5666 0 FreeSans 2560 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal5 s 1056 35982 42552 36302 0 FreeSans 2560 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal3 s 0 42168 800 42288 0 FreeSans 480 0 0 0 clk
port 10 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 complete
port 11 nsew signal output
flabel metal2 s 20626 44957 20682 45757 0 FreeSans 224 90 0 0 display_output[0]
port 12 nsew signal output
flabel metal3 s 42813 29928 43613 30048 0 FreeSans 480 0 0 0 display_output[10]
port 13 nsew signal output
flabel metal3 s 42813 23128 43613 23248 0 FreeSans 480 0 0 0 display_output[11]
port 14 nsew signal output
flabel metal3 s 42813 29248 43613 29368 0 FreeSans 480 0 0 0 display_output[12]
port 15 nsew signal output
flabel metal3 s 42813 25168 43613 25288 0 FreeSans 480 0 0 0 display_output[13]
port 16 nsew signal output
flabel metal3 s 42813 28568 43613 28688 0 FreeSans 480 0 0 0 display_output[14]
port 17 nsew signal output
flabel metal2 s 19982 44957 20038 45757 0 FreeSans 224 90 0 0 display_output[15]
port 18 nsew signal output
flabel metal2 s 21270 44957 21326 45757 0 FreeSans 224 90 0 0 display_output[1]
port 19 nsew signal output
flabel metal2 s 22558 44957 22614 45757 0 FreeSans 224 90 0 0 display_output[2]
port 20 nsew signal output
flabel metal2 s 23846 44957 23902 45757 0 FreeSans 224 90 0 0 display_output[3]
port 21 nsew signal output
flabel metal3 s 42813 24488 43613 24608 0 FreeSans 480 0 0 0 display_output[4]
port 22 nsew signal output
flabel metal3 s 42813 27888 43613 28008 0 FreeSans 480 0 0 0 display_output[5]
port 23 nsew signal output
flabel metal3 s 42813 23808 43613 23928 0 FreeSans 480 0 0 0 display_output[6]
port 24 nsew signal output
flabel metal3 s 42813 27208 43613 27328 0 FreeSans 480 0 0 0 display_output[7]
port 25 nsew signal output
flabel metal3 s 42813 25848 43613 25968 0 FreeSans 480 0 0 0 display_output[8]
port 26 nsew signal output
flabel metal3 s 42813 26528 43613 26648 0 FreeSans 480 0 0 0 display_output[9]
port 27 nsew signal output
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 input_state_FPGA[0]
port 28 nsew signal output
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 input_state_FPGA[1]
port 29 nsew signal output
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 input_state_FPGA[2]
port 30 nsew signal output
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 key_pressed
port 31 nsew signal output
flabel metal3 s 42813 5448 43613 5568 0 FreeSans 480 0 0 0 nRST
port 32 nsew signal input
rlabel metal1 21804 43520 21804 43520 0 VGND
rlabel metal1 21804 42976 21804 42976 0 VPWR
rlabel metal2 11638 1520 11638 1520 0 ColOut[0]
rlabel metal1 1380 10778 1380 10778 0 ColOut[1]
rlabel metal3 1096 12988 1096 12988 0 ColOut[2]
rlabel metal2 3358 11849 3358 11849 0 ColOut[3]
rlabel metal3 1050 15028 1050 15028 0 RowIn[0]
rlabel metal3 751 15708 751 15708 0 RowIn[1]
rlabel metal3 751 17068 751 17068 0 RowIn[2]
rlabel metal3 1050 17748 1050 17748 0 RowIn[3]
rlabel metal2 12282 35428 12282 35428 0 _0000_
rlabel metal1 13892 35734 13892 35734 0 _0001_
rlabel metal2 16146 11594 16146 11594 0 _0002_
rlabel metal1 16744 11798 16744 11798 0 _0003_
rlabel metal1 30912 12410 30912 12410 0 _0004_
rlabel metal2 12558 34680 12558 34680 0 _0005_
rlabel metal2 27600 12580 27600 12580 0 _0006_
rlabel metal1 28152 12070 28152 12070 0 _0007_
rlabel metal1 6762 29546 6762 29546 0 _0008_
rlabel metal1 4002 36346 4002 36346 0 _0009_
rlabel metal1 3082 35258 3082 35258 0 _0010_
rlabel metal1 4692 33082 4692 33082 0 _0011_
rlabel metal1 6624 32538 6624 32538 0 _0012_
rlabel metal1 4554 30906 4554 30906 0 _0013_
rlabel metal1 2852 32538 2852 32538 0 _0014_
rlabel metal2 2070 31008 2070 31008 0 _0015_
rlabel metal1 1886 28594 1886 28594 0 _0016_
rlabel metal2 2898 28730 2898 28730 0 _0017_
rlabel metal1 7222 31450 7222 31450 0 _0018_
rlabel metal1 9062 30362 9062 30362 0 _0019_
rlabel metal1 9384 31450 9384 31450 0 _0020_
rlabel metal2 9522 33252 9522 33252 0 _0021_
rlabel metal2 9706 34272 9706 34272 0 _0022_
rlabel metal1 7314 33082 7314 33082 0 _0023_
rlabel metal2 8418 35938 8418 35938 0 _0024_
rlabel metal1 10212 35802 10212 35802 0 _0025_
rlabel metal2 5566 35292 5566 35292 0 _0026_
rlabel metal2 4646 23936 4646 23936 0 _0027_
rlabel metal2 6762 21284 6762 21284 0 _0028_
rlabel metal1 4692 21590 4692 21590 0 _0029_
rlabel metal1 4600 21658 4600 21658 0 _0030_
rlabel metal1 6808 20842 6808 20842 0 _0031_
rlabel metal1 6808 18870 6808 18870 0 _0032_
rlabel metal1 9000 19754 9000 19754 0 _0033_
rlabel metal2 9798 20706 9798 20706 0 _0034_
rlabel metal1 10253 19414 10253 19414 0 _0035_
rlabel metal2 12282 19618 12282 19618 0 _0036_
rlabel metal1 12231 20502 12231 20502 0 _0037_
rlabel via1 14218 18326 14218 18326 0 _0038_
rlabel metal2 13938 17170 13938 17170 0 _0039_
rlabel metal2 13294 16966 13294 16966 0 _0040_
rlabel metal2 13846 15878 13846 15878 0 _0041_
rlabel metal1 13018 15096 13018 15096 0 _0042_
rlabel metal1 10978 15402 10978 15402 0 _0043_
rlabel metal1 9144 14382 9144 14382 0 _0044_
rlabel metal1 8602 14960 8602 14960 0 _0045_
rlabel metal1 8096 16762 8096 16762 0 _0046_
rlabel metal2 7498 17442 7498 17442 0 _0047_
rlabel metal1 4278 19278 4278 19278 0 _0048_
rlabel metal1 2640 19754 2640 19754 0 _0049_
rlabel metal1 1840 19482 1840 19482 0 _0050_
rlabel metal1 3128 20570 3128 20570 0 _0051_
rlabel metal1 7774 22474 7774 22474 0 _0052_
rlabel via1 10253 23766 10253 23766 0 _0053_
rlabel metal1 10340 23086 10340 23086 0 _0054_
rlabel metal1 10058 24106 10058 24106 0 _0055_
rlabel metal1 8004 27574 8004 27574 0 _0056_
rlabel metal1 10400 25942 10400 25942 0 _0057_
rlabel metal2 9522 26758 9522 26758 0 _0058_
rlabel metal1 9062 27574 9062 27574 0 _0059_
rlabel metal1 20844 6970 20844 6970 0 _0060_
rlabel metal1 19366 8058 19366 8058 0 _0061_
rlabel metal1 23552 9622 23552 9622 0 _0062_
rlabel metal2 22402 5372 22402 5372 0 _0063_
rlabel metal1 24794 7276 24794 7276 0 _0064_
rlabel metal1 25806 8364 25806 8364 0 _0065_
rlabel metal1 29440 6970 29440 6970 0 _0066_
rlabel metal1 30222 5746 30222 5746 0 _0067_
rlabel metal1 30038 7276 30038 7276 0 _0068_
rlabel metal2 31510 5406 31510 5406 0 _0069_
rlabel metal2 34270 8670 34270 8670 0 _0070_
rlabel metal2 34730 5780 34730 5780 0 _0071_
rlabel metal2 37398 6460 37398 6460 0 _0072_
rlabel metal1 37766 9044 37766 9044 0 _0073_
rlabel metal1 38824 9622 38824 9622 0 _0074_
rlabel metal1 6440 15538 6440 15538 0 _0075_
rlabel metal1 4324 13498 4324 13498 0 _0076_
rlabel metal1 7498 12954 7498 12954 0 _0077_
rlabel metal1 5004 14586 5004 14586 0 _0078_
rlabel metal1 3818 11050 3818 11050 0 _0079_
rlabel metal1 2162 10778 2162 10778 0 _0080_
rlabel metal1 1702 12410 1702 12410 0 _0081_
rlabel metal1 2254 11016 2254 11016 0 _0082_
rlabel metal2 1702 9112 1702 9112 0 _0083_
rlabel metal1 2990 8364 2990 8364 0 _0084_
rlabel metal2 1794 7650 1794 7650 0 _0085_
rlabel metal2 1702 6494 1702 6494 0 _0086_
rlabel metal2 3266 5542 3266 5542 0 _0087_
rlabel metal2 4094 5508 4094 5508 0 _0088_
rlabel metal1 4232 6222 4232 6222 0 _0089_
rlabel metal2 6210 5372 6210 5372 0 _0090_
rlabel metal1 7268 6358 7268 6358 0 _0091_
rlabel metal1 8096 4794 8096 4794 0 _0092_
rlabel metal2 10810 5950 10810 5950 0 _0093_
rlabel metal1 9154 8398 9154 8398 0 _0094_
rlabel metal1 10021 9146 10021 9146 0 _0095_
rlabel metal1 14214 8398 14214 8398 0 _0096_
rlabel metal1 13294 7514 13294 7514 0 _0097_
rlabel metal1 10665 6970 10665 6970 0 _0098_
rlabel metal1 9098 11322 9098 11322 0 _0099_
rlabel metal1 14766 10098 14766 10098 0 _0100_
rlabel metal2 15502 11118 15502 11118 0 _0101_
rlabel metal1 11730 10234 11730 10234 0 _0102_
rlabel metal1 14582 12410 14582 12410 0 _0103_
rlabel metal1 12282 12682 12282 12682 0 _0104_
rlabel metal2 9890 14144 9890 14144 0 _0105_
rlabel metal1 10120 12614 10120 12614 0 _0106_
rlabel metal1 16882 30906 16882 30906 0 _0107_
rlabel metal1 19228 30566 19228 30566 0 _0108_
rlabel via1 21199 29818 21199 29818 0 _0109_
rlabel metal1 24794 29818 24794 29818 0 _0110_
rlabel metal1 24600 27642 24600 27642 0 _0111_
rlabel metal2 26266 30430 26266 30430 0 _0112_
rlabel metal1 28474 27370 28474 27370 0 _0113_
rlabel metal2 28566 29410 28566 29410 0 _0114_
rlabel metal1 30176 26554 30176 26554 0 _0115_
rlabel metal1 32055 27642 32055 27642 0 _0116_
rlabel metal1 37444 29206 37444 29206 0 _0117_
rlabel metal1 36110 27370 36110 27370 0 _0118_
rlabel metal1 35328 30906 35328 30906 0 _0119_
rlabel metal1 34592 27030 34592 27030 0 _0120_
rlabel metal1 32430 30362 32430 30362 0 _0121_
rlabel via1 17519 22202 17519 22202 0 _0122_
rlabel metal2 18814 22814 18814 22814 0 _0123_
rlabel metal2 21850 24412 21850 24412 0 _0124_
rlabel metal1 22586 23834 22586 23834 0 _0125_
rlabel metal1 24932 26010 24932 26010 0 _0126_
rlabel metal1 24610 23800 24610 23800 0 _0127_
rlabel metal1 27094 23834 27094 23834 0 _0128_
rlabel metal1 28060 25466 28060 25466 0 _0129_
rlabel metal1 30360 24378 30360 24378 0 _0130_
rlabel metal1 34086 24922 34086 24922 0 _0131_
rlabel metal2 37306 24412 37306 24412 0 _0132_
rlabel metal2 37582 23902 37582 23902 0 _0133_
rlabel metal1 36747 22202 36747 22202 0 _0134_
rlabel metal2 34914 22814 34914 22814 0 _0135_
rlabel metal2 30314 22814 30314 22814 0 _0136_
rlabel metal1 9522 21658 9522 21658 0 _0137_
rlabel metal1 18906 7174 18906 7174 0 _0138_
rlabel metal1 18439 9146 18439 9146 0 _0139_
rlabel metal1 20930 10098 20930 10098 0 _0140_
rlabel metal1 22954 5882 22954 5882 0 _0141_
rlabel metal2 23506 6426 23506 6426 0 _0142_
rlabel metal2 24610 9316 24610 9316 0 _0143_
rlabel metal1 26765 6970 26765 6970 0 _0144_
rlabel metal2 28474 5610 28474 5610 0 _0145_
rlabel metal2 29762 8670 29762 8670 0 _0146_
rlabel metal1 31924 5746 31924 5746 0 _0147_
rlabel metal1 32292 8058 32292 8058 0 _0148_
rlabel metal1 33895 6970 33895 6970 0 _0149_
rlabel metal2 35466 6528 35466 6528 0 _0150_
rlabel metal2 35926 8075 35926 8075 0 _0151_
rlabel metal1 37950 10132 37950 10132 0 _0152_
rlabel metal1 15410 35258 15410 35258 0 _0153_
rlabel metal1 16238 19482 16238 19482 0 _0154_
rlabel metal2 18354 19108 18354 19108 0 _0155_
rlabel metal1 18860 17850 18860 17850 0 _0156_
rlabel metal2 20746 19108 20746 19108 0 _0157_
rlabel metal2 22494 13090 22494 13090 0 _0158_
rlabel metal1 24288 18938 24288 18938 0 _0159_
rlabel metal2 25622 13634 25622 13634 0 _0160_
rlabel metal2 26910 19992 26910 19992 0 _0161_
rlabel metal1 28382 18938 28382 18938 0 _0162_
rlabel metal2 30498 19108 30498 19108 0 _0163_
rlabel metal1 33304 18394 33304 18394 0 _0164_
rlabel metal1 35604 18394 35604 18394 0 _0165_
rlabel metal1 35604 17850 35604 17850 0 _0166_
rlabel metal1 35742 15130 35742 15130 0 _0167_
rlabel metal1 36156 12954 36156 12954 0 _0168_
rlabel metal2 30498 13396 30498 13396 0 _0169_
rlabel metal2 17342 20196 17342 20196 0 _0170_
rlabel metal1 19044 13430 19044 13430 0 _0171_
rlabel metal1 17664 15538 17664 15538 0 _0172_
rlabel metal2 22218 17306 22218 17306 0 _0173_
rlabel metal2 23138 14348 23138 14348 0 _0174_
rlabel metal1 25070 16660 25070 16660 0 _0175_
rlabel metal2 25300 13430 25300 13430 0 _0176_
rlabel metal1 28290 13430 28290 13430 0 _0177_
rlabel metal1 29210 17306 29210 17306 0 _0178_
rlabel metal1 31694 17068 31694 17068 0 _0179_
rlabel metal1 35098 17238 35098 17238 0 _0180_
rlabel metal2 41630 18292 41630 18292 0 _0181_
rlabel metal1 40434 17068 40434 17068 0 _0182_
rlabel metal1 40158 14450 40158 14450 0 _0183_
rlabel metal1 40802 12206 40802 12206 0 _0184_
rlabel metal1 34362 13396 34362 13396 0 _0185_
rlabel metal1 16974 13226 16974 13226 0 _0186_
rlabel metal2 16238 14552 16238 14552 0 _0187_
rlabel metal1 16514 16626 16514 16626 0 _0188_
rlabel metal2 22034 20060 22034 20060 0 _0189_
rlabel metal2 22770 19108 22770 19108 0 _0190_
rlabel metal1 23460 20502 23460 20502 0 _0191_
rlabel metal2 25530 17884 25530 17884 0 _0192_
rlabel metal2 27278 16286 27278 16286 0 _0193_
rlabel metal1 28888 20366 28888 20366 0 _0194_
rlabel metal1 33810 19278 33810 19278 0 _0195_
rlabel metal2 38502 19618 38502 19618 0 _0196_
rlabel metal2 40250 19618 40250 19618 0 _0197_
rlabel metal1 40940 20570 40940 20570 0 _0198_
rlabel metal1 37388 15674 37388 15674 0 _0199_
rlabel metal2 40710 13532 40710 13532 0 _0200_
rlabel metal2 32246 14620 32246 14620 0 _0201_
rlabel metal2 19182 12036 19182 12036 0 _0202_
rlabel metal2 18630 10846 18630 10846 0 _0203_
rlabel metal2 22218 12274 22218 12274 0 _0204_
rlabel metal1 22632 11322 22632 11322 0 _0205_
rlabel metal2 24518 11934 24518 11934 0 _0206_
rlabel metal1 25392 10778 25392 10778 0 _0207_
rlabel metal2 26542 10268 26542 10268 0 _0208_
rlabel metal2 30130 10268 30130 10268 0 _0209_
rlabel metal2 29854 11288 29854 11288 0 _0210_
rlabel metal1 32660 12614 32660 12614 0 _0211_
rlabel metal1 32338 10778 32338 10778 0 _0212_
rlabel metal1 34546 10132 34546 10132 0 _0213_
rlabel metal2 36110 11390 36110 11390 0 _0214_
rlabel metal2 34822 11934 34822 11934 0 _0215_
rlabel metal1 33120 11798 33120 11798 0 _0216_
rlabel metal1 17473 13702 17473 13702 0 _0217_
rlabel metal1 18676 16014 18676 16014 0 _0218_
rlabel metal2 20838 16932 20838 16932 0 _0219_
rlabel metal1 20838 13362 20838 13362 0 _0220_
rlabel metal1 23138 17034 23138 17034 0 _0221_
rlabel metal2 24150 14382 24150 14382 0 _0222_
rlabel metal2 29854 14654 29854 14654 0 _0223_
rlabel metal1 27646 17306 27646 17306 0 _0224_
rlabel metal1 31326 16218 31326 16218 0 _0225_
rlabel metal2 33810 16286 33810 16286 0 _0226_
rlabel metal1 37904 17306 37904 17306 0 _0227_
rlabel metal1 38318 17306 38318 17306 0 _0228_
rlabel metal1 37904 14586 37904 14586 0 _0229_
rlabel metal1 39698 12886 39698 12886 0 _0230_
rlabel metal2 36478 14382 36478 14382 0 _0231_
rlabel metal2 15318 36312 15318 36312 0 _0232_
rlabel metal2 15962 23256 15962 23256 0 _0233_
rlabel metal2 17618 37468 17618 37468 0 _0234_
rlabel metal2 19090 38046 19090 38046 0 _0235_
rlabel metal2 20930 37468 20930 37468 0 _0236_
rlabel metal2 22494 38692 22494 38692 0 _0237_
rlabel metal2 25346 36312 25346 36312 0 _0238_
rlabel metal2 26542 37468 26542 37468 0 _0239_
rlabel metal1 27922 35802 27922 35802 0 _0240_
rlabel metal2 28842 37162 28842 37162 0 _0241_
rlabel metal2 23414 36652 23414 36652 0 _0242_
rlabel metal2 32154 38658 32154 38658 0 _0243_
rlabel metal1 35558 37978 35558 37978 0 _0244_
rlabel metal1 34355 38726 34355 38726 0 _0245_
rlabel metal1 35328 33898 35328 33898 0 _0246_
rlabel metal1 34960 34646 34960 34646 0 _0247_
rlabel metal1 32338 36346 32338 36346 0 _0248_
rlabel metal1 17848 36210 17848 36210 0 _0249_
rlabel metal1 16606 38522 16606 38522 0 _0250_
rlabel metal1 16192 40154 16192 40154 0 _0251_
rlabel metal2 19550 42092 19550 42092 0 _0252_
rlabel metal2 22034 41922 22034 41922 0 _0253_
rlabel metal1 23644 36822 23644 36822 0 _0254_
rlabel metal2 24610 42398 24610 42398 0 _0255_
rlabel metal1 27370 34714 27370 34714 0 _0256_
rlabel metal1 29900 42330 29900 42330 0 _0257_
rlabel metal2 33166 42602 33166 42602 0 _0258_
rlabel metal1 39330 41242 39330 41242 0 _0259_
rlabel metal1 40894 38386 40894 38386 0 _0260_
rlabel metal1 40020 35258 40020 35258 0 _0261_
rlabel metal2 37582 34408 37582 34408 0 _0262_
rlabel metal1 33166 34034 33166 34034 0 _0263_
rlabel metal2 29854 35292 29854 35292 0 _0264_
rlabel metal1 15410 37978 15410 37978 0 _0265_
rlabel metal1 17342 41242 17342 41242 0 _0266_
rlabel metal1 19780 42262 19780 42262 0 _0267_
rlabel metal1 22586 41786 22586 41786 0 _0268_
rlabel metal1 24794 35258 24794 35258 0 _0269_
rlabel metal1 25576 41650 25576 41650 0 _0270_
rlabel metal2 27646 42466 27646 42466 0 _0271_
rlabel metal1 30084 40698 30084 40698 0 _0272_
rlabel metal2 34730 41956 34730 41956 0 _0273_
rlabel metal1 36793 40698 36793 40698 0 _0274_
rlabel metal1 39652 38998 39652 38998 0 _0275_
rlabel metal2 40710 36380 40710 36380 0 _0276_
rlabel metal1 37628 34646 37628 34646 0 _0277_
rlabel metal2 32430 35292 32430 35292 0 _0278_
rlabel metal1 30176 33626 30176 33626 0 _0279_
rlabel metal1 14030 34170 14030 34170 0 _0280_
rlabel metal1 16187 15402 16187 15402 0 _0281_
rlabel metal1 16279 17646 16279 17646 0 _0282_
rlabel metal1 21523 20842 21523 20842 0 _0283_
rlabel metal2 23138 22406 23138 22406 0 _0284_
rlabel metal1 24007 21590 24007 21590 0 _0285_
rlabel metal1 25801 18734 25801 18734 0 _0286_
rlabel metal1 27411 21522 27411 21522 0 _0287_
rlabel metal2 29578 21726 29578 21726 0 _0288_
rlabel metal1 32522 19720 32522 19720 0 _0289_
rlabel metal1 38175 20434 38175 20434 0 _0290_
rlabel metal1 39739 20434 39739 20434 0 _0291_
rlabel metal1 40475 21522 40475 21522 0 _0292_
rlabel via1 37577 20910 37577 20910 0 _0293_
rlabel via1 40153 21930 40153 21930 0 _0294_
rlabel metal1 30907 15062 30907 15062 0 _0295_
rlabel metal1 15175 20502 15175 20502 0 _0296_
rlabel metal1 14168 31994 14168 31994 0 _0297_
rlabel metal1 13478 23630 13478 23630 0 _0298_
rlabel metal1 12093 21590 12093 21590 0 _0299_
rlabel metal1 13294 24072 13294 24072 0 _0300_
rlabel metal1 11403 32878 11403 32878 0 _0301_
rlabel metal2 16422 34374 16422 34374 0 _0302_
rlabel metal1 18461 34646 18461 34646 0 _0303_
rlabel metal1 20373 34646 20373 34646 0 _0304_
rlabel metal1 24150 33490 24150 33490 0 _0305_
rlabel metal2 24794 33762 24794 33762 0 _0306_
rlabel metal2 25806 32538 25806 32538 0 _0307_
rlabel metal2 28290 30940 28290 30940 0 _0308_
rlabel metal1 29343 32402 29343 32402 0 _0309_
rlabel metal1 32108 31450 32108 31450 0 _0310_
rlabel metal1 40112 30362 40112 30362 0 _0311_
rlabel metal1 39928 31994 39928 31994 0 _0312_
rlabel metal2 40986 33116 40986 33116 0 _0313_
rlabel metal2 38134 32402 38134 32402 0 _0314_
rlabel metal1 33529 31790 33529 31790 0 _0315_
rlabel metal1 30217 31790 30217 31790 0 _0316_
rlabel metal2 14490 31586 14490 31586 0 _0317_
rlabel metal2 17250 33286 17250 33286 0 _0318_
rlabel metal1 17567 35054 17567 35054 0 _0319_
rlabel metal1 20879 34986 20879 34986 0 _0320_
rlabel metal1 23142 34646 23142 34646 0 _0321_
rlabel metal2 24886 31586 24886 31586 0 _0322_
rlabel metal1 26128 31450 26128 31450 0 _0323_
rlabel metal1 27554 32266 27554 32266 0 _0324_
rlabel metal2 29578 31110 29578 31110 0 _0325_
rlabel metal1 34909 32402 34909 32402 0 _0326_
rlabel metal2 38226 30498 38226 30498 0 _0327_
rlabel metal2 40986 30838 40986 30838 0 _0328_
rlabel via1 40245 33490 40245 33490 0 _0329_
rlabel metal1 37352 31994 37352 31994 0 _0330_
rlabel metal1 33207 32402 33207 32402 0 _0331_
rlabel metal2 31970 31586 31970 31586 0 _0332_
rlabel metal2 15594 32198 15594 32198 0 _0333_
rlabel via1 12829 21998 12829 21998 0 _0334_
rlabel metal2 12650 31076 12650 31076 0 _0335_
rlabel metal1 11960 29274 11960 29274 0 _0336_
rlabel metal2 13110 29988 13110 29988 0 _0337_
rlabel metal1 10166 28186 10166 28186 0 _0338_
rlabel metal2 11546 26112 11546 26112 0 _0339_
rlabel metal1 11362 27098 11362 27098 0 _0340_
rlabel metal2 11546 28288 11546 28288 0 _0341_
rlabel metal1 14398 22678 14398 22678 0 _0342_
rlabel metal2 16330 29988 16330 29988 0 _0343_
rlabel metal1 13754 26418 13754 26418 0 _0344_
rlabel metal2 19826 33762 19826 33762 0 _0345_
rlabel metal2 21390 32640 21390 32640 0 _0346_
rlabel metal2 21482 32402 21482 32402 0 _0347_
rlabel metal1 24426 32334 24426 32334 0 _0348_
rlabel metal1 40756 24242 40756 24242 0 _0349_
rlabel metal1 38226 28424 38226 28424 0 _0350_
rlabel metal2 39790 23902 39790 23902 0 _0351_
rlabel metal1 40519 27642 40519 27642 0 _0352_
rlabel metal2 37582 26078 37582 26078 0 _0353_
rlabel metal2 40710 26588 40710 26588 0 _0354_
rlabel metal1 40526 29818 40526 29818 0 _0355_
rlabel metal1 40342 23154 40342 23154 0 _0356_
rlabel metal1 40526 29682 40526 29682 0 _0357_
rlabel metal2 39146 25262 39146 25262 0 _0358_
rlabel metal2 40710 28798 40710 28798 0 _0359_
rlabel metal2 18170 32878 18170 32878 0 _0360_
rlabel metal1 18400 20978 18400 20978 0 _0361_
rlabel metal1 19320 20026 19320 20026 0 _0362_
rlabel metal1 20373 21930 20373 21930 0 _0363_
rlabel via1 21753 21998 21753 21998 0 _0364_
rlabel metal2 25622 21794 25622 21794 0 _0365_
rlabel metal1 26664 21930 26664 21930 0 _0366_
rlabel metal1 26266 20570 26266 20570 0 _0367_
rlabel metal1 29072 21114 29072 21114 0 _0368_
rlabel metal2 31142 21386 31142 21386 0 _0369_
rlabel metal2 32430 21794 32430 21794 0 _0370_
rlabel metal1 34684 22202 34684 22202 0 _0371_
rlabel metal1 35788 20026 35788 20026 0 _0372_
rlabel metal1 36160 20910 36160 20910 0 _0373_
rlabel metal1 34904 19822 34904 19822 0 _0374_
rlabel metal1 33207 20910 33207 20910 0 _0375_
rlabel metal2 15042 21692 15042 21692 0 _0376_
rlabel via1 15405 14994 15405 14994 0 _0377_
rlabel metal2 22862 27319 22862 27319 0 _0378_
rlabel metal2 17986 26758 17986 26758 0 _0379_
rlabel metal1 16928 26350 16928 26350 0 _0380_
rlabel metal1 16192 26010 16192 26010 0 _0381_
rlabel metal1 16560 26418 16560 26418 0 _0382_
rlabel metal2 16698 25500 16698 25500 0 _0383_
rlabel metal1 12650 29070 12650 29070 0 _0384_
rlabel metal2 13570 29308 13570 29308 0 _0385_
rlabel metal1 13524 29274 13524 29274 0 _0386_
rlabel metal1 20378 26860 20378 26860 0 _0387_
rlabel metal1 18768 26758 18768 26758 0 _0388_
rlabel via1 14858 25670 14858 25670 0 _0389_
rlabel metal2 14950 26214 14950 26214 0 _0390_
rlabel metal1 14996 26554 14996 26554 0 _0391_
rlabel metal2 13938 29478 13938 29478 0 _0392_
rlabel via2 14766 26027 14766 26027 0 _0393_
rlabel metal2 15042 27744 15042 27744 0 _0394_
rlabel metal1 15272 25874 15272 25874 0 _0395_
rlabel metal1 16422 26554 16422 26554 0 _0396_
rlabel metal1 6256 11798 6256 11798 0 _0397_
rlabel metal1 7314 10574 7314 10574 0 _0398_
rlabel metal1 5014 10030 5014 10030 0 _0399_
rlabel metal2 6026 7582 6026 7582 0 _0400_
rlabel metal1 5980 8466 5980 8466 0 _0401_
rlabel metal1 6854 8942 6854 8942 0 _0402_
rlabel metal1 6532 8466 6532 8466 0 _0403_
rlabel metal1 6532 8942 6532 8942 0 _0404_
rlabel metal2 9430 7786 9430 7786 0 _0405_
rlabel metal1 10902 8568 10902 8568 0 _0406_
rlabel metal2 7498 9316 7498 9316 0 _0407_
rlabel metal1 6532 8602 6532 8602 0 _0408_
rlabel metal1 6210 9690 6210 9690 0 _0409_
rlabel metal1 6026 9588 6026 9588 0 _0410_
rlabel metal1 7130 9452 7130 9452 0 _0411_
rlabel metal1 8464 8058 8464 8058 0 _0412_
rlabel metal1 11454 8330 11454 8330 0 _0413_
rlabel metal1 7682 9010 7682 9010 0 _0414_
rlabel metal1 6624 9146 6624 9146 0 _0415_
rlabel metal2 8510 10302 8510 10302 0 _0416_
rlabel metal2 12834 12002 12834 12002 0 _0417_
rlabel metal1 9844 10438 9844 10438 0 _0418_
rlabel metal1 5796 10234 5796 10234 0 _0419_
rlabel metal1 5704 10642 5704 10642 0 _0420_
rlabel metal2 5566 9758 5566 9758 0 _0421_
rlabel metal1 4370 8058 4370 8058 0 _0422_
rlabel metal2 5658 7174 5658 7174 0 _0423_
rlabel metal2 5934 9180 5934 9180 0 _0424_
rlabel metal1 6256 8602 6256 8602 0 _0425_
rlabel metal1 6210 9010 6210 9010 0 _0426_
rlabel metal1 6808 10030 6808 10030 0 _0427_
rlabel metal1 11868 11118 11868 11118 0 _0428_
rlabel metal2 7406 10336 7406 10336 0 _0429_
rlabel metal1 8602 11084 8602 11084 0 _0430_
rlabel metal1 8924 10778 8924 10778 0 _0431_
rlabel metal2 7406 11220 7406 11220 0 _0432_
rlabel metal1 5382 12750 5382 12750 0 _0433_
rlabel metal1 7222 12206 7222 12206 0 _0434_
rlabel metal1 10580 17646 10580 17646 0 _0435_
rlabel metal1 10810 17068 10810 17068 0 _0436_
rlabel metal1 10902 18088 10902 18088 0 _0437_
rlabel metal1 10718 18156 10718 18156 0 _0438_
rlabel metal1 7130 18870 7130 18870 0 _0439_
rlabel metal2 6854 19040 6854 19040 0 _0440_
rlabel metal2 11454 16966 11454 16966 0 _0441_
rlabel metal1 10580 17306 10580 17306 0 _0442_
rlabel metal1 11362 18394 11362 18394 0 _0443_
rlabel metal1 8878 13498 8878 13498 0 _0444_
rlabel metal2 12926 16354 12926 16354 0 _0445_
rlabel metal1 10948 16762 10948 16762 0 _0446_
rlabel metal1 11592 17646 11592 17646 0 _0447_
rlabel metal1 10396 17850 10396 17850 0 _0448_
rlabel metal2 10258 18156 10258 18156 0 _0449_
rlabel metal1 10074 17578 10074 17578 0 _0450_
rlabel metal1 10028 12818 10028 12818 0 _0451_
rlabel metal2 8510 20094 8510 20094 0 _0452_
rlabel metal2 8694 19618 8694 19618 0 _0453_
rlabel metal1 12972 18802 12972 18802 0 _0454_
rlabel metal1 10120 19482 10120 19482 0 _0455_
rlabel metal1 11638 20026 11638 20026 0 _0456_
rlabel metal1 12328 18734 12328 18734 0 _0457_
rlabel metal1 13616 18734 13616 18734 0 _0458_
rlabel metal1 13846 18802 13846 18802 0 _0459_
rlabel metal1 13018 16762 13018 16762 0 _0460_
rlabel metal2 12834 16932 12834 16932 0 _0461_
rlabel metal2 13018 16762 13018 16762 0 _0462_
rlabel metal1 13064 15470 13064 15470 0 _0463_
rlabel metal1 10350 15606 10350 15606 0 _0464_
rlabel metal2 10718 15742 10718 15742 0 _0465_
rlabel metal1 8326 15674 8326 15674 0 _0466_
rlabel metal1 8326 15436 8326 15436 0 _0467_
rlabel metal1 8602 16762 8602 16762 0 _0468_
rlabel metal2 8510 16388 8510 16388 0 _0469_
rlabel metal1 8410 16422 8410 16422 0 _0470_
rlabel metal1 7544 18054 7544 18054 0 _0471_
rlabel metal1 7774 17170 7774 17170 0 _0472_
rlabel metal2 4186 19873 4186 19873 0 _0473_
rlabel metal1 4600 21046 4600 21046 0 _0474_
rlabel metal2 3358 19822 3358 19822 0 _0475_
rlabel metal1 1978 19414 1978 19414 0 _0476_
rlabel metal1 7636 25262 7636 25262 0 _0477_
rlabel metal2 7774 22780 7774 22780 0 _0478_
rlabel metal1 7728 22202 7728 22202 0 _0479_
rlabel metal2 9522 24480 9522 24480 0 _0480_
rlabel metal1 8832 24378 8832 24378 0 _0481_
rlabel metal1 7682 27370 7682 27370 0 _0482_
rlabel metal1 7130 24786 7130 24786 0 _0483_
rlabel metal2 7314 25398 7314 25398 0 _0484_
rlabel metal1 7268 24854 7268 24854 0 _0485_
rlabel metal2 7130 26724 7130 26724 0 _0486_
rlabel metal1 7774 24922 7774 24922 0 _0487_
rlabel via1 7874 24106 7874 24106 0 _0488_
rlabel metal1 7774 25840 7774 25840 0 _0489_
rlabel metal2 8326 26180 8326 26180 0 _0490_
rlabel metal1 8648 24922 8648 24922 0 _0491_
rlabel metal2 8970 26180 8970 26180 0 _0492_
rlabel metal1 8188 24922 8188 24922 0 _0493_
rlabel metal2 9338 27200 9338 27200 0 _0494_
rlabel metal1 5060 13294 5060 13294 0 _0495_
rlabel metal1 5842 13260 5842 13260 0 _0496_
rlabel metal1 6624 12614 6624 12614 0 _0497_
rlabel metal1 6402 12954 6402 12954 0 _0498_
rlabel metal2 7498 12036 7498 12036 0 _0499_
rlabel metal1 8188 12070 8188 12070 0 _0500_
rlabel metal1 6026 13804 6026 13804 0 _0501_
rlabel metal1 4646 14960 4646 14960 0 _0502_
rlabel metal2 3450 11356 3450 11356 0 _0503_
rlabel metal2 3634 10948 3634 10948 0 _0504_
rlabel metal1 2622 10676 2622 10676 0 _0505_
rlabel metal1 2070 12308 2070 12308 0 _0506_
rlabel metal2 3174 10234 3174 10234 0 _0507_
rlabel metal1 5888 10438 5888 10438 0 _0508_
rlabel metal2 3450 9146 3450 9146 0 _0509_
rlabel metal1 2714 9588 2714 9588 0 _0510_
rlabel metal1 1932 8398 1932 8398 0 _0511_
rlabel metal1 1886 7344 1886 7344 0 _0512_
rlabel metal1 1702 7412 1702 7412 0 _0513_
rlabel metal1 2806 6732 2806 6732 0 _0514_
rlabel metal1 2622 6800 2622 6800 0 _0515_
rlabel metal2 3358 5916 3358 5916 0 _0516_
rlabel metal1 4094 5678 4094 5678 0 _0517_
rlabel metal2 3910 6052 3910 6052 0 _0518_
rlabel metal1 6824 6358 6824 6358 0 _0519_
rlabel via1 8610 7786 8610 7786 0 _0520_
rlabel metal1 8326 6834 8326 6834 0 _0521_
rlabel metal1 7774 6834 7774 6834 0 _0522_
rlabel metal2 8970 6052 8970 6052 0 _0523_
rlabel metal1 9292 7854 9292 7854 0 _0524_
rlabel metal1 9476 7854 9476 7854 0 _0525_
rlabel metal1 9614 8058 9614 8058 0 _0526_
rlabel metal2 13662 11696 13662 11696 0 _0527_
rlabel metal1 12650 11152 12650 11152 0 _0528_
rlabel metal2 12190 9316 12190 9316 0 _0529_
rlabel metal1 12558 8500 12558 8500 0 _0530_
rlabel metal2 10350 8262 10350 8262 0 _0531_
rlabel metal1 10488 8602 10488 8602 0 _0532_
rlabel metal2 12834 8738 12834 8738 0 _0533_
rlabel metal1 13110 7310 13110 7310 0 _0534_
rlabel metal1 12742 7344 12742 7344 0 _0535_
rlabel metal2 12834 7820 12834 7820 0 _0536_
rlabel metal1 10902 7922 10902 7922 0 _0537_
rlabel metal1 11408 7514 11408 7514 0 _0538_
rlabel metal2 8326 11322 8326 11322 0 _0539_
rlabel via1 13302 10982 13302 10982 0 _0540_
rlabel metal1 8418 11696 8418 11696 0 _0541_
rlabel metal2 13386 10438 13386 10438 0 _0542_
rlabel metal2 13754 11424 13754 11424 0 _0543_
rlabel metal2 13478 11526 13478 11526 0 _0544_
rlabel metal2 13938 11492 13938 11492 0 _0545_
rlabel metal1 12374 11220 12374 11220 0 _0546_
rlabel metal1 13432 12274 13432 12274 0 _0547_
rlabel metal1 12190 10098 12190 10098 0 _0548_
rlabel metal1 14398 12240 14398 12240 0 _0549_
rlabel metal1 12512 13974 12512 13974 0 _0550_
rlabel metal1 12926 13838 12926 13838 0 _0551_
rlabel metal1 12604 12818 12604 12818 0 _0552_
rlabel metal2 12190 14246 12190 14246 0 _0553_
rlabel metal2 12006 14212 12006 14212 0 _0554_
rlabel metal1 10856 13498 10856 13498 0 _0555_
rlabel metal1 11086 12818 11086 12818 0 _0556_
rlabel metal1 10718 12750 10718 12750 0 _0557_
rlabel metal1 20700 29614 20700 29614 0 _0558_
rlabel metal2 27646 28084 27646 28084 0 _0559_
rlabel metal1 18446 28186 18446 28186 0 _0560_
rlabel metal1 19918 29614 19918 29614 0 _0561_
rlabel metal1 19780 28186 19780 28186 0 _0562_
rlabel via1 26542 27435 26542 27435 0 _0563_
rlabel metal1 17848 27574 17848 27574 0 _0564_
rlabel metal1 18124 30634 18124 30634 0 _0565_
rlabel metal1 17664 29002 17664 29002 0 _0566_
rlabel metal1 17342 30362 17342 30362 0 _0567_
rlabel metal1 17342 30770 17342 30770 0 _0568_
rlabel metal1 20332 29206 20332 29206 0 _0569_
rlabel metal1 21206 29172 21206 29172 0 _0570_
rlabel metal1 18952 28730 18952 28730 0 _0571_
rlabel metal1 21068 29138 21068 29138 0 _0572_
rlabel metal1 19504 29750 19504 29750 0 _0573_
rlabel metal2 19734 30260 19734 30260 0 _0574_
rlabel metal1 20240 30566 20240 30566 0 _0575_
rlabel metal1 22494 28594 22494 28594 0 _0576_
rlabel metal1 22954 29104 22954 29104 0 _0577_
rlabel metal2 21850 28934 21850 28934 0 _0578_
rlabel metal2 21482 28696 21482 28696 0 _0579_
rlabel metal1 22034 28527 22034 28527 0 _0580_
rlabel metal2 21298 29478 21298 29478 0 _0581_
rlabel metal1 21390 30158 21390 30158 0 _0582_
rlabel metal1 24932 29070 24932 29070 0 _0583_
rlabel metal1 23000 28730 23000 28730 0 _0584_
rlabel metal1 23046 28492 23046 28492 0 _0585_
rlabel metal1 23598 29002 23598 29002 0 _0586_
rlabel metal1 23644 28934 23644 28934 0 _0587_
rlabel metal1 24426 29274 24426 29274 0 _0588_
rlabel metal1 24702 29580 24702 29580 0 _0589_
rlabel metal1 26542 29172 26542 29172 0 _0590_
rlabel metal2 26634 29444 26634 29444 0 _0591_
rlabel metal1 25668 29138 25668 29138 0 _0592_
rlabel metal1 24794 28084 24794 28084 0 _0593_
rlabel metal1 24886 28016 24886 28016 0 _0594_
rlabel metal1 26726 29818 26726 29818 0 _0595_
rlabel metal1 26496 29614 26496 29614 0 _0596_
rlabel metal1 26358 29818 26358 29818 0 _0597_
rlabel metal1 26818 28662 26818 28662 0 _0598_
rlabel metal2 27094 28730 27094 28730 0 _0599_
rlabel metal2 28842 27914 28842 27914 0 _0600_
rlabel metal1 28934 27472 28934 27472 0 _0601_
rlabel metal1 30774 29172 30774 29172 0 _0602_
rlabel metal2 30590 29308 30590 29308 0 _0603_
rlabel metal1 30176 29002 30176 29002 0 _0604_
rlabel metal1 30038 28730 30038 28730 0 _0605_
rlabel metal1 31326 28662 31326 28662 0 _0606_
rlabel metal1 30728 28186 30728 28186 0 _0607_
rlabel metal2 30314 27438 30314 27438 0 _0608_
rlabel metal2 23046 27200 23046 27200 0 _0609_
rlabel metal2 30406 26826 30406 26826 0 _0610_
rlabel metal2 32062 28900 32062 28900 0 _0611_
rlabel metal1 31602 28492 31602 28492 0 _0612_
rlabel metal2 32338 28220 32338 28220 0 _0613_
rlabel metal2 33534 27778 33534 27778 0 _0614_
rlabel metal1 35788 28458 35788 28458 0 _0615_
rlabel metal2 36202 28934 36202 28934 0 _0616_
rlabel metal1 36110 29172 36110 29172 0 _0617_
rlabel metal1 34638 29682 34638 29682 0 _0618_
rlabel metal1 35006 28730 35006 28730 0 _0619_
rlabel metal1 35742 27506 35742 27506 0 _0620_
rlabel metal2 36662 27200 36662 27200 0 _0621_
rlabel metal1 34408 28730 34408 28730 0 _0622_
rlabel metal1 34776 29818 34776 29818 0 _0623_
rlabel metal2 35098 30532 35098 30532 0 _0624_
rlabel metal1 35512 30362 35512 30362 0 _0625_
rlabel metal1 35006 27404 35006 27404 0 _0626_
rlabel metal1 34776 27506 34776 27506 0 _0627_
rlabel metal2 35282 27132 35282 27132 0 _0628_
rlabel metal2 34730 27642 34730 27642 0 _0629_
rlabel via2 18722 30107 18722 30107 0 _0630_
rlabel metal2 34178 29410 34178 29410 0 _0631_
rlabel metal2 33718 29988 33718 29988 0 _0632_
rlabel metal2 32982 30022 32982 30022 0 _0633_
rlabel metal1 22724 25262 22724 25262 0 _0634_
rlabel metal1 18722 24208 18722 24208 0 _0635_
rlabel metal2 18446 24837 18446 24837 0 _0636_
rlabel metal1 18630 23800 18630 23800 0 _0637_
rlabel metal1 20286 23630 20286 23630 0 _0638_
rlabel metal2 18814 23868 18814 23868 0 _0639_
rlabel metal2 17986 23052 17986 23052 0 _0640_
rlabel metal1 20286 24786 20286 24786 0 _0641_
rlabel metal1 20102 24718 20102 24718 0 _0642_
rlabel metal1 20332 23834 20332 23834 0 _0643_
rlabel metal1 19826 23834 19826 23834 0 _0644_
rlabel metal1 19642 23154 19642 23154 0 _0645_
rlabel metal2 21390 25398 21390 25398 0 _0646_
rlabel metal2 21482 26078 21482 26078 0 _0647_
rlabel metal1 21896 25942 21896 25942 0 _0648_
rlabel metal2 21666 25466 21666 25466 0 _0649_
rlabel metal1 21758 25296 21758 25296 0 _0650_
rlabel metal2 22310 24956 22310 24956 0 _0651_
rlabel metal1 23322 25942 23322 25942 0 _0652_
rlabel metal1 23690 26350 23690 26350 0 _0653_
rlabel via1 23874 26486 23874 26486 0 _0654_
rlabel metal2 23322 25500 23322 25500 0 _0655_
rlabel metal1 23230 25296 23230 25296 0 _0656_
rlabel metal1 23092 23834 23092 23834 0 _0657_
rlabel metal1 25300 24786 25300 24786 0 _0658_
rlabel metal1 25024 24650 25024 24650 0 _0659_
rlabel metal1 25208 24922 25208 24922 0 _0660_
rlabel metal1 25576 25262 25576 25262 0 _0661_
rlabel metal2 24978 25670 24978 25670 0 _0662_
rlabel metal1 26358 24106 26358 24106 0 _0663_
rlabel metal1 25898 24378 25898 24378 0 _0664_
rlabel metal1 25990 24174 25990 24174 0 _0665_
rlabel metal2 25162 24242 25162 24242 0 _0666_
rlabel metal2 29854 24446 29854 24446 0 _0667_
rlabel metal1 26818 24378 26818 24378 0 _0668_
rlabel metal2 27462 24990 27462 24990 0 _0669_
rlabel metal1 27508 23698 27508 23698 0 _0670_
rlabel metal1 29026 24820 29026 24820 0 _0671_
rlabel metal1 28934 24854 28934 24854 0 _0672_
rlabel metal1 28704 24922 28704 24922 0 _0673_
rlabel metal1 31510 24106 31510 24106 0 _0674_
rlabel metal1 30912 24378 30912 24378 0 _0675_
rlabel metal2 30498 24786 30498 24786 0 _0676_
rlabel metal1 30636 24174 30636 24174 0 _0677_
rlabel metal2 32982 24582 32982 24582 0 _0678_
rlabel metal2 33718 24718 33718 24718 0 _0679_
rlabel metal2 35374 24956 35374 24956 0 _0680_
rlabel metal1 35926 24820 35926 24820 0 _0681_
rlabel metal1 36386 24786 36386 24786 0 _0682_
rlabel metal1 35144 24174 35144 24174 0 _0683_
rlabel metal2 35650 24378 35650 24378 0 _0684_
rlabel metal1 35926 24038 35926 24038 0 _0685_
rlabel metal2 35282 22916 35282 22916 0 _0686_
rlabel via1 36570 23085 36570 23085 0 _0687_
rlabel metal1 36340 22746 36340 22746 0 _0688_
rlabel metal2 35742 23358 35742 23358 0 _0689_
rlabel metal1 35834 23052 35834 23052 0 _0690_
rlabel metal1 35374 22950 35374 22950 0 _0691_
rlabel metal2 17158 23681 17158 23681 0 _0692_
rlabel metal2 31510 23290 31510 23290 0 _0693_
rlabel metal1 31050 22950 31050 22950 0 _0694_
rlabel metal1 38042 11084 38042 11084 0 _0695_
rlabel metal1 14858 32980 14858 32980 0 _0696_
rlabel metal1 15686 34000 15686 34000 0 _0697_
rlabel metal2 15962 35938 15962 35938 0 _0698_
rlabel metal2 17158 19856 17158 19856 0 _0699_
rlabel metal1 18538 12954 18538 12954 0 _0700_
rlabel metal2 19090 15334 19090 15334 0 _0701_
rlabel metal1 19274 14382 19274 14382 0 _0702_
rlabel metal2 18814 15164 18814 15164 0 _0703_
rlabel metal1 18676 15674 18676 15674 0 _0704_
rlabel metal1 20148 15130 20148 15130 0 _0705_
rlabel metal1 19228 15674 19228 15674 0 _0706_
rlabel metal1 21804 16014 21804 16014 0 _0707_
rlabel metal2 21390 16456 21390 16456 0 _0708_
rlabel metal1 20746 16048 20746 16048 0 _0709_
rlabel metal1 20286 15674 20286 15674 0 _0710_
rlabel metal1 20654 15980 20654 15980 0 _0711_
rlabel metal1 21160 16218 21160 16218 0 _0712_
rlabel metal1 22678 15334 22678 15334 0 _0713_
rlabel via1 21865 15470 21865 15470 0 _0714_
rlabel metal2 21022 15164 21022 15164 0 _0715_
rlabel metal2 22218 15130 22218 15130 0 _0716_
rlabel metal2 21482 14552 21482 14552 0 _0717_
rlabel metal2 24794 16388 24794 16388 0 _0718_
rlabel metal2 25070 16252 25070 16252 0 _0719_
rlabel metal2 24242 16388 24242 16388 0 _0720_
rlabel metal2 20838 15912 20838 15912 0 _0721_
rlabel metal2 24150 16422 24150 16422 0 _0722_
rlabel metal1 23828 16762 23828 16762 0 _0723_
rlabel metal1 26496 15470 26496 15470 0 _0724_
rlabel metal1 27232 15470 27232 15470 0 _0725_
rlabel metal1 25530 15538 25530 15538 0 _0726_
rlabel metal2 26266 15113 26266 15113 0 _0727_
rlabel metal2 26450 15436 26450 15436 0 _0728_
rlabel metal1 25438 15062 25438 15062 0 _0729_
rlabel metal1 24702 15062 24702 15062 0 _0730_
rlabel via1 29302 15606 29302 15606 0 _0731_
rlabel metal2 28658 15028 28658 15028 0 _0732_
rlabel metal1 28750 14994 28750 14994 0 _0733_
rlabel metal1 27922 15606 27922 15606 0 _0734_
rlabel metal1 29302 15946 29302 15946 0 _0735_
rlabel metal1 29164 14858 29164 14858 0 _0736_
rlabel metal2 30222 17340 30222 17340 0 _0737_
rlabel metal1 32706 17204 32706 17204 0 _0738_
rlabel metal1 29440 16558 29440 16558 0 _0739_
rlabel metal1 29348 16490 29348 16490 0 _0740_
rlabel metal2 28198 16932 28198 16932 0 _0741_
rlabel metal1 28520 16762 28520 16762 0 _0742_
rlabel metal1 33258 17204 33258 17204 0 _0743_
rlabel metal2 33534 17306 33534 17306 0 _0744_
rlabel metal1 32752 16558 32752 16558 0 _0745_
rlabel metal2 31786 15980 31786 15980 0 _0746_
rlabel metal1 33028 16626 33028 16626 0 _0747_
rlabel metal2 32246 16286 32246 16286 0 _0748_
rlabel metal1 35328 17510 35328 17510 0 _0749_
rlabel metal1 34454 17272 34454 17272 0 _0750_
rlabel metal1 34270 17136 34270 17136 0 _0751_
rlabel metal2 34086 16762 34086 16762 0 _0752_
rlabel metal1 33994 16592 33994 16592 0 _0753_
rlabel metal1 42136 18326 42136 18326 0 _0754_
rlabel metal1 41814 18156 41814 18156 0 _0755_
rlabel metal2 41722 17544 41722 17544 0 _0756_
rlabel metal1 35236 16694 35236 16694 0 _0757_
rlabel metal2 37582 16490 37582 16490 0 _0758_
rlabel metal1 38088 17034 38088 17034 0 _0759_
rlabel metal2 40158 16932 40158 16932 0 _0760_
rlabel via1 40065 16082 40065 16082 0 _0761_
rlabel metal1 40618 16116 40618 16116 0 _0762_
rlabel metal2 40526 16252 40526 16252 0 _0763_
rlabel metal2 40250 16745 40250 16745 0 _0764_
rlabel metal1 39284 14382 39284 14382 0 _0765_
rlabel metal2 39606 15028 39606 15028 0 _0766_
rlabel metal2 39146 15946 39146 15946 0 _0767_
rlabel metal1 38686 14314 38686 14314 0 _0768_
rlabel viali 38226 14383 38226 14383 0 _0769_
rlabel metal1 39468 13294 39468 13294 0 _0770_
rlabel metal2 39422 13226 39422 13226 0 _0771_
rlabel metal1 39146 13838 39146 13838 0 _0772_
rlabel metal1 39928 13158 39928 13158 0 _0773_
rlabel metal1 39468 14042 39468 14042 0 _0774_
rlabel metal2 34362 14076 34362 14076 0 _0775_
rlabel metal1 38318 13498 38318 13498 0 _0776_
rlabel metal1 35006 14518 35006 14518 0 _0777_
rlabel metal1 17664 23630 17664 23630 0 _0778_
rlabel metal1 16238 23630 16238 23630 0 _0779_
rlabel metal2 16422 23868 16422 23868 0 _0780_
rlabel metal1 18676 38726 18676 38726 0 _0781_
rlabel metal1 30958 36312 30958 36312 0 _0782_
rlabel metal1 30669 36006 30669 36006 0 _0783_
rlabel metal2 31142 36550 31142 36550 0 _0784_
rlabel metal1 34316 36006 34316 36006 0 _0785_
rlabel metal1 34316 36142 34316 36142 0 _0786_
rlabel metal1 33902 36074 33902 36074 0 _0787_
rlabel metal1 35834 36278 35834 36278 0 _0788_
rlabel metal1 38456 36006 38456 36006 0 _0789_
rlabel metal1 39330 36176 39330 36176 0 _0790_
rlabel metal1 37398 36074 37398 36074 0 _0791_
rlabel metal2 39054 36550 39054 36550 0 _0792_
rlabel metal1 39882 36720 39882 36720 0 _0793_
rlabel metal1 39790 36788 39790 36788 0 _0794_
rlabel metal2 38594 37162 38594 37162 0 _0795_
rlabel metal1 38502 37706 38502 37706 0 _0796_
rlabel metal1 39744 38522 39744 38522 0 _0797_
rlabel metal2 39698 38862 39698 38862 0 _0798_
rlabel metal1 38962 38964 38962 38964 0 _0799_
rlabel metal1 38410 38386 38410 38386 0 _0800_
rlabel metal1 37628 41514 37628 41514 0 _0801_
rlabel metal1 37812 41514 37812 41514 0 _0802_
rlabel metal1 36892 40086 36892 40086 0 _0803_
rlabel metal1 36570 39984 36570 39984 0 _0804_
rlabel metal2 34086 42194 34086 42194 0 _0805_
rlabel metal1 34224 42602 34224 42602 0 _0806_
rlabel metal1 32982 41548 32982 41548 0 _0807_
rlabel metal2 33258 42058 33258 42058 0 _0808_
rlabel viali 31418 42197 31418 42197 0 _0809_
rlabel metal2 31878 41786 31878 41786 0 _0810_
rlabel metal1 32430 41650 32430 41650 0 _0811_
rlabel metal2 31142 40800 31142 40800 0 _0812_
rlabel metal1 28750 41480 28750 41480 0 _0813_
rlabel metal1 28106 41242 28106 41242 0 _0814_
rlabel via2 28106 40477 28106 40477 0 _0815_
rlabel metal2 28566 40834 28566 40834 0 _0816_
rlabel metal1 26450 41106 26450 41106 0 _0817_
rlabel metal1 26174 41038 26174 41038 0 _0818_
rlabel metal1 29118 40460 29118 40460 0 _0819_
rlabel metal2 26082 40766 26082 40766 0 _0820_
rlabel metal1 25300 38930 25300 38930 0 _0821_
rlabel metal1 24840 38930 24840 38930 0 _0822_
rlabel metal2 25254 39100 25254 39100 0 _0823_
rlabel via1 25346 39406 25346 39406 0 _0824_
rlabel metal1 23552 41242 23552 41242 0 _0825_
rlabel metal1 23414 40970 23414 40970 0 _0826_
rlabel metal2 24610 40256 24610 40256 0 _0827_
rlabel metal1 20838 40460 20838 40460 0 _0828_
rlabel metal2 21942 41786 21942 41786 0 _0829_
rlabel metal1 21390 43078 21390 43078 0 _0830_
rlabel metal1 21206 41072 21206 41072 0 _0831_
rlabel metal1 21482 41446 21482 41446 0 _0832_
rlabel metal2 18906 40732 18906 40732 0 _0833_
rlabel metal1 20562 40562 20562 40562 0 _0834_
rlabel metal2 18722 39236 18722 39236 0 _0835_
rlabel metal2 20378 40834 20378 40834 0 _0836_
rlabel metal2 20746 40188 20746 40188 0 _0837_
rlabel metal1 22034 40052 22034 40052 0 _0838_
rlabel metal1 24840 40018 24840 40018 0 _0839_
rlabel metal2 24794 39610 24794 39610 0 _0840_
rlabel metal1 25760 40018 25760 40018 0 _0841_
rlabel metal1 29210 40426 29210 40426 0 _0842_
rlabel metal1 28014 40052 28014 40052 0 _0843_
rlabel metal1 28612 40494 28612 40494 0 _0844_
rlabel metal1 33258 41650 33258 41650 0 _0845_
rlabel metal1 32338 41140 32338 41140 0 _0846_
rlabel metal2 32798 40970 32798 40970 0 _0847_
rlabel metal1 37444 39406 37444 39406 0 _0848_
rlabel metal2 37674 39100 37674 39100 0 _0849_
rlabel metal2 37858 38284 37858 38284 0 _0850_
rlabel metal1 37766 37230 37766 37230 0 _0851_
rlabel metal1 37122 36142 37122 36142 0 _0852_
rlabel metal2 37214 36448 37214 36448 0 _0853_
rlabel metal2 37490 36839 37490 36839 0 _0854_
rlabel metal2 31602 36924 31602 36924 0 _0855_
rlabel metal2 30682 36992 30682 36992 0 _0856_
rlabel metal1 30866 36788 30866 36788 0 _0857_
rlabel metal1 36478 38998 36478 38998 0 _0858_
rlabel metal2 18814 39644 18814 39644 0 _0859_
rlabel via1 19734 38930 19734 38930 0 _0860_
rlabel metal1 20102 38318 20102 38318 0 _0861_
rlabel metal1 19872 38386 19872 38386 0 _0862_
rlabel metal1 20010 38454 20010 38454 0 _0863_
rlabel metal1 21206 38930 21206 38930 0 _0864_
rlabel metal2 20838 40460 20838 40460 0 _0865_
rlabel metal1 21206 38998 21206 38998 0 _0866_
rlabel metal2 21298 38148 21298 38148 0 _0867_
rlabel metal2 21206 38012 21206 38012 0 _0868_
rlabel metal2 21850 39134 21850 39134 0 _0869_
rlabel metal2 22586 40154 22586 40154 0 _0870_
rlabel metal1 22402 39406 22402 39406 0 _0871_
rlabel metal1 22678 38318 22678 38318 0 _0872_
rlabel metal2 22678 38828 22678 38828 0 _0873_
rlabel metal2 24426 39236 24426 39236 0 _0874_
rlabel metal1 25254 38284 25254 38284 0 _0875_
rlabel metal1 25254 39474 25254 39474 0 _0876_
rlabel metal2 25622 39134 25622 39134 0 _0877_
rlabel metal1 25806 36890 25806 36890 0 _0878_
rlabel metal2 26726 38522 26726 38522 0 _0879_
rlabel metal2 26082 40154 26082 40154 0 _0880_
rlabel metal2 27002 39134 27002 39134 0 _0881_
rlabel metal2 27278 38148 27278 38148 0 _0882_
rlabel metal2 27186 38012 27186 38012 0 _0883_
rlabel metal2 28290 38148 28290 38148 0 _0884_
rlabel metal2 27922 40154 27922 40154 0 _0885_
rlabel metal2 28382 39406 28382 39406 0 _0886_
rlabel metal2 28474 36992 28474 36992 0 _0887_
rlabel metal1 28612 38318 28612 38318 0 _0888_
rlabel metal1 28474 40596 28474 40596 0 _0889_
rlabel metal1 28704 38998 28704 38998 0 _0890_
rlabel metal2 29578 38080 29578 38080 0 _0891_
rlabel metal1 32154 39338 32154 39338 0 _0892_
rlabel metal1 30774 38964 30774 38964 0 _0893_
rlabel metal2 33074 40834 33074 40834 0 _0894_
rlabel metal1 32752 39610 32752 39610 0 _0895_
rlabel metal1 25024 37162 25024 37162 0 _0896_
rlabel metal1 32108 39610 32108 39610 0 _0897_
rlabel metal1 34684 40154 34684 40154 0 _0898_
rlabel metal2 32430 40222 32430 40222 0 _0899_
rlabel metal2 32430 39066 32430 39066 0 _0900_
rlabel metal1 32292 38386 32292 38386 0 _0901_
rlabel metal2 34362 38760 34362 38760 0 _0902_
rlabel metal1 36202 38896 36202 38896 0 _0903_
rlabel metal1 38180 38862 38180 38862 0 _0904_
rlabel metal1 35374 38862 35374 38862 0 _0905_
rlabel metal1 36064 37842 36064 37842 0 _0906_
rlabel metal1 34224 38522 34224 38522 0 _0907_
rlabel metal1 38042 37774 38042 37774 0 _0908_
rlabel metal2 35098 38012 35098 38012 0 _0909_
rlabel metal1 35006 39440 35006 39440 0 _0910_
rlabel metal1 35052 38522 35052 38522 0 _0911_
rlabel metal1 35098 37196 35098 37196 0 _0912_
rlabel metal2 36386 36924 36386 36924 0 _0913_
rlabel metal1 37260 36210 37260 36210 0 _0914_
rlabel metal2 36478 36516 36478 36516 0 _0915_
rlabel metal2 36018 35870 36018 35870 0 _0916_
rlabel metal1 36018 35666 36018 35666 0 _0917_
rlabel metal1 34638 36346 34638 36346 0 _0918_
rlabel metal1 35512 36618 35512 36618 0 _0919_
rlabel metal1 35098 35700 35098 35700 0 _0920_
rlabel metal2 35190 35615 35190 35615 0 _0921_
rlabel metal1 35190 36890 35190 36890 0 _0922_
rlabel metal1 31418 36686 31418 36686 0 _0923_
rlabel metal1 32016 36890 32016 36890 0 _0924_
rlabel metal1 32614 36210 32614 36210 0 _0925_
rlabel metal1 19550 36788 19550 36788 0 _0926_
rlabel metal1 16652 34102 16652 34102 0 _0927_
rlabel metal1 17112 37434 17112 37434 0 _0928_
rlabel metal1 17342 40154 17342 40154 0 _0929_
rlabel metal1 19964 42670 19964 42670 0 _0930_
rlabel metal1 22816 35802 22816 35802 0 _0931_
rlabel metal2 24886 36006 24886 36006 0 _0932_
rlabel metal1 25806 42534 25806 42534 0 _0933_
rlabel metal1 27968 33626 27968 33626 0 _0934_
rlabel metal1 30084 39610 30084 39610 0 _0935_
rlabel metal1 33994 41242 33994 41242 0 _0936_
rlabel metal2 39330 40596 39330 40596 0 _0937_
rlabel metal1 41262 37978 41262 37978 0 _0938_
rlabel metal1 40802 34170 40802 34170 0 _0939_
rlabel metal1 38916 33626 38916 33626 0 _0940_
rlabel metal1 34408 33626 34408 33626 0 _0941_
rlabel metal2 30222 34850 30222 34850 0 _0942_
rlabel metal2 16238 37638 16238 37638 0 _0943_
rlabel metal2 17802 40868 17802 40868 0 _0944_
rlabel metal1 20516 42534 20516 42534 0 _0945_
rlabel metal1 23046 41514 23046 41514 0 _0946_
rlabel metal1 25530 34714 25530 34714 0 _0947_
rlabel metal1 26910 33626 26910 33626 0 _0948_
rlabel metal1 27830 34170 27830 34170 0 _0949_
rlabel metal1 30728 39610 30728 39610 0 _0950_
rlabel metal2 35190 41344 35190 41344 0 _0951_
rlabel metal1 38088 40970 38088 40970 0 _0952_
rlabel metal2 40342 38624 40342 38624 0 _0953_
rlabel metal1 41032 34714 41032 34714 0 _0954_
rlabel metal1 38042 33626 38042 33626 0 _0955_
rlabel metal1 33442 33626 33442 33626 0 _0956_
rlabel metal1 30958 33626 30958 33626 0 _0957_
rlabel metal2 14674 34544 14674 34544 0 _0958_
rlabel via4 38732 27608 38732 27608 0 _0959_
rlabel metal1 14904 24378 14904 24378 0 _0960_
rlabel metal1 15640 22066 15640 22066 0 _0961_
rlabel metal1 13478 22542 13478 22542 0 _0962_
rlabel metal2 15226 30090 15226 30090 0 _0963_
rlabel metal2 16238 26044 16238 26044 0 _0964_
rlabel metal1 20148 20026 20148 20026 0 _0965_
rlabel metal1 17158 21590 17158 21590 0 _0966_
rlabel metal1 16698 21590 16698 21590 0 _0967_
rlabel via2 17158 16099 17158 16099 0 _0968_
rlabel metal1 18446 18394 18446 18394 0 _0969_
rlabel metal1 22494 21658 22494 21658 0 _0970_
rlabel viali 23886 31790 23886 31790 0 _0971_
rlabel metal2 40894 24735 40894 24735 0 _0972_
rlabel metal2 38502 28271 38502 28271 0 _0973_
rlabel metal1 39054 23086 39054 23086 0 _0974_
rlabel via2 39330 27421 39330 27421 0 _0975_
rlabel metal1 32936 19890 32936 19890 0 _0976_
rlabel metal1 39054 26758 39054 26758 0 _0977_
rlabel metal1 40664 20502 40664 20502 0 _0978_
rlabel metal1 41492 23698 41492 23698 0 _0979_
rlabel metal1 38456 22746 38456 22746 0 _0980_
rlabel metal2 40066 26214 40066 26214 0 _0981_
rlabel metal1 31418 15538 31418 15538 0 _0982_
rlabel via2 16054 20995 16054 20995 0 _0983_
rlabel metal2 21574 33796 21574 33796 0 _0984_
rlabel metal1 13846 23154 13846 23154 0 _0985_
rlabel metal1 12466 22542 12466 22542 0 _0986_
rlabel metal1 13570 24174 13570 24174 0 _0987_
rlabel metal2 15134 25534 15134 25534 0 _0988_
rlabel metal2 14950 24956 14950 24956 0 _0989_
rlabel metal1 14674 24820 14674 24820 0 _0990_
rlabel metal2 14214 23868 14214 23868 0 _0991_
rlabel metal1 17296 29002 17296 29002 0 _0992_
rlabel metal1 17480 29750 17480 29750 0 _0993_
rlabel metal1 18078 29138 18078 29138 0 _0994_
rlabel metal1 17158 27098 17158 27098 0 _0995_
rlabel metal1 19228 29818 19228 29818 0 _0996_
rlabel metal1 29210 26860 29210 26860 0 _0997_
rlabel metal2 22034 27710 22034 27710 0 _0998_
rlabel metal1 20010 33490 20010 33490 0 _0999_
rlabel metal1 21022 32470 21022 32470 0 _1000_
rlabel metal1 21022 32368 21022 32368 0 _1001_
rlabel metal2 22126 31314 22126 31314 0 _1002_
rlabel metal1 21988 31790 21988 31790 0 _1003_
rlabel metal1 24242 30906 24242 30906 0 _1004_
rlabel metal2 24058 32232 24058 32232 0 _1005_
rlabel metal1 40710 25160 40710 25160 0 _1006_
rlabel metal1 40618 24922 40618 24922 0 _1007_
rlabel metal2 37674 28577 37674 28577 0 _1008_
rlabel metal1 38088 28186 38088 28186 0 _1009_
rlabel via2 39514 24123 39514 24123 0 _1010_
rlabel metal1 39238 23290 39238 23290 0 _1011_
rlabel metal1 40434 27982 40434 27982 0 _1012_
rlabel metal1 39606 27574 39606 27574 0 _1013_
rlabel metal1 37490 26316 37490 26316 0 _1014_
rlabel metal1 37398 26384 37398 26384 0 _1015_
rlabel metal2 34178 26707 34178 26707 0 _1016_
rlabel metal1 40572 26010 40572 26010 0 _1017_
rlabel metal1 37076 30226 37076 30226 0 _1018_
rlabel metal1 40112 29614 40112 29614 0 _1019_
rlabel metal1 40158 22984 40158 22984 0 _1020_
rlabel metal1 40342 22984 40342 22984 0 _1021_
rlabel metal1 36570 29614 36570 29614 0 _1022_
rlabel metal1 38732 29750 38732 29750 0 _1023_
rlabel metal2 39330 26214 39330 26214 0 _1024_
rlabel metal1 39514 25976 39514 25976 0 _1025_
rlabel metal1 32016 29138 32016 29138 0 _1026_
rlabel metal1 32890 28934 32890 28934 0 _1027_
rlabel metal1 18676 29274 18676 29274 0 _1028_
rlabel metal1 35236 24786 35236 24786 0 _1029_
rlabel metal1 30544 23834 30544 23834 0 _1030_
rlabel metal1 13524 25126 13524 25126 0 _1031_
rlabel metal1 7084 29138 7084 29138 0 _1032_
rlabel metal1 5934 16218 5934 16218 0 _1033_
rlabel via2 28106 12835 28106 12835 0 _1034_
rlabel metal2 17986 26112 17986 26112 0 _1035_
rlabel metal1 17756 26350 17756 26350 0 _1036_
rlabel metal1 20838 26384 20838 26384 0 _1037_
rlabel metal1 17526 16116 17526 16116 0 _1038_
rlabel metal1 35144 11118 35144 11118 0 _1039_
rlabel metal1 19642 12886 19642 12886 0 _1040_
rlabel metal2 20838 38046 20838 38046 0 _1041_
rlabel metal2 8970 24004 8970 24004 0 _1042_
rlabel metal2 9062 21726 9062 21726 0 _1043_
rlabel metal2 9062 11084 9062 11084 0 _1044_
rlabel metal1 29854 36584 29854 36584 0 _1045_
rlabel metal1 4600 28526 4600 28526 0 _1046_
rlabel metal2 5842 30464 5842 30464 0 _1047_
rlabel metal1 6210 33932 6210 33932 0 _1048_
rlabel metal1 5888 34170 5888 34170 0 _1049_
rlabel metal1 5704 30838 5704 30838 0 _1050_
rlabel metal2 6578 30396 6578 30396 0 _1051_
rlabel metal1 6072 28730 6072 28730 0 _1052_
rlabel metal1 4140 27438 4140 27438 0 _1053_
rlabel metal2 4646 27982 4646 27982 0 _1054_
rlabel metal1 6808 20230 6808 20230 0 _1055_
rlabel via1 5103 26350 5103 26350 0 _1056_
rlabel metal1 5382 25806 5382 25806 0 _1057_
rlabel metal2 4002 24208 4002 24208 0 _1058_
rlabel metal1 6164 20026 6164 20026 0 _1059_
rlabel metal1 6624 23698 6624 23698 0 _1060_
rlabel metal2 4554 25024 4554 25024 0 _1061_
rlabel metal1 4922 26928 4922 26928 0 _1062_
rlabel metal1 4370 26996 4370 26996 0 _1063_
rlabel metal1 4646 26928 4646 26928 0 _1064_
rlabel metal1 5290 29614 5290 29614 0 _1065_
rlabel metal1 4830 24752 4830 24752 0 _1066_
rlabel metal2 2530 24174 2530 24174 0 _1067_
rlabel metal2 39192 12750 39192 12750 0 _1068_
rlabel metal1 26542 11628 26542 11628 0 _1069_
rlabel metal1 24058 11594 24058 11594 0 _1070_
rlabel metal1 33626 12138 33626 12138 0 _1071_
rlabel metal2 27002 12070 27002 12070 0 _1072_
rlabel metal1 27968 12682 27968 12682 0 _1073_
rlabel metal2 21666 9180 21666 9180 0 _1074_
rlabel metal2 24518 8126 24518 8126 0 _1075_
rlabel metal1 27278 7922 27278 7922 0 _1076_
rlabel metal1 28244 7378 28244 7378 0 _1077_
rlabel metal1 29992 7446 29992 7446 0 _1078_
rlabel metal1 33902 7446 33902 7446 0 _1079_
rlabel metal1 35650 7310 35650 7310 0 _1080_
rlabel metal1 36662 8466 36662 8466 0 _1081_
rlabel metal2 38594 9367 38594 9367 0 _1082_
rlabel metal1 38134 9520 38134 9520 0 _1083_
rlabel metal2 37674 9860 37674 9860 0 _1084_
rlabel metal1 35512 7378 35512 7378 0 _1085_
rlabel metal1 35604 9554 35604 9554 0 _1086_
rlabel metal1 35466 9656 35466 9656 0 _1087_
rlabel metal1 23092 8602 23092 8602 0 _1088_
rlabel metal1 21666 9520 21666 9520 0 _1089_
rlabel metal1 22034 11084 22034 11084 0 _1090_
rlabel metal1 22494 9078 22494 9078 0 _1091_
rlabel metal1 20056 9554 20056 9554 0 _1092_
rlabel metal2 19550 9248 19550 9248 0 _1093_
rlabel metal1 20746 9486 20746 9486 0 _1094_
rlabel metal2 22310 9724 22310 9724 0 _1095_
rlabel metal1 23598 9996 23598 9996 0 _1096_
rlabel metal2 24978 7174 24978 7174 0 _1097_
rlabel metal1 24610 10030 24610 10030 0 _1098_
rlabel metal2 27002 8262 27002 8262 0 _1099_
rlabel metal2 27186 9078 27186 9078 0 _1100_
rlabel metal1 28382 10132 28382 10132 0 _1101_
rlabel metal2 28198 7582 28198 7582 0 _1102_
rlabel metal2 27370 9758 27370 9758 0 _1103_
rlabel metal1 27646 9418 27646 9418 0 _1104_
rlabel metal1 29578 9962 29578 9962 0 _1105_
rlabel via1 28106 10031 28106 10031 0 _1106_
rlabel metal1 30866 10030 30866 10030 0 _1107_
rlabel metal2 29854 8500 29854 8500 0 _1108_
rlabel metal1 30958 10166 30958 10166 0 _1109_
rlabel metal1 32246 7344 32246 7344 0 _1110_
rlabel metal2 32706 9792 32706 9792 0 _1111_
rlabel metal2 31234 9894 31234 9894 0 _1112_
rlabel metal2 32614 9350 32614 9350 0 _1113_
rlabel metal2 32246 9622 32246 9622 0 _1114_
rlabel metal1 32735 8942 32735 8942 0 _1115_
rlabel metal1 33580 9146 33580 9146 0 _1116_
rlabel metal2 36018 7854 36018 7854 0 _1117_
rlabel metal1 36202 7174 36202 7174 0 _1118_
rlabel metal1 35696 10234 35696 10234 0 _1119_
rlabel metal1 35144 10710 35144 10710 0 _1120_
rlabel metal1 37582 8602 37582 8602 0 _1121_
rlabel metal1 36294 8976 36294 8976 0 _1122_
rlabel metal1 36018 10676 36018 10676 0 _1123_
rlabel viali 35925 10642 35925 10642 0 _1124_
rlabel metal1 35328 10778 35328 10778 0 _1125_
rlabel metal2 35558 11424 35558 11424 0 _1126_
rlabel metal1 22126 12376 22126 12376 0 _1127_
rlabel metal1 6440 29682 6440 29682 0 _1128_
rlabel metal1 6670 28730 6670 28730 0 _1129_
rlabel metal2 5934 29852 5934 29852 0 _1130_
rlabel metal1 5336 28186 5336 28186 0 _1131_
rlabel metal2 5244 32300 5244 32300 0 _1132_
rlabel metal1 5934 31790 5934 31790 0 _1133_
rlabel metal2 5566 29716 5566 29716 0 _1134_
rlabel metal1 7682 31280 7682 31280 0 _1135_
rlabel metal1 7590 31246 7590 31246 0 _1136_
rlabel metal1 8924 30294 8924 30294 0 _1137_
rlabel metal1 9338 29818 9338 29818 0 _1138_
rlabel metal1 10028 32402 10028 32402 0 _1139_
rlabel metal2 9614 31790 9614 31790 0 _1140_
rlabel metal2 9522 31195 9522 31195 0 _1141_
rlabel metal1 9798 32946 9798 32946 0 _1142_
rlabel metal1 9706 32810 9706 32810 0 _1143_
rlabel metal2 9154 34000 9154 34000 0 _1144_
rlabel metal2 11086 33660 11086 33660 0 _1145_
rlabel metal1 10258 33932 10258 33932 0 _1146_
rlabel metal1 7636 34986 7636 34986 0 _1147_
rlabel metal1 8326 32878 8326 32878 0 _1148_
rlabel metal1 8878 35598 8878 35598 0 _1149_
rlabel metal1 7268 35258 7268 35258 0 _1150_
rlabel metal1 6854 36176 6854 36176 0 _1151_
rlabel metal1 9660 35054 9660 35054 0 _1152_
rlabel metal1 9614 35258 9614 35258 0 _1153_
rlabel metal2 5566 35904 5566 35904 0 _1154_
rlabel metal1 5474 36142 5474 36142 0 _1155_
rlabel metal1 2346 33592 2346 33592 0 _1156_
rlabel metal2 5382 35836 5382 35836 0 _1157_
rlabel metal1 4048 35258 4048 35258 0 _1158_
rlabel metal1 4508 36142 4508 36142 0 _1159_
rlabel metal1 3910 34612 3910 34612 0 _1160_
rlabel metal1 3772 34714 3772 34714 0 _1161_
rlabel metal2 3358 35258 3358 35258 0 _1162_
rlabel metal1 5382 32742 5382 32742 0 _1163_
rlabel metal1 4324 32946 4324 32946 0 _1164_
rlabel metal1 4048 32878 4048 32878 0 _1165_
rlabel metal1 5658 32504 5658 32504 0 _1166_
rlabel metal2 5658 32436 5658 32436 0 _1167_
rlabel metal2 5474 32606 5474 32606 0 _1168_
rlabel metal1 4830 29138 4830 29138 0 _1169_
rlabel metal2 4784 31348 4784 31348 0 _1170_
rlabel metal1 4186 32198 4186 32198 0 _1171_
rlabel metal1 4094 30634 4094 30634 0 _1172_
rlabel metal1 4784 29274 4784 29274 0 _1173_
rlabel metal1 4784 28730 4784 28730 0 _1174_
rlabel metal1 5520 29818 5520 29818 0 _1175_
rlabel metal2 5474 30566 5474 30566 0 _1176_
rlabel metal2 2438 32878 2438 32878 0 _1177_
rlabel metal2 2254 32844 2254 32844 0 _1178_
rlabel metal2 2438 30498 2438 30498 0 _1179_
rlabel metal2 1794 29376 1794 29376 0 _1180_
rlabel metal1 2346 30600 2346 30600 0 _1181_
rlabel metal1 2254 30736 2254 30736 0 _1182_
rlabel metal2 2438 29342 2438 29342 0 _1183_
rlabel metal1 2346 29104 2346 29104 0 _1184_
rlabel metal1 2254 29206 2254 29206 0 _1185_
rlabel metal1 3772 28662 3772 28662 0 _1186_
rlabel metal1 4922 21488 4922 21488 0 _1187_
rlabel metal1 6210 20842 6210 20842 0 _1188_
rlabel metal2 5658 23698 5658 23698 0 _1189_
rlabel metal1 5382 24242 5382 24242 0 _1190_
rlabel metal1 6348 20570 6348 20570 0 _1191_
rlabel metal2 6210 21114 6210 21114 0 _1192_
rlabel metal1 5842 17068 5842 17068 0 _1193_
rlabel metal2 5658 16932 5658 16932 0 _1194_
rlabel metal1 5244 17306 5244 17306 0 _1195_
rlabel metal1 5428 21114 5428 21114 0 _1196_
rlabel metal1 6072 17306 6072 17306 0 _1197_
rlabel via2 4922 17187 4922 17187 0 _1198_
rlabel metal2 5474 16796 5474 16796 0 _1199_
rlabel metal1 5566 16660 5566 16660 0 _1200_
rlabel metal2 5290 16898 5290 16898 0 _1201_
rlabel metal1 5980 16626 5980 16626 0 _1202_
rlabel metal1 5796 17850 5796 17850 0 _1203_
rlabel metal1 7498 23732 7498 23732 0 _1204_
rlabel metal1 8602 24820 8602 24820 0 _1205_
rlabel metal2 7314 21726 7314 21726 0 _1206_
rlabel metal1 17388 25738 17388 25738 0 _1207_
rlabel metal2 14858 28118 14858 28118 0 _1208_
rlabel metal2 14674 28050 14674 28050 0 _1209_
rlabel metal1 21206 26384 21206 26384 0 _1210_
rlabel metal1 33258 24650 33258 24650 0 _1211_
rlabel metal2 17618 24956 17618 24956 0 _1212_
rlabel metal2 15686 25568 15686 25568 0 _1213_
rlabel metal2 18538 26826 18538 26826 0 _1214_
rlabel metal1 18216 26962 18216 26962 0 _1215_
rlabel metal3 575 41956 575 41956 0 clk
rlabel metal1 15778 13430 15778 13430 0 clknet_0_clk
rlabel metal1 16652 14994 16652 14994 0 clknet_2_0__leaf_clk
rlabel metal1 14628 37162 14628 37162 0 clknet_2_1__leaf_clk
rlabel metal1 38180 16558 38180 16558 0 clknet_2_2__leaf_clk
rlabel metal1 33902 34680 33902 34680 0 clknet_2_3__leaf_clk
rlabel metal2 1518 11424 1518 11424 0 clknet_leaf_0_clk
rlabel metal1 2714 35700 2714 35700 0 clknet_leaf_10_clk
rlabel metal2 14766 39712 14766 39712 0 clknet_leaf_11_clk
rlabel metal2 19458 42398 19458 42398 0 clknet_leaf_12_clk
rlabel metal1 14766 36142 14766 36142 0 clknet_leaf_13_clk
rlabel metal1 20286 32946 20286 32946 0 clknet_leaf_14_clk
rlabel metal1 24564 27506 24564 27506 0 clknet_leaf_15_clk
rlabel metal2 29762 33728 29762 33728 0 clknet_leaf_16_clk
rlabel metal1 24288 40018 24288 40018 0 clknet_leaf_17_clk
rlabel metal2 29118 38964 29118 38964 0 clknet_leaf_18_clk
rlabel metal2 33994 38998 33994 38998 0 clknet_leaf_19_clk
rlabel metal2 2714 14688 2714 14688 0 clknet_leaf_1_clk
rlabel metal1 39376 41650 39376 41650 0 clknet_leaf_20_clk
rlabel metal2 39606 35904 39606 35904 0 clknet_leaf_21_clk
rlabel metal1 37306 32266 37306 32266 0 clknet_leaf_22_clk
rlabel metal1 39514 23766 39514 23766 0 clknet_leaf_23_clk
rlabel metal1 32200 31790 32200 31790 0 clknet_leaf_24_clk
rlabel metal2 28474 21250 28474 21250 0 clknet_leaf_25_clk
rlabel metal2 31970 15538 31970 15538 0 clknet_leaf_26_clk
rlabel metal1 40158 21998 40158 21998 0 clknet_leaf_27_clk
rlabel metal2 35282 17017 35282 17017 0 clknet_leaf_28_clk
rlabel metal1 35512 13362 35512 13362 0 clknet_leaf_29_clk
rlabel metal1 2208 16014 2208 16014 0 clknet_leaf_2_clk
rlabel metal1 38410 7888 38410 7888 0 clknet_leaf_30_clk
rlabel metal1 33350 9486 33350 9486 0 clknet_leaf_31_clk
rlabel metal2 28750 5984 28750 5984 0 clknet_leaf_32_clk
rlabel metal2 27922 12818 27922 12818 0 clknet_leaf_33_clk
rlabel metal1 24334 14450 24334 14450 0 clknet_leaf_34_clk
rlabel metal1 17710 19380 17710 19380 0 clknet_leaf_35_clk
rlabel metal1 16146 11186 16146 11186 0 clknet_leaf_36_clk
rlabel metal1 19918 6834 19918 6834 0 clknet_leaf_37_clk
rlabel metal1 11730 13294 11730 13294 0 clknet_leaf_38_clk
rlabel metal1 1610 5746 1610 5746 0 clknet_leaf_39_clk
rlabel metal1 9660 22066 9660 22066 0 clknet_leaf_3_clk
rlabel metal2 14398 16218 14398 16218 0 clknet_leaf_4_clk
rlabel metal2 18906 21760 18906 21760 0 clknet_leaf_5_clk
rlabel metal1 14858 30294 14858 30294 0 clknet_leaf_6_clk
rlabel metal2 9982 23936 9982 23936 0 clknet_leaf_7_clk
rlabel metal2 2714 31416 2714 31416 0 clknet_leaf_8_clk
rlabel metal1 4922 33524 4922 33524 0 clknet_leaf_9_clk
rlabel metal3 751 25908 751 25908 0 complete
rlabel metal1 20700 43418 20700 43418 0 display_output[0]
rlabel via2 41998 30005 41998 30005 0 display_output[10]
rlabel metal2 42182 22831 42182 22831 0 display_output[11]
rlabel metal3 42512 29308 42512 29308 0 display_output[12]
rlabel metal2 41538 25177 41538 25177 0 display_output[13]
rlabel metal2 42090 28815 42090 28815 0 display_output[14]
rlabel metal2 20286 44251 20286 44251 0 display_output[15]
rlabel metal2 21574 44251 21574 44251 0 display_output[1]
rlabel metal2 22770 44251 22770 44251 0 display_output[2]
rlabel metal2 24058 44251 24058 44251 0 display_output[3]
rlabel via2 41538 24565 41538 24565 0 display_output[4]
rlabel via2 41722 27931 41722 27931 0 display_output[5]
rlabel metal2 40250 23953 40250 23953 0 display_output[6]
rlabel metal2 42090 27557 42090 27557 0 display_output[7]
rlabel metal2 42090 25959 42090 25959 0 display_output[8]
rlabel metal2 42090 26673 42090 26673 0 display_output[9]
rlabel metal2 14398 25534 14398 25534 0 equal_input
rlabel metal1 14628 34510 14628 34510 0 gencon_inst.ALU_finish
rlabel metal1 16238 37162 16238 37162 0 gencon_inst.ALU_in1\[0\]
rlabel metal2 41170 37315 41170 37315 0 gencon_inst.ALU_in1\[10\]
rlabel metal2 41354 34884 41354 34884 0 gencon_inst.ALU_in1\[11\]
rlabel metal1 38778 33490 38778 33490 0 gencon_inst.ALU_in1\[12\]
rlabel metal1 34362 33490 34362 33490 0 gencon_inst.ALU_in1\[13\]
rlabel metal2 31602 33762 31602 33762 0 gencon_inst.ALU_in1\[14\]
rlabel metal2 15870 34442 15870 34442 0 gencon_inst.ALU_in1\[15\]
rlabel metal1 18078 40154 18078 40154 0 gencon_inst.ALU_in1\[1\]
rlabel metal2 21390 34204 21390 34204 0 gencon_inst.ALU_in1\[2\]
rlabel metal1 24840 35802 24840 35802 0 gencon_inst.ALU_in1\[3\]
rlabel metal1 25714 34646 25714 34646 0 gencon_inst.ALU_in1\[4\]
rlabel metal1 26864 33558 26864 33558 0 gencon_inst.ALU_in1\[5\]
rlabel metal1 28566 32980 28566 32980 0 gencon_inst.ALU_in1\[6\]
rlabel metal1 31142 39338 31142 39338 0 gencon_inst.ALU_in1\[7\]
rlabel metal1 35190 41174 35190 41174 0 gencon_inst.ALU_in1\[8\]
rlabel metal1 39284 40086 39284 40086 0 gencon_inst.ALU_in1\[9\]
rlabel metal2 16054 34884 16054 34884 0 gencon_inst.ALU_in2\[0\]
rlabel metal1 41722 32470 41722 32470 0 gencon_inst.ALU_in2\[10\]
rlabel metal2 41262 35156 41262 35156 0 gencon_inst.ALU_in2\[11\]
rlabel metal1 38410 33082 38410 33082 0 gencon_inst.ALU_in2\[12\]
rlabel metal2 34454 32096 34454 32096 0 gencon_inst.ALU_in2\[13\]
rlabel metal2 31510 33728 31510 33728 0 gencon_inst.ALU_in2\[14\]
rlabel metal2 15502 32402 15502 32402 0 gencon_inst.ALU_in2\[15\]
rlabel metal1 19826 35020 19826 35020 0 gencon_inst.ALU_in2\[1\]
rlabel metal2 20930 35360 20930 35360 0 gencon_inst.ALU_in2\[2\]
rlabel metal1 22724 33830 22724 33830 0 gencon_inst.ALU_in2\[3\]
rlabel metal1 25484 33830 25484 33830 0 gencon_inst.ALU_in2\[4\]
rlabel metal1 26542 33490 26542 33490 0 gencon_inst.ALU_in2\[5\]
rlabel metal1 28566 33490 28566 33490 0 gencon_inst.ALU_in2\[6\]
rlabel metal2 30682 32538 30682 32538 0 gencon_inst.ALU_in2\[7\]
rlabel metal1 34822 41072 34822 41072 0 gencon_inst.ALU_in2\[8\]
rlabel metal1 39698 40154 39698 40154 0 gencon_inst.ALU_in2\[9\]
rlabel metal1 18630 30736 18630 30736 0 gencon_inst.ALU_out\[0\]
rlabel metal2 37766 37553 37766 37553 0 gencon_inst.ALU_out\[10\]
rlabel via2 35742 38811 35742 38811 0 gencon_inst.ALU_out\[11\]
rlabel metal1 36846 33422 36846 33422 0 gencon_inst.ALU_out\[12\]
rlabel metal1 36800 34442 36800 34442 0 gencon_inst.ALU_out\[13\]
rlabel viali 33259 29614 33259 29614 0 gencon_inst.ALU_out\[14\]
rlabel metal1 18814 36006 18814 36006 0 gencon_inst.ALU_out\[15\]
rlabel metal2 20562 36737 20562 36737 0 gencon_inst.ALU_out\[1\]
rlabel metal1 22724 37434 22724 37434 0 gencon_inst.ALU_out\[2\]
rlabel metal1 24058 38794 24058 38794 0 gencon_inst.ALU_out\[3\]
rlabel metal1 27462 36686 27462 36686 0 gencon_inst.ALU_out\[4\]
rlabel metal1 27968 37094 27968 37094 0 gencon_inst.ALU_out\[5\]
rlabel metal2 30130 34833 30130 34833 0 gencon_inst.ALU_out\[6\]
rlabel metal1 30130 36550 30130 36550 0 gencon_inst.ALU_out\[7\]
rlabel metal2 23046 35955 23046 35955 0 gencon_inst.ALU_out\[8\]
rlabel metal2 33902 38641 33902 38641 0 gencon_inst.ALU_out\[9\]
rlabel metal2 13110 33252 13110 33252 0 gencon_inst.addOrSub
rlabel metal2 16790 36550 16790 36550 0 gencon_inst.add_calc.diffSign
rlabel metal2 40986 39236 40986 39236 0 gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1
rlabel metal2 42182 36788 42182 36788 0 gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1
rlabel metal1 39008 36142 39008 36142 0 gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1
rlabel metal1 34454 35598 34454 35598 0 gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1
rlabel metal2 31510 34918 31510 34918 0 gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1
rlabel metal2 18814 40800 18814 40800 0 gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1
rlabel metal1 21344 42330 21344 42330 0 gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1
rlabel metal1 23276 41990 23276 41990 0 gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1
rlabel metal1 26864 35598 26864 35598 0 gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1
rlabel metal1 26450 41208 26450 41208 0 gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1
rlabel metal2 29026 42364 29026 42364 0 gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1
rlabel metal1 31372 41786 31372 41786 0 gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1
rlabel metal1 34362 42670 34362 42670 0 gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1
rlabel metal2 37490 41854 37490 41854 0 gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1
rlabel metal1 17802 38998 17802 38998 0 gencon_inst.add_calc.main.a0.in1
rlabel metal1 16882 38828 16882 38828 0 gencon_inst.add_calc.main.in2\[0\]
rlabel metal2 42182 38964 42182 38964 0 gencon_inst.add_calc.main.in2\[10\]
rlabel metal1 41745 36686 41745 36686 0 gencon_inst.add_calc.main.in2\[11\]
rlabel metal1 39514 35700 39514 35700 0 gencon_inst.add_calc.main.in2\[12\]
rlabel metal2 33810 34612 33810 34612 0 gencon_inst.add_calc.main.in2\[13\]
rlabel metal1 30314 36176 30314 36176 0 gencon_inst.add_calc.main.in2\[14\]
rlabel metal2 16882 40868 16882 40868 0 gencon_inst.add_calc.main.in2\[1\]
rlabel metal1 21206 42262 21206 42262 0 gencon_inst.add_calc.main.in2\[2\]
rlabel metal1 23920 41106 23920 41106 0 gencon_inst.add_calc.main.in2\[3\]
rlabel metal1 25438 37230 25438 37230 0 gencon_inst.add_calc.main.in2\[4\]
rlabel metal1 26174 42330 26174 42330 0 gencon_inst.add_calc.main.in2\[5\]
rlabel metal1 28980 35258 28980 35258 0 gencon_inst.add_calc.main.in2\[6\]
rlabel metal2 31786 42466 31786 42466 0 gencon_inst.add_calc.main.in2\[7\]
rlabel metal2 33902 43044 33902 43044 0 gencon_inst.add_calc.main.in2\[8\]
rlabel metal1 38732 42126 38732 42126 0 gencon_inst.add_calc.main.in2\[9\]
rlabel metal1 13800 34170 13800 34170 0 gencon_inst.add_calc.next_finish
rlabel metal1 17158 36686 17158 36686 0 gencon_inst.add_calc.sameSignVal
rlabel metal2 12374 33252 12374 33252 0 gencon_inst.add_calc.start
rlabel metal1 13731 35802 13731 35802 0 gencon_inst.add_calc.state\[0\]
rlabel metal2 18814 37723 18814 37723 0 gencon_inst.add_calc.state\[1\]
rlabel metal1 15226 36346 15226 36346 0 gencon_inst.add_calc.state\[2\]
rlabel metal1 15410 27982 15410 27982 0 gencon_inst.gencon_state\[0\]
rlabel metal1 19550 26894 19550 26894 0 gencon_inst.gencon_state\[1\]
rlabel via1 17789 26282 17789 26282 0 gencon_inst.gencon_state\[2\]
rlabel metal1 19734 26452 19734 26452 0 gencon_inst.gencon_state\[3\]
rlabel metal1 15502 25330 15502 25330 0 gencon_inst.key_read
rlabel metal1 7636 27846 7636 27846 0 gencon_inst.keypad_input\[0\]
rlabel metal1 9522 26010 9522 26010 0 gencon_inst.keypad_input\[1\]
rlabel metal1 9062 26758 9062 26758 0 gencon_inst.keypad_input\[2\]
rlabel metal2 9062 27676 9062 27676 0 gencon_inst.keypad_input\[3\]
rlabel metal2 19826 29410 19826 29410 0 gencon_inst.latched_keypad_input\[0\]
rlabel metal1 19596 24786 19596 24786 0 gencon_inst.latched_keypad_input\[1\]
rlabel metal1 20930 28526 20930 28526 0 gencon_inst.latched_keypad_input\[2\]
rlabel metal1 13846 28526 13846 28526 0 gencon_inst.latched_keypad_input\[3\]
rlabel metal1 13708 31246 13708 31246 0 gencon_inst.latched_operator_input\[0\]
rlabel metal2 13570 30464 13570 30464 0 gencon_inst.latched_operator_input\[1\]
rlabel metal1 13708 30022 13708 30022 0 gencon_inst.latched_operator_input\[2\]
rlabel metal1 17158 15674 17158 15674 0 gencon_inst.mult_calc.INn1\[0\]
rlabel metal1 41699 21454 41699 21454 0 gencon_inst.mult_calc.INn1\[10\]
rlabel metal2 41354 21828 41354 21828 0 gencon_inst.mult_calc.INn1\[11\]
rlabel metal2 38686 22100 38686 22100 0 gencon_inst.mult_calc.INn1\[12\]
rlabel metal1 41308 22202 41308 22202 0 gencon_inst.mult_calc.INn1\[13\]
rlabel metal2 31878 15300 31878 15300 0 gencon_inst.mult_calc.INn1\[14\]
rlabel metal1 16422 20366 16422 20366 0 gencon_inst.mult_calc.INn1\[15\]
rlabel metal1 18446 17748 18446 17748 0 gencon_inst.mult_calc.INn1\[1\]
rlabel metal1 22770 21114 22770 21114 0 gencon_inst.mult_calc.INn1\[2\]
rlabel metal1 24564 22066 24564 22066 0 gencon_inst.mult_calc.INn1\[3\]
rlabel metal1 25254 22542 25254 22542 0 gencon_inst.mult_calc.INn1\[4\]
rlabel metal2 26726 19108 26726 19108 0 gencon_inst.mult_calc.INn1\[5\]
rlabel metal1 28658 23630 28658 23630 0 gencon_inst.mult_calc.INn1\[6\]
rlabel metal1 30406 21658 30406 21658 0 gencon_inst.mult_calc.INn1\[7\]
rlabel metal1 33350 19924 33350 19924 0 gencon_inst.mult_calc.INn1\[8\]
rlabel metal2 39054 20026 39054 20026 0 gencon_inst.mult_calc.INn1\[9\]
rlabel metal1 19826 11866 19826 11866 0 gencon_inst.mult_calc.INn2\[0\]
rlabel metal2 32706 11458 32706 11458 0 gencon_inst.mult_calc.INn2\[10\]
rlabel metal1 34132 20230 34132 20230 0 gencon_inst.mult_calc.INn2\[11\]
rlabel metal1 34914 20774 34914 20774 0 gencon_inst.mult_calc.INn2\[12\]
rlabel metal1 36524 19686 36524 19686 0 gencon_inst.mult_calc.INn2\[13\]
rlabel metal1 33672 20774 33672 20774 0 gencon_inst.mult_calc.INn2\[14\]
rlabel metal1 15824 21114 15824 21114 0 gencon_inst.mult_calc.INn2\[15\]
rlabel metal1 21114 21454 21114 21454 0 gencon_inst.mult_calc.INn2\[1\]
rlabel metal1 20930 11798 20930 11798 0 gencon_inst.mult_calc.INn2\[2\]
rlabel metal2 22816 16932 22816 16932 0 gencon_inst.mult_calc.INn2\[3\]
rlabel metal1 26588 21454 26588 21454 0 gencon_inst.mult_calc.INn2\[4\]
rlabel metal1 27554 21862 27554 21862 0 gencon_inst.mult_calc.INn2\[5\]
rlabel metal1 27784 21046 27784 21046 0 gencon_inst.mult_calc.INn2\[6\]
rlabel metal2 27232 17238 27232 17238 0 gencon_inst.mult_calc.INn2\[7\]
rlabel metal1 32108 20774 32108 20774 0 gencon_inst.mult_calc.INn2\[8\]
rlabel via2 33534 21845 33534 21845 0 gencon_inst.mult_calc.INn2\[9\]
rlabel metal2 18446 14484 18446 14484 0 gencon_inst.mult_calc.adderSave\[0\]
rlabel metal2 41446 17850 41446 17850 0 gencon_inst.mult_calc.adderSave\[10\]
rlabel metal1 39928 17714 39928 17714 0 gencon_inst.mult_calc.adderSave\[11\]
rlabel metal1 39560 14926 39560 14926 0 gencon_inst.mult_calc.adderSave\[12\]
rlabel metal1 38916 12274 38916 12274 0 gencon_inst.mult_calc.adderSave\[13\]
rlabel metal1 35098 14042 35098 14042 0 gencon_inst.mult_calc.adderSave\[14\]
rlabel metal1 19964 15878 19964 15878 0 gencon_inst.mult_calc.adderSave\[1\]
rlabel metal2 22126 16830 22126 16830 0 gencon_inst.mult_calc.adderSave\[2\]
rlabel metal2 21666 14348 21666 14348 0 gencon_inst.mult_calc.adderSave\[3\]
rlabel metal1 24610 17714 24610 17714 0 gencon_inst.mult_calc.adderSave\[4\]
rlabel metal2 25622 14484 25622 14484 0 gencon_inst.mult_calc.adderSave\[5\]
rlabel metal1 30314 14892 30314 14892 0 gencon_inst.mult_calc.adderSave\[6\]
rlabel metal2 28750 17340 28750 17340 0 gencon_inst.mult_calc.adderSave\[7\]
rlabel metal1 30176 16422 30176 16422 0 gencon_inst.mult_calc.adderSave\[8\]
rlabel metal2 35282 16388 35282 16388 0 gencon_inst.mult_calc.adderSave\[9\]
rlabel metal1 20470 11186 20470 11186 0 gencon_inst.mult_calc.compCount.in2\[0\]
rlabel metal1 32706 9078 32706 9078 0 gencon_inst.mult_calc.compCount.in2\[10\]
rlabel metal1 35604 9486 35604 9486 0 gencon_inst.mult_calc.compCount.in2\[11\]
rlabel metal1 37398 11322 37398 11322 0 gencon_inst.mult_calc.compCount.in2\[12\]
rlabel metal1 36340 11866 36340 11866 0 gencon_inst.mult_calc.compCount.in2\[13\]
rlabel metal1 34822 12750 34822 12750 0 gencon_inst.mult_calc.compCount.in2\[14\]
rlabel metal1 20010 9622 20010 9622 0 gencon_inst.mult_calc.compCount.in2\[1\]
rlabel metal2 21482 10914 21482 10914 0 gencon_inst.mult_calc.compCount.in2\[2\]
rlabel metal2 24150 11356 24150 11356 0 gencon_inst.mult_calc.compCount.in2\[3\]
rlabel metal2 25530 9860 25530 9860 0 gencon_inst.mult_calc.compCount.in2\[4\]
rlabel metal1 26680 11186 26680 11186 0 gencon_inst.mult_calc.compCount.in2\[5\]
rlabel metal2 28014 10642 28014 10642 0 gencon_inst.mult_calc.compCount.in2\[6\]
rlabel metal2 29118 9656 29118 9656 0 gencon_inst.mult_calc.compCount.in2\[7\]
rlabel metal1 31464 11254 31464 11254 0 gencon_inst.mult_calc.compCount.in2\[8\]
rlabel metal1 33994 12750 33994 12750 0 gencon_inst.mult_calc.compCount.in2\[9\]
rlabel metal1 34408 7174 34408 7174 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1
rlabel metal2 33258 5882 33258 5882 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1
rlabel metal2 37030 6324 37030 6324 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1
rlabel metal2 37398 8058 37398 8058 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1
rlabel metal1 37766 9452 37766 9452 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[14\].thingy.in1
rlabel metal1 21482 9010 21482 9010 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
rlabel metal2 20378 8466 20378 8466 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1
rlabel metal1 21758 8840 21758 8840 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1
rlabel metal1 22862 6630 22862 6630 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1
rlabel metal1 26128 8058 26128 8058 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1
rlabel metal1 25254 7854 25254 7854 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1
rlabel metal1 28336 7310 28336 7310 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1
rlabel metal1 31234 6290 31234 6290 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1
rlabel metal1 31142 7310 31142 7310 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1
rlabel metal1 32890 5134 32890 5134 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1
rlabel metal2 20194 6868 20194 6868 0 gencon_inst.mult_calc.countSave\[0\]
rlabel metal2 33902 8092 33902 8092 0 gencon_inst.mult_calc.countSave\[10\]
rlabel metal1 34730 6834 34730 6834 0 gencon_inst.mult_calc.countSave\[11\]
rlabel metal1 37352 6426 37352 6426 0 gencon_inst.mult_calc.countSave\[12\]
rlabel metal1 38594 7990 38594 7990 0 gencon_inst.mult_calc.countSave\[13\]
rlabel metal1 40020 10574 40020 10574 0 gencon_inst.mult_calc.countSave\[14\]
rlabel metal1 19182 7922 19182 7922 0 gencon_inst.mult_calc.countSave\[1\]
rlabel metal2 22218 10404 22218 10404 0 gencon_inst.mult_calc.countSave\[2\]
rlabel metal1 21942 6290 21942 6290 0 gencon_inst.mult_calc.countSave\[3\]
rlabel metal1 25530 6426 25530 6426 0 gencon_inst.mult_calc.countSave\[4\]
rlabel metal1 25944 9486 25944 9486 0 gencon_inst.mult_calc.countSave\[5\]
rlabel metal1 28152 6766 28152 6766 0 gencon_inst.mult_calc.countSave\[6\]
rlabel metal2 29946 5780 29946 5780 0 gencon_inst.mult_calc.countSave\[7\]
rlabel metal1 29486 8398 29486 8398 0 gencon_inst.mult_calc.countSave\[8\]
rlabel metal1 33488 5746 33488 5746 0 gencon_inst.mult_calc.countSave\[9\]
rlabel metal2 17250 19244 17250 19244 0 gencon_inst.mult_calc.diffSign
rlabel metal1 17020 13362 17020 13362 0 gencon_inst.mult_calc.finish
rlabel metal1 40986 19346 40986 19346 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1
rlabel metal2 41078 18802 41078 18802 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2
rlabel metal2 42182 20026 42182 20026 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1
rlabel metal1 41952 17170 41952 17170 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2
rlabel metal2 39514 14144 39514 14144 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1
rlabel metal2 41446 15300 41446 15300 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2
rlabel metal2 42182 13668 42182 13668 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1
rlabel metal1 40986 12750 40986 12750 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2
rlabel metal1 34178 14246 34178 14246 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in1
rlabel metal2 33074 13702 33074 13702 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in2
rlabel metal1 18906 16558 18906 16558 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1
rlabel metal1 19780 15470 19780 15470 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2
rlabel metal2 21850 16626 21850 16626 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1
rlabel metal2 22034 16626 22034 16626 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2
rlabel metal2 23782 19516 23782 19516 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1
rlabel metal2 22402 14212 22402 14212 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2
rlabel metal2 25806 20740 25806 20740 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1
rlabel metal1 26220 17102 26220 17102 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2
rlabel metal1 27278 17850 27278 17850 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1
rlabel metal2 26726 14076 26726 14076 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2
rlabel metal1 28658 15878 28658 15878 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1
rlabel metal2 28382 14586 28382 14586 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2
rlabel metal2 30130 20910 30130 20910 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1
rlabel metal1 30544 17646 30544 17646 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2
rlabel metal2 32154 19924 32154 19924 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1
rlabel metal1 32936 17714 32936 17714 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2
rlabel metal1 37444 18802 37444 18802 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
rlabel metal1 35052 17578 35052 17578 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2
rlabel metal2 18906 14892 18906 14892 0 gencon_inst.mult_calc.main.a0.in1
rlabel metal2 20562 14926 20562 14926 0 gencon_inst.mult_calc.main.a0.in2
rlabel metal2 28566 13328 28566 13328 0 gencon_inst.mult_calc.next_finish
rlabel metal1 19366 19278 19366 19278 0 gencon_inst.mult_calc.out\[0\]
rlabel metal1 36294 18394 36294 18394 0 gencon_inst.mult_calc.out\[10\]
rlabel metal1 36432 18598 36432 18598 0 gencon_inst.mult_calc.out\[11\]
rlabel metal1 37076 15674 37076 15674 0 gencon_inst.mult_calc.out\[12\]
rlabel metal1 37076 13430 37076 13430 0 gencon_inst.mult_calc.out\[13\]
rlabel metal1 32062 13838 32062 13838 0 gencon_inst.mult_calc.out\[14\]
rlabel metal1 18538 20570 18538 20570 0 gencon_inst.mult_calc.out\[15\]
rlabel metal1 19964 18394 19964 18394 0 gencon_inst.mult_calc.out\[1\]
rlabel metal1 21298 19278 21298 19278 0 gencon_inst.mult_calc.out\[2\]
rlabel metal1 23736 13430 23736 13430 0 gencon_inst.mult_calc.out\[3\]
rlabel metal1 25530 19482 25530 19482 0 gencon_inst.mult_calc.out\[4\]
rlabel metal1 25944 14042 25944 14042 0 gencon_inst.mult_calc.out\[5\]
rlabel metal1 27784 20570 27784 20570 0 gencon_inst.mult_calc.out\[6\]
rlabel metal1 29716 19278 29716 19278 0 gencon_inst.mult_calc.out\[7\]
rlabel metal1 31234 18734 31234 18734 0 gencon_inst.mult_calc.out\[8\]
rlabel metal1 33718 18394 33718 18394 0 gencon_inst.mult_calc.out\[9\]
rlabel metal2 16514 15572 16514 15572 0 gencon_inst.mult_calc.start
rlabel via1 17595 11322 17595 11322 0 gencon_inst.mult_calc.state\[0\]
rlabel metal1 30590 12138 30590 12138 0 gencon_inst.mult_calc.state\[2\]
rlabel metal1 19274 11594 19274 11594 0 gencon_inst.mult_calc.state\[3\]
rlabel metal1 34086 14926 34086 14926 0 gencon_inst.mult_calc.state\[4\]
rlabel metal2 14490 27778 14490 27778 0 gencon_inst.next_state\[0\]
rlabel metal1 15594 27098 15594 27098 0 gencon_inst.next_state\[1\]
rlabel metal2 15870 25500 15870 25500 0 gencon_inst.next_state\[2\]
rlabel metal1 15134 28186 15134 28186 0 gencon_inst.next_state\[3\]
rlabel metal1 17986 31994 17986 31994 0 gencon_inst.operand1\[0\]
rlabel metal2 39054 29580 39054 29580 0 gencon_inst.operand1\[10\]
rlabel metal3 40365 33252 40365 33252 0 gencon_inst.operand1\[11\]
rlabel metal1 37260 31654 37260 31654 0 gencon_inst.operand1\[12\]
rlabel metal2 33856 29138 33856 29138 0 gencon_inst.operand1\[13\]
rlabel metal1 34086 28934 34086 28934 0 gencon_inst.operand1\[14\]
rlabel metal1 16468 31450 16468 31450 0 gencon_inst.operand1\[15\]
rlabel metal2 19458 28832 19458 28832 0 gencon_inst.operand1\[1\]
rlabel metal1 21206 28560 21206 28560 0 gencon_inst.operand1\[2\]
rlabel metal2 23276 34918 23276 34918 0 gencon_inst.operand1\[3\]
rlabel metal2 25254 30226 25254 30226 0 gencon_inst.operand1\[4\]
rlabel metal2 26818 30804 26818 30804 0 gencon_inst.operand1\[5\]
rlabel metal1 27600 32402 27600 32402 0 gencon_inst.operand1\[6\]
rlabel metal2 30130 30124 30130 30124 0 gencon_inst.operand1\[7\]
rlabel metal1 35006 32810 35006 32810 0 gencon_inst.operand1\[8\]
rlabel metal2 38410 28628 38410 28628 0 gencon_inst.operand1\[9\]
rlabel metal1 18170 20842 18170 20842 0 gencon_inst.operand2\[0\]
rlabel metal1 34868 21930 34868 21930 0 gencon_inst.operand2\[10\]
rlabel metal1 41722 33490 41722 33490 0 gencon_inst.operand2\[11\]
rlabel metal1 35098 21590 35098 21590 0 gencon_inst.operand2\[12\]
rlabel metal1 33166 20502 33166 20502 0 gencon_inst.operand2\[13\]
rlabel metal1 32798 21862 32798 21862 0 gencon_inst.operand2\[14\]
rlabel metal1 15410 21998 15410 21998 0 gencon_inst.operand2\[15\]
rlabel metal1 19504 31722 19504 31722 0 gencon_inst.operand2\[1\]
rlabel metal2 20746 23528 20746 23528 0 gencon_inst.operand2\[2\]
rlabel metal1 21114 22678 21114 22678 0 gencon_inst.operand2\[3\]
rlabel metal1 25300 33490 25300 33490 0 gencon_inst.operand2\[4\]
rlabel metal1 26358 32436 26358 32436 0 gencon_inst.operand2\[5\]
rlabel metal1 25990 20502 25990 20502 0 gencon_inst.operand2\[6\]
rlabel metal1 30268 32402 30268 32402 0 gencon_inst.operand2\[7\]
rlabel metal1 32614 26010 32614 26010 0 gencon_inst.operand2\[8\]
rlabel metal1 32660 21386 32660 21386 0 gencon_inst.operand2\[9\]
rlabel metal1 13156 30566 13156 30566 0 gencon_inst.operator_input\[0\]
rlabel metal1 12512 25874 12512 25874 0 gencon_inst.operator_input\[1\]
rlabel metal1 12788 25874 12788 25874 0 gencon_inst.operator_input\[2\]
rlabel metal1 13248 23834 13248 23834 0 gencon_inst.prev_operator_input\[0\]
rlabel metal1 13248 23086 13248 23086 0 gencon_inst.prev_operator_input\[1\]
rlabel metal1 13110 24378 13110 24378 0 gencon_inst.prev_operator_input\[2\]
rlabel metal1 14030 21862 14030 21862 0 gencon_inst.prev_read_input
rlabel metal2 11178 21760 11178 21760 0 gencon_inst.read_input
rlabel metal1 3105 13498 3105 13498 0 input_ctrl_inst.RowMid\[0\]
rlabel metal1 3795 14382 3795 14382 0 input_ctrl_inst.RowMid\[1\]
rlabel metal1 3795 16626 3795 16626 0 input_ctrl_inst.RowMid\[2\]
rlabel metal1 3795 17646 3795 17646 0 input_ctrl_inst.RowMid\[3\]
rlabel metal2 4830 16116 4830 16116 0 input_ctrl_inst.RowSync\[0\]
rlabel metal2 4646 16048 4646 16048 0 input_ctrl_inst.RowSync\[1\]
rlabel metal2 5382 16847 5382 16847 0 input_ctrl_inst.RowSync\[2\]
rlabel metal1 5060 17578 5060 17578 0 input_ctrl_inst.RowSync\[3\]
rlabel metal2 5750 16439 5750 16439 0 input_ctrl_inst.col_index\[0\]
rlabel metal1 3864 7854 3864 7854 0 input_ctrl_inst.col_index\[10\]
rlabel metal1 3864 7718 3864 7718 0 input_ctrl_inst.col_index\[11\]
rlabel metal1 5612 6630 5612 6630 0 input_ctrl_inst.col_index\[12\]
rlabel metal1 6394 6698 6394 6698 0 input_ctrl_inst.col_index\[13\]
rlabel metal1 5888 6086 5888 6086 0 input_ctrl_inst.col_index\[14\]
rlabel metal1 6992 5134 6992 5134 0 input_ctrl_inst.col_index\[15\]
rlabel metal2 7498 6426 7498 6426 0 input_ctrl_inst.col_index\[16\]
rlabel metal2 9154 5508 9154 5508 0 input_ctrl_inst.col_index\[17\]
rlabel metal1 8802 6698 8802 6698 0 input_ctrl_inst.col_index\[18\]
rlabel metal1 9154 7786 9154 7786 0 input_ctrl_inst.col_index\[19\]
rlabel metal1 6486 20366 6486 20366 0 input_ctrl_inst.col_index\[1\]
rlabel metal2 11270 8126 11270 8126 0 input_ctrl_inst.col_index\[20\]
rlabel metal2 12466 7922 12466 7922 0 input_ctrl_inst.col_index\[21\]
rlabel metal1 12880 7446 12880 7446 0 input_ctrl_inst.col_index\[22\]
rlabel metal2 11914 7140 11914 7140 0 input_ctrl_inst.col_index\[23\]
rlabel metal2 9706 11118 9706 11118 0 input_ctrl_inst.col_index\[24\]
rlabel metal1 12972 11050 12972 11050 0 input_ctrl_inst.col_index\[25\]
rlabel metal1 12466 11594 12466 11594 0 input_ctrl_inst.col_index\[26\]
rlabel metal2 13294 10268 13294 10268 0 input_ctrl_inst.col_index\[27\]
rlabel metal1 13570 12172 13570 12172 0 input_ctrl_inst.col_index\[28\]
rlabel metal1 12466 12308 12466 12308 0 input_ctrl_inst.col_index\[29\]
rlabel metal2 6118 16626 6118 16626 0 input_ctrl_inst.col_index\[2\]
rlabel metal1 12650 12138 12650 12138 0 input_ctrl_inst.col_index\[30\]
rlabel metal1 12006 12274 12006 12274 0 input_ctrl_inst.col_index\[31\]
rlabel metal1 6440 16762 6440 16762 0 input_ctrl_inst.col_index\[3\]
rlabel metal1 5382 10574 5382 10574 0 input_ctrl_inst.col_index\[4\]
rlabel metal1 4462 12818 4462 12818 0 input_ctrl_inst.col_index\[5\]
rlabel metal1 3588 12750 3588 12750 0 input_ctrl_inst.col_index\[6\]
rlabel metal2 4186 10982 4186 10982 0 input_ctrl_inst.col_index\[7\]
rlabel metal1 3634 9078 3634 9078 0 input_ctrl_inst.col_index\[8\]
rlabel metal2 3634 7582 3634 7582 0 input_ctrl_inst.col_index\[9\]
rlabel metal1 8326 29478 8326 29478 0 input_ctrl_inst.debounce_cnt\[0\]
rlabel metal1 4784 36006 4784 36006 0 input_ctrl_inst.debounce_cnt\[10\]
rlabel metal1 4876 34986 4876 34986 0 input_ctrl_inst.debounce_cnt\[11\]
rlabel metal2 5382 33966 5382 33966 0 input_ctrl_inst.debounce_cnt\[12\]
rlabel metal1 5888 33558 5888 33558 0 input_ctrl_inst.debounce_cnt\[13\]
rlabel metal1 5198 32300 5198 32300 0 input_ctrl_inst.debounce_cnt\[14\]
rlabel metal1 2806 30192 2806 30192 0 input_ctrl_inst.debounce_cnt\[15\]
rlabel metal1 3496 31246 3496 31246 0 input_ctrl_inst.debounce_cnt\[16\]
rlabel metal1 2300 29546 2300 29546 0 input_ctrl_inst.debounce_cnt\[17\]
rlabel metal2 4186 29427 4186 29427 0 input_ctrl_inst.debounce_cnt\[18\]
rlabel metal2 10442 30396 10442 30396 0 input_ctrl_inst.debounce_cnt\[1\]
rlabel metal2 8786 31042 8786 31042 0 input_ctrl_inst.debounce_cnt\[2\]
rlabel metal1 8970 31212 8970 31212 0 input_ctrl_inst.debounce_cnt\[3\]
rlabel metal1 10580 32878 10580 32878 0 input_ctrl_inst.debounce_cnt\[4\]
rlabel metal1 9936 34714 9936 34714 0 input_ctrl_inst.debounce_cnt\[5\]
rlabel metal1 8556 34170 8556 34170 0 input_ctrl_inst.debounce_cnt\[6\]
rlabel metal1 7130 35054 7130 35054 0 input_ctrl_inst.debounce_cnt\[7\]
rlabel metal1 9982 35598 9982 35598 0 input_ctrl_inst.debounce_cnt\[8\]
rlabel metal1 6946 34918 6946 34918 0 input_ctrl_inst.debounce_cnt\[9\]
rlabel metal1 7636 23698 7636 23698 0 input_ctrl_inst.decoded_key\[0\]
rlabel metal1 7291 21318 7291 21318 0 input_ctrl_inst.decoded_key\[1\]
rlabel metal1 9890 24752 9890 24752 0 input_ctrl_inst.decoded_key\[2\]
rlabel metal1 5014 22406 5014 22406 0 input_ctrl_inst.decoded_key\[3\]
rlabel metal1 3634 23596 3634 23596 0 input_ctrl_inst.input_control_state\[0\]
rlabel metal1 3726 24174 3726 24174 0 input_ctrl_inst.input_control_state\[1\]
rlabel metal1 5014 26282 5014 26282 0 input_ctrl_inst.input_control_state\[2\]
rlabel metal1 3367 26554 3367 26554 0 input_ctrl_inst.next_state\[0\]
rlabel metal2 2162 23834 2162 23834 0 input_ctrl_inst.next_state\[1\]
rlabel metal1 5152 26554 5152 26554 0 input_ctrl_inst.next_state\[2\]
rlabel metal2 8878 21284 8878 21284 0 input_ctrl_inst.read_input_flag
rlabel metal1 9614 18088 9614 18088 0 input_ctrl_inst.scan_timer\[0\]
rlabel metal1 12926 15436 12926 15436 0 input_ctrl_inst.scan_timer\[10\]
rlabel metal1 11822 16524 11822 16524 0 input_ctrl_inst.scan_timer\[11\]
rlabel metal1 10534 14926 10534 14926 0 input_ctrl_inst.scan_timer\[12\]
rlabel metal1 9890 15538 9890 15538 0 input_ctrl_inst.scan_timer\[13\]
rlabel metal2 9430 16218 9430 16218 0 input_ctrl_inst.scan_timer\[14\]
rlabel metal1 8970 17510 8970 17510 0 input_ctrl_inst.scan_timer\[15\]
rlabel metal1 4508 20026 4508 20026 0 input_ctrl_inst.scan_timer\[16\]
rlabel metal1 3772 20026 3772 20026 0 input_ctrl_inst.scan_timer\[17\]
rlabel metal1 3864 19822 3864 19822 0 input_ctrl_inst.scan_timer\[18\]
rlabel metal1 4186 20910 4186 20910 0 input_ctrl_inst.scan_timer\[19\]
rlabel metal2 8878 19550 8878 19550 0 input_ctrl_inst.scan_timer\[1\]
rlabel metal1 10902 21012 10902 21012 0 input_ctrl_inst.scan_timer\[2\]
rlabel metal2 10902 19108 10902 19108 0 input_ctrl_inst.scan_timer\[3\]
rlabel metal2 13202 19176 13202 19176 0 input_ctrl_inst.scan_timer\[4\]
rlabel metal1 13248 20570 13248 20570 0 input_ctrl_inst.scan_timer\[5\]
rlabel metal2 12558 17952 12558 17952 0 input_ctrl_inst.scan_timer\[6\]
rlabel metal1 13938 17748 13938 17748 0 input_ctrl_inst.scan_timer\[7\]
rlabel metal1 12742 17204 12742 17204 0 input_ctrl_inst.scan_timer\[8\]
rlabel metal2 12788 16422 12788 16422 0 input_ctrl_inst.scan_timer\[9\]
rlabel metal1 1472 24650 1472 24650 0 input_state_FPGA[0]
rlabel metal3 1142 23188 1142 23188 0 input_state_FPGA[1]
rlabel metal1 1472 21862 1472 21862 0 input_state_FPGA[2]
rlabel metal3 751 27948 751 27948 0 key_pressed
rlabel metal2 42090 5559 42090 5559 0 nRST
rlabel metal1 1702 13362 1702 13362 0 net1
rlabel metal1 1702 25942 1702 25942 0 net10
rlabel metal1 34638 19210 34638 19210 0 net100
rlabel metal2 41722 20196 41722 20196 0 net101
rlabel metal2 38410 14314 38410 14314 0 net102
rlabel metal1 19964 14314 19964 14314 0 net103
rlabel metal1 17204 12206 17204 12206 0 net104
rlabel metal2 36570 13838 36570 13838 0 net105
rlabel metal1 21574 42194 21574 42194 0 net106
rlabel metal1 32890 42262 32890 42262 0 net107
rlabel metal2 40250 40902 40250 40902 0 net108
rlabel metal1 17802 36822 17802 36822 0 net109
rlabel metal1 20976 43282 20976 43282 0 net11
rlabel metal1 19918 42772 19918 42772 0 net110
rlabel metal1 24978 37264 24978 37264 0 net111
rlabel metal1 33718 42092 33718 42092 0 net112
rlabel metal1 41630 38930 41630 38930 0 net113
rlabel metal1 13524 35666 13524 35666 0 net114
rlabel metal2 34178 37536 34178 37536 0 net115
rlabel metal1 5152 16490 5152 16490 0 net116
rlabel metal1 6946 12240 6946 12240 0 net117
rlabel metal2 14030 24446 14030 24446 0 net118
rlabel metal1 16698 16218 16698 16218 0 net119
rlabel via1 41814 30906 41814 30906 0 net12
rlabel metal1 4607 13974 4607 13974 0 net120
rlabel metal2 10350 13600 10350 13600 0 net121
rlabel metal1 3135 12886 3135 12886 0 net122
rlabel metal1 6532 19686 6532 19686 0 net123
rlabel metal2 2438 22848 2438 22848 0 net124
rlabel metal2 7958 15266 7958 15266 0 net125
rlabel metal1 20937 6698 20937 6698 0 net126
rlabel metal1 17342 11832 17342 11832 0 net127
rlabel metal1 15909 16490 15909 16490 0 net128
rlabel metal1 20785 19754 20785 19754 0 net129
rlabel metal1 39790 22644 39790 22644 0 net13
rlabel metal2 17986 6595 17986 6595 0 net130
rlabel metal2 2806 28322 2806 28322 0 net131
rlabel metal1 10534 31831 10534 31831 0 net132
rlabel metal2 12742 28050 12742 28050 0 net133
rlabel metal1 17303 25194 17303 25194 0 net134
rlabel metal1 19741 32470 19741 32470 0 net135
rlabel metal2 16146 39678 16146 39678 0 net136
rlabel metal2 20286 41888 20286 41888 0 net137
rlabel metal2 22034 34357 22034 34357 0 net138
rlabel metal2 22862 13770 22862 13770 0 net139
rlabel metal1 42044 32402 42044 32402 0 net14
rlabel metal1 21926 13226 21926 13226 0 net140
rlabel metal1 28389 14314 28389 14314 0 net141
rlabel metal2 30406 13600 30406 13600 0 net142
rlabel metal1 25077 20502 25077 20502 0 net143
rlabel metal1 28849 17578 28849 17578 0 net144
rlabel metal1 32062 17170 32062 17170 0 net145
rlabel metal1 35006 9445 35006 9445 0 net146
rlabel metal1 35420 12954 35420 12954 0 net147
rlabel metal1 36655 12886 36655 12886 0 net148
rlabel metal2 41630 16116 41630 16116 0 net149
rlabel metal2 40618 25296 40618 25296 0 net15
rlabel metal1 41860 15402 41860 15402 0 net150
rlabel metal2 41446 10251 41446 10251 0 net151
rlabel metal1 26089 27370 26089 27370 0 net152
rlabel metal1 23835 38998 23835 38998 0 net153
rlabel metal1 29946 36713 29946 36713 0 net154
rlabel metal1 31234 34544 31234 34544 0 net155
rlabel metal1 40427 27370 40427 27370 0 net156
rlabel metal2 33810 25432 33810 25432 0 net157
rlabel metal2 34362 42466 34362 42466 0 net158
rlabel metal1 38173 41514 38173 41514 0 net159
rlabel metal1 40342 29172 40342 29172 0 net16
rlabel metal2 41814 33473 41814 33473 0 net160
rlabel metal2 3082 17340 3082 17340 0 net161
rlabel metal2 2990 16252 2990 16252 0 net162
rlabel metal2 3818 14756 3818 14756 0 net163
rlabel metal1 2300 14042 2300 14042 0 net164
rlabel metal2 14490 22644 14490 22644 0 net165
rlabel metal2 32798 15266 32798 15266 0 net166
rlabel metal1 30176 21862 30176 21862 0 net167
rlabel metal1 17296 17714 17296 17714 0 net168
rlabel metal1 40848 20434 40848 20434 0 net169
rlabel metal1 20010 43282 20010 43282 0 net17
rlabel metal1 32982 14994 32982 14994 0 net170
rlabel metal1 22356 21522 22356 21522 0 net171
rlabel metal1 26680 19346 26680 19346 0 net172
rlabel metal2 3450 20604 3450 20604 0 net173
rlabel metal1 2341 20910 2341 20910 0 net174
rlabel metal1 14076 23698 14076 23698 0 net175
rlabel metal1 24840 20978 24840 20978 0 net176
rlabel metal1 41814 20570 41814 20570 0 net177
rlabel metal1 33442 19686 33442 19686 0 net178
rlabel metal2 39606 19550 39606 19550 0 net179
rlabel metal1 21298 43214 21298 43214 0 net18
rlabel metal2 18170 15776 18170 15776 0 net180
rlabel metal1 40940 18938 40940 18938 0 net181
rlabel metal1 21942 20434 21942 20434 0 net182
rlabel metal2 29946 21114 29946 21114 0 net183
rlabel metal1 14214 24106 14214 24106 0 net184
rlabel metal1 26634 18258 26634 18258 0 net185
rlabel metal1 17480 17306 17480 17306 0 net186
rlabel metal1 34178 19414 34178 19414 0 net187
rlabel metal1 23414 21862 23414 21862 0 net188
rlabel metal2 41538 19958 41538 19958 0 net189
rlabel metal1 23046 33082 23046 33082 0 net19
rlabel metal2 12650 22848 12650 22848 0 net190
rlabel metal1 25024 20842 25024 20842 0 net191
rlabel metal1 10396 27370 10396 27370 0 net192
rlabel metal1 38226 18938 38226 18938 0 net193
rlabel metal2 17986 14790 17986 14790 0 net194
rlabel metal1 40388 29546 40388 29546 0 net195
rlabel metal2 2806 23868 2806 23868 0 net196
rlabel metal1 16192 20842 16192 20842 0 net197
rlabel metal1 23276 18734 23276 18734 0 net198
rlabel metal2 15594 21828 15594 21828 0 net199
rlabel metal1 1748 14382 1748 14382 0 net2
rlabel metal2 23506 33201 23506 33201 0 net20
rlabel via1 14393 20842 14393 20842 0 net200
rlabel metal2 4554 20706 4554 20706 0 net201
rlabel metal1 5244 19346 5244 19346 0 net202
rlabel metal1 40802 33966 40802 33966 0 net203
rlabel metal1 9108 6290 9108 6290 0 net204
rlabel metal1 41124 31858 41124 31858 0 net205
rlabel metal1 20746 35598 20746 35598 0 net206
rlabel metal1 21896 33626 21896 33626 0 net207
rlabel metal2 17802 19312 17802 19312 0 net208
rlabel metal1 37904 22950 37904 22950 0 net209
rlabel metal2 41354 24582 41354 24582 0 net21
rlabel metal2 28106 32606 28106 32606 0 net210
rlabel metal1 42044 33626 42044 33626 0 net211
rlabel metal1 35466 32538 35466 32538 0 net212
rlabel metal1 27646 16660 27646 16660 0 net213
rlabel metal1 24932 33082 24932 33082 0 net214
rlabel metal1 13754 29614 13754 29614 0 net215
rlabel metal2 38870 10234 38870 10234 0 net216
rlabel metal2 38594 10404 38594 10404 0 net217
rlabel metal1 15134 31314 15134 31314 0 net218
rlabel metal1 41124 14042 41124 14042 0 net219
rlabel metal2 38870 28220 38870 28220 0 net22
rlabel metal1 37904 16082 37904 16082 0 net220
rlabel metal2 36846 7174 36846 7174 0 net221
rlabel metal1 28336 30906 28336 30906 0 net222
rlabel metal2 27738 31314 27738 31314 0 net223
rlabel metal1 24518 34986 24518 34986 0 net224
rlabel metal2 38594 32300 38594 32300 0 net225
rlabel metal1 41170 29070 41170 29070 0 net226
rlabel metal2 36478 7174 36478 7174 0 net227
rlabel metal1 20240 7446 20240 7446 0 net228
rlabel metal1 33994 31314 33994 31314 0 net229
rlabel metal2 40066 23630 40066 23630 0 net23
rlabel metal1 37766 31892 37766 31892 0 net230
rlabel metal1 26174 32470 26174 32470 0 net231
rlabel metal1 22678 10778 22678 10778 0 net232
rlabel metal2 37490 8670 37490 8670 0 net233
rlabel metal1 38870 8568 38870 8568 0 net234
rlabel metal1 28382 6970 28382 6970 0 net235
rlabel metal2 28474 6800 28474 6800 0 net236
rlabel metal2 25162 9180 25162 9180 0 net237
rlabel metal1 26634 8602 26634 8602 0 net238
rlabel metal1 18814 11220 18814 11220 0 net239
rlabel metal1 39698 27472 39698 27472 0 net24
rlabel metal1 19228 21114 19228 21114 0 net240
rlabel metal2 31694 31076 31694 31076 0 net241
rlabel metal1 29946 6290 29946 6290 0 net242
rlabel metal1 25024 7378 25024 7378 0 net243
rlabel metal1 25674 6970 25674 6970 0 net244
rlabel metal1 4048 19346 4048 19346 0 net245
rlabel metal1 13846 35632 13846 35632 0 net246
rlabel metal1 22632 5610 22632 5610 0 net247
rlabel metal1 21804 5882 21804 5882 0 net248
rlabel metal2 16790 33150 16790 33150 0 net249
rlabel metal2 39054 25959 39054 25959 0 net25
rlabel metal1 30958 31450 30958 31450 0 net250
rlabel metal1 19872 8058 19872 8058 0 net251
rlabel metal2 2898 26044 2898 26044 0 net252
rlabel metal1 17940 19754 17940 19754 0 net253
rlabel metal1 29946 8262 29946 8262 0 net254
rlabel metal1 30866 7514 30866 7514 0 net255
rlabel metal1 16790 34034 16790 34034 0 net256
rlabel metal1 26772 31314 26772 31314 0 net257
rlabel metal1 25208 31450 25208 31450 0 net258
rlabel metal1 27876 16490 27876 16490 0 net259
rlabel metal2 41078 26146 41078 26146 0 net26
rlabel metal2 23874 34068 23874 34068 0 net260
rlabel metal2 23966 33762 23966 33762 0 net261
rlabel metal1 13524 31858 13524 31858 0 net262
rlabel metal2 13938 32606 13938 32606 0 net263
rlabel metal1 32982 5882 32982 5882 0 net264
rlabel metal1 21390 22644 21390 22644 0 net265
rlabel metal1 37674 26384 37674 26384 0 net266
rlabel metal1 19964 11730 19964 11730 0 net267
rlabel metal2 19550 11628 19550 11628 0 net268
rlabel metal1 33304 8058 33304 8058 0 net269
rlabel metal2 1426 24956 1426 24956 0 net27
rlabel metal1 12604 29138 12604 29138 0 net270
rlabel metal1 10258 26248 10258 26248 0 net271
rlabel metal1 18032 35802 18032 35802 0 net272
rlabel metal2 39330 12376 39330 12376 0 net273
rlabel metal1 39238 11832 39238 11832 0 net274
rlabel metal1 10074 31246 10074 31246 0 net275
rlabel metal1 35190 6630 35190 6630 0 net276
rlabel metal1 14628 34918 14628 34918 0 net277
rlabel metal1 41262 13906 41262 13906 0 net278
rlabel metal1 29118 17238 29118 17238 0 net279
rlabel metal2 1426 23494 1426 23494 0 net28
rlabel metal1 32062 5338 32062 5338 0 net280
rlabel metal2 19182 34816 19182 34816 0 net281
rlabel metal1 10304 27302 10304 27302 0 net282
rlabel metal1 39560 10030 39560 10030 0 net283
rlabel metal2 8418 5066 8418 5066 0 net284
rlabel metal1 37122 12818 37122 12818 0 net285
rlabel metal1 17710 12274 17710 12274 0 net286
rlabel metal1 40526 15402 40526 15402 0 net287
rlabel metal2 40894 14756 40894 14756 0 net288
rlabel metal1 26036 13838 26036 13838 0 net289
rlabel metal2 1426 22202 1426 22202 0 net29
rlabel metal1 30866 42330 30866 42330 0 net290
rlabel metal1 19596 16558 19596 16558 0 net291
rlabel metal1 40342 31892 40342 31892 0 net292
rlabel metal1 24334 10676 24334 10676 0 net293
rlabel metal2 29762 17374 29762 17374 0 net294
rlabel metal2 35098 13226 35098 13226 0 net295
rlabel metal1 33856 13430 33856 13430 0 net296
rlabel metal2 35282 5372 35282 5372 0 net297
rlabel metal1 33212 21522 33212 21522 0 net298
rlabel metal1 9568 28730 9568 28730 0 net299
rlabel metal1 1702 16626 1702 16626 0 net3
rlabel metal1 1702 28118 1702 28118 0 net30
rlabel metal2 34822 17408 34822 17408 0 net300
rlabel metal1 38456 14790 38456 14790 0 net301
rlabel metal2 13018 30940 13018 30940 0 net302
rlabel metal2 25530 16796 25530 16796 0 net303
rlabel metal2 24426 17000 24426 17000 0 net304
rlabel metal1 32430 17544 32430 17544 0 net305
rlabel metal2 31142 17442 31142 17442 0 net306
rlabel via2 33810 21301 33810 21301 0 net307
rlabel metal1 21574 22508 21574 22508 0 net308
rlabel metal1 15686 35156 15686 35156 0 net309
rlabel metal2 35282 37026 35282 37026 0 net31
rlabel metal1 14904 35734 14904 35734 0 net310
rlabel metal2 17066 40528 17066 40528 0 net311
rlabel metal1 35328 9962 35328 9962 0 net312
rlabel metal2 33902 9758 33902 9758 0 net313
rlabel metal1 8418 22406 8418 22406 0 net314
rlabel metal1 23184 41106 23184 41106 0 net315
rlabel metal1 20378 41786 20378 41786 0 net316
rlabel metal1 3128 12682 3128 12682 0 net317
rlabel metal1 39560 41242 39560 41242 0 net318
rlabel metal1 25622 20366 25622 20366 0 net319
rlabel metal1 20424 38726 20424 38726 0 net32
rlabel metal1 24886 13192 24886 13192 0 net320
rlabel metal2 14214 35428 14214 35428 0 net321
rlabel metal1 30544 35734 30544 35734 0 net322
rlabel metal1 22218 14042 22218 14042 0 net323
rlabel metal2 23782 14178 23782 14178 0 net324
rlabel metal1 25760 42670 25760 42670 0 net325
rlabel metal2 22586 16762 22586 16762 0 net326
rlabel metal2 20930 17850 20930 17850 0 net327
rlabel metal1 33672 42330 33672 42330 0 net328
rlabel metal1 41998 17680 41998 17680 0 net329
rlabel metal1 34730 21624 34730 21624 0 net33
rlabel metal1 40204 18326 40204 18326 0 net330
rlabel metal1 40664 35054 40664 35054 0 net331
rlabel metal1 29118 10642 29118 10642 0 net332
rlabel metal1 29532 9622 29532 9622 0 net333
rlabel metal2 41446 39168 41446 39168 0 net334
rlabel metal1 30268 32470 30268 32470 0 net335
rlabel metal1 40480 17238 40480 17238 0 net336
rlabel metal2 40526 16796 40526 16796 0 net337
rlabel metal1 20700 42670 20700 42670 0 net338
rlabel metal1 25024 37094 25024 37094 0 net339
rlabel metal1 16882 21454 16882 21454 0 net34
rlabel metal1 32752 10642 32752 10642 0 net340
rlabel metal2 31970 10472 31970 10472 0 net341
rlabel metal1 35558 20502 35558 20502 0 net342
rlabel metal1 16698 12172 16698 12172 0 net343
rlabel metal1 17802 20842 17802 20842 0 net344
rlabel metal1 19039 20502 19039 20502 0 net345
rlabel metal1 35650 32742 35650 32742 0 net346
rlabel metal2 19918 36448 19918 36448 0 net347
rlabel metal2 41262 30736 41262 30736 0 net348
rlabel metal2 40158 34850 40158 34850 0 net349
rlabel metal2 10442 35564 10442 35564 0 net35
rlabel metal1 19826 10778 19826 10778 0 net350
rlabel metal1 7636 22066 7636 22066 0 net351
rlabel metal1 34592 12614 34592 12614 0 net352
rlabel metal2 13570 17034 13570 17034 0 net353
rlabel metal1 28244 42194 28244 42194 0 net354
rlabel metal1 25116 21522 25116 21522 0 net355
rlabel metal1 40480 39338 40480 39338 0 net356
rlabel metal1 35236 41514 35236 41514 0 net357
rlabel metal1 30222 30566 30222 30566 0 net358
rlabel metal1 36754 19856 36754 19856 0 net359
rlabel metal1 7774 31416 7774 31416 0 net36
rlabel metal1 37720 41242 37720 41242 0 net360
rlabel metal2 41078 36992 41078 36992 0 net361
rlabel metal1 33488 35666 33488 35666 0 net362
rlabel metal1 8372 14994 8372 14994 0 net363
rlabel metal1 23184 41582 23184 41582 0 net364
rlabel metal1 27554 10778 27554 10778 0 net365
rlabel metal2 31234 20400 31234 20400 0 net366
rlabel metal2 30498 40698 30498 40698 0 net367
rlabel metal2 34362 34782 34362 34782 0 net368
rlabel metal1 14766 33830 14766 33830 0 net369
rlabel metal1 2622 32334 2622 32334 0 net37
rlabel metal1 35282 22032 35282 22032 0 net370
rlabel metal2 27738 13498 27738 13498 0 net371
rlabel metal2 29118 14144 29118 14144 0 net372
rlabel metal1 31050 33558 31050 33558 0 net373
rlabel metal1 36524 21318 36524 21318 0 net374
rlabel metal1 10212 20434 10212 20434 0 net375
rlabel metal1 20700 33626 20700 33626 0 net376
rlabel metal1 26634 42330 26634 42330 0 net377
rlabel metal1 22816 12070 22816 12070 0 net378
rlabel metal1 38318 35666 38318 35666 0 net379
rlabel metal2 8142 32674 8142 32674 0 net38
rlabel metal1 12236 20910 12236 20910 0 net380
rlabel metal1 35558 12070 35558 12070 0 net381
rlabel metal1 23276 11050 23276 11050 0 net382
rlabel metal1 4876 4794 4876 4794 0 net383
rlabel metal2 26082 17238 26082 17238 0 net384
rlabel metal2 23230 36992 23230 36992 0 net385
rlabel metal1 38824 29818 38824 29818 0 net386
rlabel metal1 21574 14348 21574 14348 0 net387
rlabel metal2 36754 11968 36754 11968 0 net388
rlabel metal1 8372 18394 8372 18394 0 net389
rlabel metal2 39882 29308 39882 29308 0 net39
rlabel metal2 21482 17578 21482 17578 0 net390
rlabel metal1 31050 16218 31050 16218 0 net391
rlabel metal1 26358 10710 26358 10710 0 net392
rlabel metal1 28520 20910 28520 20910 0 net393
rlabel metal1 1794 8500 1794 8500 0 net394
rlabel metal1 19596 15130 19596 15130 0 net395
rlabel metal1 30682 11730 30682 11730 0 net396
rlabel metal2 24426 18258 24426 18258 0 net397
rlabel metal2 12650 15164 12650 15164 0 net398
rlabel metal1 35144 14314 35144 14314 0 net399
rlabel metal1 1702 17714 1702 17714 0 net4
rlabel metal1 18722 33456 18722 33456 0 net40
rlabel metal1 25208 12070 25208 12070 0 net400
rlabel metal2 9614 24412 9614 24412 0 net401
rlabel metal1 3174 10642 3174 10642 0 net402
rlabel metal1 6302 5202 6302 5202 0 net403
rlabel metal1 25709 35054 25709 35054 0 net404
rlabel metal2 38870 17374 38870 17374 0 net405
rlabel metal2 35006 17408 35006 17408 0 net406
rlabel metal1 19826 13226 19826 13226 0 net407
rlabel metal1 18630 33082 18630 33082 0 net408
rlabel metal1 33580 12818 33580 12818 0 net409
rlabel metal1 17986 21114 17986 21114 0 net41
rlabel metal2 10166 33354 10166 33354 0 net410
rlabel metal1 10120 15130 10120 15130 0 net411
rlabel metal2 19918 16082 19918 16082 0 net412
rlabel metal1 6026 35734 6026 35734 0 net413
rlabel metal1 16376 37978 16376 37978 0 net414
rlabel metal1 38226 17136 38226 17136 0 net415
rlabel metal2 32614 32096 32614 32096 0 net416
rlabel metal1 11362 12750 11362 12750 0 net417
rlabel metal1 8878 11798 8878 11798 0 net418
rlabel metal1 10258 22746 10258 22746 0 net419
rlabel metal1 19228 21658 19228 21658 0 net42
rlabel metal1 28336 34714 28336 34714 0 net420
rlabel metal1 39836 31790 39836 31790 0 net421
rlabel metal1 36340 33626 36340 33626 0 net422
rlabel metal1 12282 10030 12282 10030 0 net423
rlabel metal1 10074 35734 10074 35734 0 net424
rlabel metal2 5750 6154 5750 6154 0 net425
rlabel metal1 2990 30736 2990 30736 0 net426
rlabel metal1 3358 29206 3358 29206 0 net427
rlabel metal1 12052 8942 12052 8942 0 net428
rlabel metal2 2254 7854 2254 7854 0 net429
rlabel metal1 18170 30566 18170 30566 0 net43
rlabel metal1 18814 37434 18814 37434 0 net430
rlabel metal1 2760 29070 2760 29070 0 net431
rlabel metal1 10028 33966 10028 33966 0 net432
rlabel metal1 8602 32810 8602 32810 0 net433
rlabel metal1 14720 11322 14720 11322 0 net434
rlabel metal2 16054 32266 16054 32266 0 net435
rlabel metal1 22080 37774 22080 37774 0 net436
rlabel metal1 35880 35258 35880 35258 0 net437
rlabel metal2 16790 29852 16790 29852 0 net438
rlabel metal1 32798 36142 32798 36142 0 net439
rlabel metal1 18538 30838 18538 30838 0 net44
rlabel metal2 29394 15555 29394 15555 0 net440
rlabel metal1 13386 12818 13386 12818 0 net441
rlabel metal1 17342 38250 17342 38250 0 net442
rlabel metal1 29716 37842 29716 37842 0 net443
rlabel metal1 36616 37978 36616 37978 0 net444
rlabel metal1 28980 35734 28980 35734 0 net445
rlabel metal1 9338 8534 9338 8534 0 net446
rlabel metal1 23598 38386 23598 38386 0 net447
rlabel metal1 9706 30158 9706 30158 0 net448
rlabel metal1 26450 36754 26450 36754 0 net449
rlabel metal1 35512 27506 35512 27506 0 net45
rlabel metal1 7590 21658 7590 21658 0 net450
rlabel metal2 19274 34612 19274 34612 0 net46
rlabel metal1 21344 35598 21344 35598 0 net47
rlabel metal2 34270 33116 34270 33116 0 net48
rlabel metal2 41998 33762 41998 33762 0 net49
rlabel metal2 41998 6086 41998 6086 0 net5
rlabel metal1 34776 21522 34776 21522 0 net50
rlabel metal2 20654 22236 20654 22236 0 net51
rlabel metal2 20654 32912 20654 32912 0 net52
rlabel metal2 39422 23137 39422 23137 0 net53
rlabel metal2 19918 23358 19918 23358 0 net54
rlabel metal1 27738 24650 27738 24650 0 net55
rlabel metal1 28014 27982 28014 27982 0 net56
rlabel metal1 36294 26996 36294 26996 0 net57
rlabel metal1 13754 10574 13754 10574 0 net58
rlabel metal2 13202 8670 13202 8670 0 net59
rlabel metal1 11592 2414 11592 2414 0 net6
rlabel metal1 20102 30192 20102 30192 0 net60
rlabel metal1 36662 29070 36662 29070 0 net61
rlabel metal1 21436 36210 21436 36210 0 net62
rlabel metal1 34914 41004 34914 41004 0 net63
rlabel metal1 41630 34510 41630 34510 0 net64
rlabel metal2 41906 34238 41906 34238 0 net65
rlabel metal1 18400 24650 18400 24650 0 net66
rlabel viali 33168 24786 33168 24786 0 net67
rlabel metal1 19044 28662 19044 28662 0 net68
rlabel via1 36480 26962 36480 26962 0 net69
rlabel metal1 1702 10574 1702 10574 0 net7
rlabel via1 28200 28050 28200 28050 0 net70
rlabel metal2 19090 28254 19090 28254 0 net71
rlabel metal1 20194 29478 20194 29478 0 net72
rlabel metal1 15318 26894 15318 26894 0 net73
rlabel metal1 29440 25126 29440 25126 0 net74
rlabel metal1 5980 10030 5980 10030 0 net75
rlabel metal1 19596 31858 19596 31858 0 net76
rlabel metal1 32200 25806 32200 25806 0 net77
rlabel metal2 20194 7650 20194 7650 0 net78
rlabel metal1 19918 16558 19918 16558 0 net79
rlabel metal1 1702 13940 1702 13940 0 net8
rlabel metal1 35282 13226 35282 13226 0 net80
rlabel metal1 37490 17034 37490 17034 0 net81
rlabel metal1 7866 20434 7866 20434 0 net82
rlabel metal1 6210 17782 6210 17782 0 net83
rlabel metal1 5750 19788 5750 19788 0 net84
rlabel metal1 20010 38794 20010 38794 0 net85
rlabel metal1 19412 9010 19412 9010 0 net86
rlabel metal1 32246 7854 32246 7854 0 net87
rlabel metal1 19964 8874 19964 8874 0 net88
rlabel metal1 34730 16558 34730 16558 0 net89
rlabel metal1 5152 11662 5152 11662 0 net9
rlabel metal1 35374 15062 35374 15062 0 net90
rlabel metal1 20608 14382 20608 14382 0 net91
rlabel metal2 2714 25330 2714 25330 0 net92
rlabel metal1 14812 27302 14812 27302 0 net93
rlabel metal1 20286 7888 20286 7888 0 net94
rlabel metal2 19550 14858 19550 14858 0 net95
rlabel metal2 38962 10302 38962 10302 0 net96
rlabel metal1 35006 13362 35006 13362 0 net97
rlabel metal1 24978 18904 24978 18904 0 net98
rlabel metal1 19596 11662 19596 11662 0 net99
<< properties >>
string FIXED_BBOX 0 0 43613 45757
<< end >>

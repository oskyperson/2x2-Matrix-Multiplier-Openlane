VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO outel8227
  CLASS BLOCK ;
  FOREIGN outel8227 ;
  ORIGIN 0.000 0.000 ;
  SIZE 187.910 BY 198.630 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 187.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END cs
  PIN dataBusIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 183.910 105.440 187.910 106.040 ;
    END
  END dataBusIn[0]
  PIN dataBusIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 183.910 108.840 187.910 109.440 ;
    END
  END dataBusIn[1]
  PIN dataBusIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 183.910 112.240 187.910 112.840 ;
    END
  END dataBusIn[2]
  PIN dataBusIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 194.630 148.490 198.630 ;
    END
  END dataBusIn[3]
  PIN dataBusIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 194.630 145.270 198.630 ;
    END
  END dataBusIn[4]
  PIN dataBusIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 183.910 81.640 187.910 82.240 ;
    END
  END dataBusIn[5]
  PIN dataBusIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 183.910 122.440 187.910 123.040 ;
    END
  END dataBusIn[6]
  PIN dataBusIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 183.910 119.040 187.910 119.640 ;
    END
  END dataBusIn[7]
  PIN dataBusOut[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END dataBusOut[0]
  PIN dataBusOut[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END dataBusOut[1]
  PIN dataBusOut[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END dataBusOut[2]
  PIN dataBusOut[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END dataBusOut[3]
  PIN dataBusOut[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END dataBusOut[4]
  PIN dataBusOut[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END dataBusOut[5]
  PIN dataBusOut[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END dataBusOut[6]
  PIN dataBusOut[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END dataBusOut[7]
  PIN dataBusSelect
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END dataBusSelect
  PIN gpio[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END gpio[0]
  PIN gpio[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 194.630 116.290 198.630 ;
    END
  END gpio[10]
  PIN gpio[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 194.630 125.950 198.630 ;
    END
  END gpio[11]
  PIN gpio[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 194.630 113.070 198.630 ;
    END
  END gpio[12]
  PIN gpio[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 194.630 119.510 198.630 ;
    END
  END gpio[13]
  PIN gpio[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 194.630 129.170 198.630 ;
    END
  END gpio[14]
  PIN gpio[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 194.630 122.730 198.630 ;
    END
  END gpio[15]
  PIN gpio[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END gpio[16]
  PIN gpio[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gpio[17]
  PIN gpio[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END gpio[18]
  PIN gpio[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END gpio[19]
  PIN gpio[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END gpio[1]
  PIN gpio[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END gpio[20]
  PIN gpio[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.246500 ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 183.910 78.240 187.910 78.840 ;
    END
  END gpio[21]
  PIN gpio[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END gpio[22]
  PIN gpio[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpio[23]
  PIN gpio[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END gpio[24]
  PIN gpio[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END gpio[25]
  PIN gpio[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END gpio[2]
  PIN gpio[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END gpio[3]
  PIN gpio[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END gpio[4]
  PIN gpio[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END gpio[5]
  PIN gpio[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END gpio[6]
  PIN gpio[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END gpio[7]
  PIN gpio[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 194.630 135.610 198.630 ;
    END
  END gpio[8]
  PIN gpio[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 194.630 132.390 198.630 ;
    END
  END gpio[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 183.910 17.040 187.910 17.640 ;
    END
  END nrst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 182.350 187.870 ;
      LAYER li1 ;
        RECT 5.520 10.795 182.160 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.240 182.550 187.920 ;
      LAYER met2 ;
        RECT 6.530 194.350 112.510 194.630 ;
        RECT 113.350 194.350 115.730 194.630 ;
        RECT 116.570 194.350 118.950 194.630 ;
        RECT 119.790 194.350 122.170 194.630 ;
        RECT 123.010 194.350 125.390 194.630 ;
        RECT 126.230 194.350 128.610 194.630 ;
        RECT 129.450 194.350 131.830 194.630 ;
        RECT 132.670 194.350 135.050 194.630 ;
        RECT 135.890 194.350 144.710 194.630 ;
        RECT 145.550 194.350 147.930 194.630 ;
        RECT 148.770 194.350 182.530 194.630 ;
        RECT 6.530 4.280 182.530 194.350 ;
        RECT 6.530 4.000 41.670 4.280 ;
        RECT 42.510 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 99.630 4.280 ;
        RECT 100.470 4.000 102.850 4.280 ;
        RECT 103.690 4.000 106.070 4.280 ;
        RECT 106.910 4.000 109.290 4.280 ;
        RECT 110.130 4.000 112.510 4.280 ;
        RECT 113.350 4.000 182.530 4.280 ;
      LAYER met3 ;
        RECT 4.000 177.840 183.910 187.845 ;
        RECT 4.400 176.440 183.910 177.840 ;
        RECT 4.000 164.240 183.910 176.440 ;
        RECT 4.400 162.840 183.910 164.240 ;
        RECT 4.000 160.840 183.910 162.840 ;
        RECT 4.400 159.440 183.910 160.840 ;
        RECT 4.000 157.440 183.910 159.440 ;
        RECT 4.400 156.040 183.910 157.440 ;
        RECT 4.000 154.040 183.910 156.040 ;
        RECT 4.400 152.640 183.910 154.040 ;
        RECT 4.000 150.640 183.910 152.640 ;
        RECT 4.400 149.240 183.910 150.640 ;
        RECT 4.000 147.240 183.910 149.240 ;
        RECT 4.400 145.840 183.910 147.240 ;
        RECT 4.000 143.840 183.910 145.840 ;
        RECT 4.400 142.440 183.910 143.840 ;
        RECT 4.000 140.440 183.910 142.440 ;
        RECT 4.400 139.040 183.910 140.440 ;
        RECT 4.000 123.440 183.910 139.040 ;
        RECT 4.000 122.040 183.510 123.440 ;
        RECT 4.000 120.040 183.910 122.040 ;
        RECT 4.000 118.640 183.510 120.040 ;
        RECT 4.000 113.240 183.910 118.640 ;
        RECT 4.000 111.840 183.510 113.240 ;
        RECT 4.000 109.840 183.910 111.840 ;
        RECT 4.000 108.440 183.510 109.840 ;
        RECT 4.000 106.440 183.910 108.440 ;
        RECT 4.000 105.040 183.510 106.440 ;
        RECT 4.000 82.640 183.910 105.040 ;
        RECT 4.000 81.240 183.510 82.640 ;
        RECT 4.000 79.240 183.910 81.240 ;
        RECT 4.000 77.840 183.510 79.240 ;
        RECT 4.000 18.040 183.910 77.840 ;
        RECT 4.000 16.640 183.510 18.040 ;
        RECT 4.000 10.715 183.910 16.640 ;
      LAYER met4 ;
        RECT 13.175 15.135 20.640 174.585 ;
        RECT 23.040 15.135 23.940 174.585 ;
        RECT 26.340 15.135 174.240 174.585 ;
        RECT 176.640 15.135 177.265 174.585 ;
  END
END outel8227
END LIBRARY


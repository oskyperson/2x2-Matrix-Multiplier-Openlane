magic
tech sky130A
magscale 1 2
timestamp 1727302560
<< viali >>
rect 20821 37281 20855 37315
rect 23581 37281 23615 37315
rect 17601 37213 17635 37247
rect 23857 37213 23891 37247
rect 29101 37213 29135 37247
rect 29837 37213 29871 37247
rect 17417 37145 17451 37179
rect 20545 37145 20579 37179
rect 21833 37145 21867 37179
rect 17785 37077 17819 37111
rect 20177 37077 20211 37111
rect 20637 37077 20671 37111
rect 29285 37077 29319 37111
rect 29929 37077 29963 37111
rect 15485 36873 15519 36907
rect 15117 36805 15151 36839
rect 17417 36805 17451 36839
rect 21833 36805 21867 36839
rect 14933 36737 14967 36771
rect 15209 36737 15243 36771
rect 15577 36737 15611 36771
rect 15761 36737 15795 36771
rect 15853 36737 15887 36771
rect 16037 36737 16071 36771
rect 16313 36737 16347 36771
rect 16497 36737 16531 36771
rect 16681 36737 16715 36771
rect 16835 36737 16869 36771
rect 17049 36737 17083 36771
rect 17325 36737 17359 36771
rect 17509 36737 17543 36771
rect 17627 36737 17661 36771
rect 18049 36747 18083 36781
rect 18245 36737 18279 36771
rect 18613 36737 18647 36771
rect 18889 36737 18923 36771
rect 19073 36737 19107 36771
rect 23857 36737 23891 36771
rect 9321 36669 9355 36703
rect 11069 36669 11103 36703
rect 11345 36669 11379 36703
rect 12633 36669 12667 36703
rect 12909 36669 12943 36703
rect 14657 36669 14691 36703
rect 14749 36669 14783 36703
rect 15485 36669 15519 36703
rect 15669 36669 15703 36703
rect 16405 36669 16439 36703
rect 17785 36669 17819 36703
rect 18337 36669 18371 36703
rect 18429 36669 18463 36703
rect 19349 36669 19383 36703
rect 19625 36669 19659 36703
rect 21373 36669 21407 36703
rect 23581 36669 23615 36703
rect 15853 36601 15887 36635
rect 18981 36601 19015 36635
rect 15301 36533 15335 36567
rect 17141 36533 17175 36567
rect 18797 36533 18831 36567
rect 13277 36329 13311 36363
rect 16957 36329 16991 36363
rect 19257 36329 19291 36363
rect 22845 36329 22879 36363
rect 24409 36329 24443 36363
rect 25237 36329 25271 36363
rect 9413 36261 9447 36295
rect 10149 36193 10183 36227
rect 13369 36193 13403 36227
rect 13645 36193 13679 36227
rect 14197 36193 14231 36227
rect 16773 36193 16807 36227
rect 18705 36193 18739 36227
rect 18797 36193 18831 36227
rect 18981 36193 19015 36227
rect 19901 36193 19935 36227
rect 20177 36193 20211 36227
rect 21925 36193 21959 36227
rect 22569 36193 22603 36227
rect 23489 36193 23523 36227
rect 25053 36193 25087 36227
rect 25789 36193 25823 36227
rect 7205 36125 7239 36159
rect 7389 36125 7423 36159
rect 9321 36125 9355 36159
rect 9689 36125 9723 36159
rect 9873 36125 9907 36159
rect 12633 36125 12667 36159
rect 12817 36125 12851 36159
rect 12909 36125 12943 36159
rect 13001 36125 13035 36159
rect 13737 36125 13771 36159
rect 14289 36125 14323 36159
rect 19073 36125 19107 36159
rect 19441 36125 19475 36159
rect 19717 36125 19751 36159
rect 22385 36125 22419 36159
rect 23213 36125 23247 36159
rect 24869 36125 24903 36159
rect 9597 36057 9631 36091
rect 10425 36057 10459 36091
rect 12173 36057 12207 36091
rect 14749 36057 14783 36091
rect 16497 36057 16531 36091
rect 18429 36057 18463 36091
rect 24777 36057 24811 36091
rect 25605 36057 25639 36091
rect 7297 35989 7331 36023
rect 9321 35989 9355 36023
rect 9781 35989 9815 36023
rect 14657 35989 14691 36023
rect 18797 35989 18831 36023
rect 19625 35989 19659 36023
rect 22017 35989 22051 36023
rect 22477 35989 22511 36023
rect 23305 35989 23339 36023
rect 25697 35989 25731 36023
rect 10517 35785 10551 35819
rect 11529 35785 11563 35819
rect 11897 35785 11931 35819
rect 12725 35785 12759 35819
rect 14473 35785 14507 35819
rect 14933 35785 14967 35819
rect 15853 35785 15887 35819
rect 18153 35785 18187 35819
rect 21465 35785 21499 35819
rect 24501 35785 24535 35819
rect 17417 35717 17451 35751
rect 18705 35717 18739 35751
rect 22661 35717 22695 35751
rect 24961 35717 24995 35751
rect 6377 35649 6411 35683
rect 8769 35649 8803 35683
rect 8953 35649 8987 35683
rect 9229 35649 9263 35683
rect 9781 35649 9815 35683
rect 9965 35649 9999 35683
rect 10149 35649 10183 35683
rect 10333 35649 10367 35683
rect 10885 35649 10919 35683
rect 12357 35649 12391 35683
rect 12541 35649 12575 35683
rect 12909 35649 12943 35683
rect 13001 35649 13035 35683
rect 13553 35649 13587 35683
rect 14105 35649 14139 35683
rect 14381 35649 14415 35683
rect 14565 35649 14599 35683
rect 14841 35649 14875 35683
rect 15025 35649 15059 35683
rect 15117 35649 15151 35683
rect 15301 35649 15335 35683
rect 15669 35649 15703 35683
rect 16129 35649 16163 35683
rect 16681 35649 16715 35683
rect 16865 35649 16899 35683
rect 16957 35649 16991 35683
rect 17233 35649 17267 35683
rect 17785 35649 17819 35683
rect 18429 35649 18463 35683
rect 20913 35649 20947 35683
rect 21373 35649 21407 35683
rect 24409 35649 24443 35683
rect 24869 35649 24903 35683
rect 6653 35581 6687 35615
rect 9137 35581 9171 35615
rect 9597 35581 9631 35615
rect 10057 35581 10091 35615
rect 10977 35581 11011 35615
rect 11989 35581 12023 35615
rect 12081 35581 12115 35615
rect 13277 35581 13311 35615
rect 13369 35581 13403 35615
rect 13829 35581 13863 35615
rect 15393 35581 15427 35615
rect 15485 35581 15519 35615
rect 16221 35581 16255 35615
rect 17049 35581 17083 35615
rect 17693 35581 17727 35615
rect 20453 35581 20487 35615
rect 21005 35581 21039 35615
rect 21097 35581 21131 35615
rect 22385 35581 22419 35615
rect 25053 35581 25087 35615
rect 8125 35445 8159 35479
rect 8769 35445 8803 35479
rect 11161 35445 11195 35479
rect 13185 35445 13219 35479
rect 13737 35445 13771 35479
rect 13921 35445 13955 35479
rect 14289 35445 14323 35479
rect 16405 35445 16439 35479
rect 20545 35445 20579 35479
rect 6009 35241 6043 35275
rect 6745 35241 6779 35275
rect 7849 35241 7883 35275
rect 8953 35241 8987 35275
rect 9321 35241 9355 35275
rect 10517 35241 10551 35275
rect 11989 35241 12023 35275
rect 13369 35241 13403 35275
rect 15577 35241 15611 35275
rect 17877 35241 17911 35275
rect 7297 35173 7331 35207
rect 8493 35173 8527 35207
rect 11161 35173 11195 35207
rect 13277 35173 13311 35207
rect 13737 35173 13771 35207
rect 16865 35173 16899 35207
rect 7481 35105 7515 35139
rect 9229 35105 9263 35139
rect 10885 35105 10919 35139
rect 11345 35105 11379 35139
rect 13093 35105 13127 35139
rect 15117 35105 15151 35139
rect 15485 35105 15519 35139
rect 17417 35105 17451 35139
rect 18337 35105 18371 35139
rect 21005 35105 21039 35139
rect 23305 35105 23339 35139
rect 5825 35037 5859 35071
rect 6009 35037 6043 35071
rect 6101 35037 6135 35071
rect 6285 35037 6319 35071
rect 6377 35037 6411 35071
rect 6469 35037 6503 35071
rect 7113 35037 7147 35071
rect 7389 35037 7423 35071
rect 7665 35037 7699 35071
rect 7947 35037 7981 35071
rect 8125 35037 8159 35071
rect 8309 35037 8343 35071
rect 8401 35037 8435 35071
rect 8585 35037 8619 35071
rect 8953 35037 8987 35071
rect 9137 35037 9171 35071
rect 9505 35037 9539 35071
rect 10241 35037 10275 35071
rect 10793 35037 10827 35071
rect 11529 35037 11563 35071
rect 11621 35037 11655 35071
rect 12081 35037 12115 35071
rect 12265 35037 12299 35071
rect 12449 35037 12483 35071
rect 13369 35037 13403 35071
rect 13461 35037 13495 35071
rect 13553 35037 13587 35071
rect 14657 35037 14691 35071
rect 14841 35037 14875 35071
rect 14933 35037 14967 35071
rect 15393 35037 15427 35071
rect 15669 35037 15703 35071
rect 15761 35037 15795 35071
rect 16221 35037 16255 35071
rect 16497 35037 16531 35071
rect 17141 35037 17175 35071
rect 17509 35037 17543 35071
rect 19073 35037 19107 35071
rect 20269 35037 20303 35071
rect 23029 35037 23063 35071
rect 27261 35037 27295 35071
rect 27537 35037 27571 35071
rect 8033 34969 8067 35003
rect 9689 34969 9723 35003
rect 10517 34969 10551 35003
rect 13737 34969 13771 35003
rect 16037 34969 16071 35003
rect 19441 34969 19475 35003
rect 20177 34969 20211 35003
rect 21281 34969 21315 35003
rect 24041 34969 24075 35003
rect 25145 34969 25179 35003
rect 25881 34969 25915 35003
rect 6929 34901 6963 34935
rect 8769 34901 8803 34935
rect 10333 34901 10367 34935
rect 14749 34901 14783 34935
rect 15301 34901 15335 34935
rect 16405 34901 16439 34935
rect 27077 34901 27111 34935
rect 27445 34901 27479 34935
rect 6101 34697 6135 34731
rect 6745 34697 6779 34731
rect 7389 34697 7423 34731
rect 9229 34697 9263 34731
rect 9965 34697 9999 34731
rect 12725 34697 12759 34731
rect 12909 34697 12943 34731
rect 15209 34697 15243 34731
rect 16497 34697 16531 34731
rect 16681 34697 16715 34731
rect 17417 34697 17451 34731
rect 18245 34697 18279 34731
rect 22293 34697 22327 34731
rect 25513 34697 25547 34731
rect 7113 34629 7147 34663
rect 7573 34629 7607 34663
rect 8677 34629 8711 34663
rect 13093 34629 13127 34663
rect 19349 34629 19383 34663
rect 19901 34629 19935 34663
rect 21649 34629 21683 34663
rect 22385 34629 22419 34663
rect 24593 34629 24627 34663
rect 6009 34561 6043 34595
rect 6193 34561 6227 34595
rect 6837 34561 6871 34595
rect 7021 34561 7055 34595
rect 7297 34561 7331 34595
rect 7389 34561 7423 34595
rect 7481 34561 7515 34595
rect 7665 34561 7699 34595
rect 7757 34561 7791 34595
rect 7941 34561 7975 34595
rect 8217 34561 8251 34595
rect 8309 34561 8343 34595
rect 8493 34561 8527 34595
rect 9045 34561 9079 34595
rect 9873 34561 9907 34595
rect 10057 34561 10091 34595
rect 12265 34561 12299 34595
rect 12357 34561 12391 34595
rect 12541 34561 12575 34595
rect 12817 34561 12851 34595
rect 15485 34561 15519 34595
rect 17141 34561 17175 34595
rect 17325 34561 17359 34595
rect 17509 34561 17543 34595
rect 17601 34561 17635 34595
rect 17785 34561 17819 34595
rect 18061 34561 18095 34595
rect 18429 34561 18463 34595
rect 19165 34561 19199 34595
rect 19441 34561 19475 34595
rect 25329 34561 25363 34595
rect 26249 34561 26283 34595
rect 26433 34561 26467 34595
rect 27445 34561 27479 34595
rect 8861 34493 8895 34527
rect 15393 34493 15427 34527
rect 15577 34493 15611 34527
rect 15669 34493 15703 34527
rect 16037 34493 16071 34527
rect 16865 34493 16899 34527
rect 16957 34493 16991 34527
rect 17049 34493 17083 34527
rect 19625 34493 19659 34527
rect 22569 34493 22603 34527
rect 22845 34493 22879 34527
rect 26157 34493 26191 34527
rect 27997 34493 28031 34527
rect 29929 34493 29963 34527
rect 6561 34425 6595 34459
rect 16313 34425 16347 34459
rect 7757 34357 7791 34391
rect 13093 34357 13127 34391
rect 19165 34357 19199 34391
rect 28181 34357 28215 34391
rect 29665 34357 29699 34391
rect 7849 34153 7883 34187
rect 9873 34153 9907 34187
rect 11805 34153 11839 34187
rect 12909 34153 12943 34187
rect 13829 34153 13863 34187
rect 14105 34153 14139 34187
rect 15301 34153 15335 34187
rect 16221 34153 16255 34187
rect 23121 34153 23155 34187
rect 7021 34085 7055 34119
rect 8401 34085 8435 34119
rect 10149 34085 10183 34119
rect 14473 34085 14507 34119
rect 14657 34085 14691 34119
rect 15209 34085 15243 34119
rect 16865 34085 16899 34119
rect 17509 34085 17543 34119
rect 18797 34085 18831 34119
rect 6469 34017 6503 34051
rect 7481 34017 7515 34051
rect 8309 34017 8343 34051
rect 9505 34017 9539 34051
rect 10057 34017 10091 34051
rect 11437 34017 11471 34051
rect 13093 34017 13127 34051
rect 13921 34017 13955 34051
rect 15117 34017 15151 34051
rect 15853 34017 15887 34051
rect 16589 34017 16623 34051
rect 17049 34017 17083 34051
rect 18705 34017 18739 34051
rect 19257 34017 19291 34051
rect 23673 34017 23707 34051
rect 24409 34017 24443 34051
rect 26341 34017 26375 34051
rect 28365 34017 28399 34051
rect 4721 33949 4755 33983
rect 6653 33949 6687 33983
rect 6837 33949 6871 33983
rect 6929 33949 6963 33983
rect 7205 33949 7239 33983
rect 7665 33949 7699 33983
rect 8033 33949 8067 33983
rect 8125 33949 8159 33983
rect 8677 33949 8711 33983
rect 9622 33949 9656 33983
rect 10241 33949 10275 33983
rect 10333 33949 10367 33983
rect 10793 33949 10827 33983
rect 10885 33949 10919 33983
rect 10977 33949 11011 33983
rect 11529 33949 11563 33983
rect 12265 33949 12299 33983
rect 12449 33949 12483 33983
rect 12725 33949 12759 33983
rect 13185 33949 13219 33983
rect 13645 33949 13679 33983
rect 13737 33949 13771 33983
rect 14381 33949 14415 33983
rect 14565 33949 14599 33983
rect 14841 33949 14875 33983
rect 15209 33949 15243 33983
rect 15301 33949 15335 33983
rect 15485 33949 15519 33983
rect 15577 33949 15611 33983
rect 16037 33949 16071 33983
rect 16497 33949 16531 33983
rect 17141 33949 17175 33983
rect 17877 33949 17911 33983
rect 18061 33949 18095 33983
rect 18153 33949 18187 33983
rect 18245 33949 18279 33983
rect 18429 33949 18463 33983
rect 18889 33949 18923 33983
rect 18981 33949 19015 33983
rect 21649 33949 21683 33983
rect 22017 33949 22051 33983
rect 22385 33949 22419 33983
rect 23489 33949 23523 33983
rect 23581 33949 23615 33983
rect 24225 33949 24259 33983
rect 24777 33949 24811 33983
rect 30389 33949 30423 33983
rect 32781 33949 32815 33983
rect 4997 33881 5031 33915
rect 8309 33881 8343 33915
rect 8401 33881 8435 33915
rect 11069 33881 11103 33915
rect 14933 33881 14967 33915
rect 18613 33881 18647 33915
rect 19533 33881 19567 33915
rect 21833 33881 21867 33915
rect 21925 33881 21959 33915
rect 26203 33881 26237 33915
rect 26617 33881 26651 33915
rect 29653 33881 29687 33915
rect 6653 33813 6687 33847
rect 7389 33813 7423 33847
rect 8585 33813 8619 33847
rect 11253 33813 11287 33847
rect 13553 33813 13587 33847
rect 15761 33813 15795 33847
rect 21005 33813 21039 33847
rect 22201 33813 22235 33847
rect 24041 33813 24075 33847
rect 28089 33813 28123 33847
rect 29009 33813 29043 33847
rect 29745 33813 29779 33847
rect 30205 33813 30239 33847
rect 32597 33813 32631 33847
rect 5089 33609 5123 33643
rect 6377 33609 6411 33643
rect 7757 33609 7791 33643
rect 11529 33609 11563 33643
rect 16129 33609 16163 33643
rect 18061 33609 18095 33643
rect 21833 33609 21867 33643
rect 29377 33609 29411 33643
rect 33885 33609 33919 33643
rect 5917 33541 5951 33575
rect 6653 33541 6687 33575
rect 10333 33541 10367 33575
rect 11345 33541 11379 33575
rect 13185 33541 13219 33575
rect 16313 33541 16347 33575
rect 16681 33541 16715 33575
rect 18153 33541 18187 33575
rect 19073 33541 19107 33575
rect 24777 33541 24811 33575
rect 27169 33541 27203 33575
rect 5273 33473 5307 33507
rect 5457 33473 5491 33507
rect 5641 33473 5675 33507
rect 5825 33473 5859 33507
rect 6193 33473 6227 33507
rect 6561 33473 6595 33507
rect 6745 33473 6779 33507
rect 6929 33473 6963 33507
rect 7113 33473 7147 33507
rect 7297 33473 7331 33507
rect 7573 33473 7607 33507
rect 7849 33473 7883 33507
rect 10149 33473 10183 33507
rect 10241 33473 10275 33507
rect 10517 33473 10551 33507
rect 11161 33473 11195 33507
rect 11713 33473 11747 33507
rect 11989 33473 12023 33507
rect 12173 33473 12207 33507
rect 12449 33473 12483 33507
rect 13093 33473 13127 33507
rect 13369 33473 13403 33507
rect 13553 33473 13587 33507
rect 13645 33473 13679 33507
rect 13829 33473 13863 33507
rect 14013 33473 14047 33507
rect 14197 33473 14231 33507
rect 14381 33473 14415 33507
rect 14473 33473 14507 33507
rect 14565 33473 14599 33507
rect 14749 33473 14783 33507
rect 14933 33473 14967 33507
rect 15025 33473 15059 33507
rect 15393 33473 15427 33507
rect 15945 33473 15979 33507
rect 16129 33473 16163 33507
rect 16221 33473 16255 33507
rect 16865 33473 16899 33507
rect 18245 33473 18279 33507
rect 18613 33473 18647 33507
rect 18705 33473 18739 33507
rect 18889 33473 18923 33507
rect 19533 33473 19567 33507
rect 19717 33473 19751 33507
rect 20177 33473 20211 33507
rect 23581 33473 23615 33507
rect 24225 33473 24259 33507
rect 26341 33473 26375 33507
rect 27353 33473 27387 33507
rect 27445 33473 27479 33507
rect 29469 33473 29503 33507
rect 31677 33473 31711 33507
rect 32137 33473 32171 33507
rect 5549 33405 5583 33439
rect 8125 33405 8159 33439
rect 9873 33405 9907 33439
rect 10977 33405 11011 33439
rect 12357 33405 12391 33439
rect 12817 33405 12851 33439
rect 13921 33405 13955 33439
rect 15301 33405 15335 33439
rect 17785 33405 17819 33439
rect 18981 33405 19015 33439
rect 19349 33405 19383 33439
rect 19809 33405 19843 33439
rect 23305 33405 23339 33439
rect 24501 33405 24535 33439
rect 26525 33405 26559 33439
rect 27721 33405 27755 33439
rect 29193 33405 29227 33439
rect 29653 33405 29687 33439
rect 31401 33405 31435 33439
rect 32413 33405 32447 33439
rect 6101 33337 6135 33371
rect 9965 33337 9999 33371
rect 15209 33337 15243 33371
rect 15577 33337 15611 33371
rect 6193 33269 6227 33303
rect 15117 33269 15151 33303
rect 21603 33269 21637 33303
rect 23673 33269 23707 33303
rect 26249 33269 26283 33303
rect 26985 33269 27019 33303
rect 4537 33065 4571 33099
rect 5273 33065 5307 33099
rect 5457 33065 5491 33099
rect 6469 33065 6503 33099
rect 6561 33065 6595 33099
rect 7297 33065 7331 33099
rect 7849 33065 7883 33099
rect 9413 33065 9447 33099
rect 12173 33065 12207 33099
rect 19533 33065 19567 33099
rect 24501 33065 24535 33099
rect 25237 33065 25271 33099
rect 31401 33065 31435 33099
rect 32045 33065 32079 33099
rect 3985 32997 4019 33031
rect 4721 32997 4755 33031
rect 5687 32997 5721 33031
rect 9965 32997 9999 33031
rect 24041 32997 24075 33031
rect 27629 32997 27663 33031
rect 28273 32997 28307 33031
rect 29561 32997 29595 33031
rect 4813 32929 4847 32963
rect 4905 32929 4939 32963
rect 5549 32929 5583 32963
rect 6653 32929 6687 32963
rect 22116 32929 22150 32963
rect 22385 32929 22419 32963
rect 25145 32929 25179 32963
rect 25329 32929 25363 32963
rect 29285 32929 29319 32963
rect 31309 32929 31343 32963
rect 32321 32929 32355 32963
rect 33057 32929 33091 32963
rect 4169 32861 4203 32895
rect 4261 32861 4295 32895
rect 5089 32861 5123 32895
rect 5365 32861 5399 32895
rect 5825 32861 5859 32895
rect 6009 32861 6043 32895
rect 6101 32861 6135 32895
rect 6285 32861 6319 32895
rect 6837 32861 6871 32895
rect 7113 32861 7147 32895
rect 7297 32861 7331 32895
rect 7573 32861 7607 32895
rect 8033 32861 8067 32895
rect 8125 32861 8159 32895
rect 8309 32861 8343 32895
rect 8401 32861 8435 32895
rect 9321 32861 9355 32895
rect 9505 32861 9539 32895
rect 10057 32861 10091 32895
rect 10149 32861 10183 32895
rect 10333 32861 10367 32895
rect 11253 32861 11287 32895
rect 11989 32861 12023 32895
rect 14105 32861 14139 32895
rect 19441 32861 19475 32895
rect 20268 32861 20302 32895
rect 20361 32861 20395 32895
rect 21833 32861 21867 32895
rect 24225 32861 24259 32895
rect 24409 32861 24443 32895
rect 24928 32861 24962 32895
rect 25421 32861 25455 32895
rect 25513 32861 25547 32895
rect 25881 32861 25915 32895
rect 27813 32861 27847 32895
rect 27905 32861 27939 32895
rect 27997 32861 28031 32895
rect 28181 32861 28215 32895
rect 28457 32861 28491 32895
rect 28549 32861 28583 32895
rect 28825 32861 28859 32895
rect 29101 32861 29135 32895
rect 31585 32861 31619 32895
rect 31953 32861 31987 32895
rect 32229 32861 32263 32895
rect 32413 32861 32447 32895
rect 32505 32861 32539 32895
rect 3985 32793 4019 32827
rect 4353 32793 4387 32827
rect 4569 32793 4603 32827
rect 6561 32793 6595 32827
rect 9781 32793 9815 32827
rect 11805 32793 11839 32827
rect 14381 32793 14415 32827
rect 16129 32793 16163 32827
rect 19717 32793 19751 32827
rect 19901 32793 19935 32827
rect 22017 32793 22051 32827
rect 28641 32793 28675 32827
rect 28917 32793 28951 32827
rect 31033 32793 31067 32827
rect 31677 32793 31711 32827
rect 31769 32793 31803 32827
rect 32781 32793 32815 32827
rect 7021 32725 7055 32759
rect 10057 32725 10091 32759
rect 10241 32725 10275 32759
rect 11161 32725 11195 32759
rect 19349 32725 19383 32759
rect 19993 32725 20027 32759
rect 21649 32725 21683 32759
rect 23857 32725 23891 32759
rect 24869 32725 24903 32759
rect 25053 32725 25087 32759
rect 27307 32725 27341 32759
rect 4905 32521 4939 32555
rect 6009 32521 6043 32555
rect 6745 32521 6779 32555
rect 6837 32521 6871 32555
rect 18245 32521 18279 32555
rect 19717 32521 19751 32555
rect 19901 32521 19935 32555
rect 21557 32521 21591 32555
rect 22753 32521 22787 32555
rect 23489 32521 23523 32555
rect 25421 32521 25455 32555
rect 27629 32521 27663 32555
rect 27997 32521 28031 32555
rect 29377 32521 29411 32555
rect 30389 32521 30423 32555
rect 30757 32521 30791 32555
rect 31217 32521 31251 32555
rect 31585 32521 31619 32555
rect 31769 32521 31803 32555
rect 33425 32521 33459 32555
rect 1501 32453 1535 32487
rect 6561 32453 6595 32487
rect 7389 32453 7423 32487
rect 9045 32453 9079 32487
rect 10609 32453 10643 32487
rect 10977 32453 11011 32487
rect 16313 32453 16347 32487
rect 22109 32453 22143 32487
rect 22201 32453 22235 32487
rect 23259 32453 23293 32487
rect 24777 32453 24811 32487
rect 27353 32453 27387 32487
rect 28181 32453 28215 32487
rect 29929 32453 29963 32487
rect 30021 32453 30055 32487
rect 31401 32453 31435 32487
rect 32459 32453 32493 32487
rect 32689 32453 32723 32487
rect 3525 32385 3559 32419
rect 4813 32385 4847 32419
rect 4997 32385 5031 32419
rect 5273 32385 5307 32419
rect 5641 32385 5675 32419
rect 6377 32385 6411 32419
rect 7021 32385 7055 32419
rect 7297 32385 7331 32419
rect 7481 32385 7515 32419
rect 7573 32385 7607 32419
rect 7757 32385 7791 32419
rect 7849 32385 7883 32419
rect 8033 32385 8067 32419
rect 8769 32385 8803 32419
rect 11805 32385 11839 32419
rect 12449 32385 12483 32419
rect 15577 32385 15611 32419
rect 15853 32385 15887 32419
rect 16129 32385 16163 32419
rect 16221 32385 16255 32419
rect 16497 32385 16531 32419
rect 17785 32385 17819 32419
rect 18153 32385 18187 32419
rect 18429 32385 18463 32419
rect 18981 32385 19015 32419
rect 19165 32385 19199 32419
rect 19257 32385 19291 32419
rect 19349 32385 19383 32419
rect 19441 32385 19475 32419
rect 19842 32385 19876 32419
rect 20361 32385 20395 32419
rect 21465 32385 21499 32419
rect 21649 32385 21683 32419
rect 21833 32385 21867 32419
rect 21926 32385 21960 32419
rect 22298 32385 22332 32419
rect 22937 32385 22971 32419
rect 23029 32385 23063 32419
rect 23121 32385 23155 32419
rect 23397 32385 23431 32419
rect 24225 32385 24259 32419
rect 24409 32385 24443 32419
rect 25237 32385 25271 32419
rect 26617 32385 26651 32419
rect 27261 32385 27295 32419
rect 28457 32385 28491 32419
rect 29193 32385 29227 32419
rect 29285 32385 29319 32419
rect 29653 32385 29687 32419
rect 29801 32385 29835 32419
rect 30159 32385 30193 32419
rect 31125 32385 31159 32419
rect 31309 32385 31343 32419
rect 31677 32385 31711 32419
rect 32597 32385 32631 32419
rect 32781 32385 32815 32419
rect 32965 32385 32999 32419
rect 33057 32385 33091 32419
rect 33241 32385 33275 32419
rect 3249 32317 3283 32351
rect 5549 32317 5583 32351
rect 5733 32317 5767 32351
rect 7205 32317 7239 32351
rect 12081 32317 12115 32351
rect 17693 32317 17727 32351
rect 17877 32317 17911 32351
rect 17969 32317 18003 32351
rect 24041 32317 24075 32351
rect 25145 32317 25179 32351
rect 26157 32317 26191 32351
rect 26341 32317 26375 32351
rect 26433 32317 26467 32351
rect 26525 32317 26559 32351
rect 26985 32317 27019 32351
rect 27470 32317 27504 32351
rect 28733 32317 28767 32351
rect 30573 32317 30607 32351
rect 30665 32317 30699 32351
rect 30941 32317 30975 32351
rect 31033 32317 31067 32351
rect 32321 32317 32355 32351
rect 12265 32249 12299 32283
rect 15761 32249 15795 32283
rect 18429 32249 18463 32283
rect 19625 32249 19659 32283
rect 28273 32249 28307 32283
rect 29009 32249 29043 32283
rect 30297 32249 30331 32283
rect 5089 32181 5123 32215
rect 5457 32181 5491 32215
rect 5825 32181 5859 32215
rect 7573 32181 7607 32215
rect 7849 32181 7883 32215
rect 10517 32181 10551 32215
rect 11621 32181 11655 32215
rect 11989 32181 12023 32215
rect 15393 32181 15427 32215
rect 15945 32181 15979 32215
rect 17509 32181 17543 32215
rect 20269 32181 20303 32215
rect 22477 32181 22511 32215
rect 24593 32181 24627 32215
rect 25237 32181 25271 32215
rect 25513 32181 25547 32215
rect 26801 32181 26835 32215
rect 27813 32181 27847 32215
rect 27997 32181 28031 32215
rect 28641 32181 28675 32215
rect 29561 32181 29595 32215
rect 31953 32181 31987 32215
rect 2329 31977 2363 32011
rect 3157 31977 3191 32011
rect 6377 31977 6411 32011
rect 7113 31977 7147 32011
rect 8033 31977 8067 32011
rect 9413 31977 9447 32011
rect 13737 31977 13771 32011
rect 17601 31977 17635 32011
rect 21557 31977 21591 32011
rect 22753 31977 22787 32011
rect 24409 31977 24443 32011
rect 27905 31977 27939 32011
rect 29745 31977 29779 32011
rect 30113 31977 30147 32011
rect 30389 31977 30423 32011
rect 31493 31977 31527 32011
rect 32229 31977 32263 32011
rect 32597 31977 32631 32011
rect 5549 31909 5583 31943
rect 6653 31909 6687 31943
rect 9597 31909 9631 31943
rect 9965 31909 9999 31943
rect 10793 31909 10827 31943
rect 15393 31909 15427 31943
rect 15485 31909 15519 31943
rect 21649 31909 21683 31943
rect 22569 31909 22603 31943
rect 24685 31909 24719 31943
rect 29561 31909 29595 31943
rect 30757 31909 30791 31943
rect 32781 31909 32815 31943
rect 3801 31841 3835 31875
rect 6285 31841 6319 31875
rect 7481 31841 7515 31875
rect 7665 31841 7699 31875
rect 8677 31841 8711 31875
rect 10057 31841 10091 31875
rect 13093 31841 13127 31875
rect 13369 31841 13403 31875
rect 24777 31841 24811 31875
rect 26341 31841 26375 31875
rect 27353 31841 27387 31875
rect 28549 31841 28583 31875
rect 31125 31841 31159 31875
rect 2513 31773 2547 31807
rect 2697 31773 2731 31807
rect 2789 31773 2823 31807
rect 3341 31773 3375 31807
rect 3525 31773 3559 31807
rect 3617 31773 3651 31807
rect 5825 31773 5859 31807
rect 5917 31773 5951 31807
rect 6561 31773 6595 31807
rect 6745 31773 6779 31807
rect 6837 31773 6871 31807
rect 7357 31773 7391 31807
rect 7573 31773 7607 31807
rect 7849 31773 7883 31807
rect 8125 31773 8159 31807
rect 8493 31773 8527 31807
rect 9229 31773 9263 31807
rect 9505 31773 9539 31807
rect 9781 31773 9815 31807
rect 10609 31773 10643 31807
rect 10972 31773 11006 31807
rect 11069 31773 11103 31807
rect 11289 31773 11323 31807
rect 11437 31773 11471 31807
rect 13645 31773 13679 31807
rect 15117 31773 15151 31807
rect 15301 31773 15335 31807
rect 15577 31773 15611 31807
rect 15761 31773 15795 31807
rect 17877 31773 17911 31807
rect 19355 31773 19389 31807
rect 19441 31773 19475 31807
rect 19533 31773 19567 31807
rect 19625 31773 19659 31807
rect 19809 31773 19843 31807
rect 19901 31773 19935 31807
rect 19993 31773 20027 31807
rect 22017 31773 22051 31807
rect 22293 31773 22327 31807
rect 22845 31773 22879 31807
rect 23029 31773 23063 31807
rect 23489 31773 23523 31807
rect 24133 31773 24167 31807
rect 24593 31773 24627 31807
rect 24869 31773 24903 31807
rect 25053 31773 25087 31807
rect 25605 31773 25639 31807
rect 25697 31773 25731 31807
rect 25881 31773 25915 31807
rect 25973 31773 26007 31807
rect 26249 31773 26283 31807
rect 26433 31773 26467 31807
rect 26525 31773 26559 31807
rect 26801 31773 26835 31807
rect 26985 31773 27019 31807
rect 27169 31773 27203 31807
rect 27261 31773 27295 31807
rect 27445 31773 27479 31807
rect 27629 31773 27663 31807
rect 28090 31773 28124 31807
rect 28181 31773 28215 31807
rect 28273 31773 28307 31807
rect 30021 31773 30055 31807
rect 30481 31773 30515 31807
rect 30938 31773 30972 31807
rect 31217 31773 31251 31807
rect 32045 31773 32079 31807
rect 32229 31773 32263 31807
rect 29699 31739 29733 31773
rect 4077 31705 4111 31739
rect 9045 31705 9079 31739
rect 11161 31705 11195 31739
rect 17601 31705 17635 31739
rect 22385 31705 22419 31739
rect 22569 31705 22603 31739
rect 23121 31705 23155 31739
rect 23673 31705 23707 31739
rect 28411 31705 28445 31739
rect 29101 31705 29135 31739
rect 29929 31705 29963 31739
rect 31493 31705 31527 31739
rect 32413 31705 32447 31739
rect 5641 31637 5675 31671
rect 8309 31637 8343 31671
rect 10333 31637 10367 31671
rect 11621 31637 11655 31671
rect 17785 31637 17819 31671
rect 20269 31637 20303 31671
rect 24041 31637 24075 31671
rect 25237 31637 25271 31671
rect 25421 31637 25455 31671
rect 26065 31637 26099 31671
rect 28825 31637 28859 31671
rect 31309 31637 31343 31671
rect 32613 31637 32647 31671
rect 4537 31433 4571 31467
rect 6745 31433 6779 31467
rect 6929 31433 6963 31467
rect 9597 31433 9631 31467
rect 9781 31433 9815 31467
rect 10609 31433 10643 31467
rect 11253 31433 11287 31467
rect 19901 31433 19935 31467
rect 25697 31433 25731 31467
rect 26985 31433 27019 31467
rect 30849 31433 30883 31467
rect 31033 31433 31067 31467
rect 32505 31433 32539 31467
rect 33057 31433 33091 31467
rect 2237 31365 2271 31399
rect 2421 31365 2455 31399
rect 4169 31365 4203 31399
rect 7573 31365 7607 31399
rect 15025 31365 15059 31399
rect 21005 31365 21039 31399
rect 24685 31365 24719 31399
rect 25329 31365 25363 31399
rect 25421 31365 25455 31399
rect 25789 31365 25823 31399
rect 25973 31365 26007 31399
rect 27137 31365 27171 31399
rect 27353 31365 27387 31399
rect 31753 31365 31787 31399
rect 31953 31365 31987 31399
rect 32965 31365 32999 31399
rect 2053 31297 2087 31331
rect 2329 31297 2363 31331
rect 4445 31297 4479 31331
rect 4813 31297 4847 31331
rect 4905 31297 4939 31331
rect 4997 31297 5031 31331
rect 5181 31297 5215 31331
rect 5641 31297 5675 31331
rect 6377 31297 6411 31331
rect 6561 31297 6595 31331
rect 7113 31297 7147 31331
rect 7389 31297 7423 31331
rect 8309 31297 8343 31331
rect 8493 31297 8527 31331
rect 8585 31297 8619 31331
rect 8953 31297 8987 31331
rect 9137 31297 9171 31331
rect 9229 31297 9263 31331
rect 9413 31297 9447 31331
rect 9722 31297 9756 31331
rect 10793 31297 10827 31331
rect 10977 31297 11011 31331
rect 11161 31297 11195 31331
rect 11345 31297 11379 31331
rect 11713 31297 11747 31331
rect 12357 31297 12391 31331
rect 14933 31297 14967 31331
rect 15393 31297 15427 31331
rect 17141 31297 17175 31331
rect 18613 31297 18647 31331
rect 18797 31297 18831 31331
rect 18889 31297 18923 31331
rect 19001 31297 19035 31331
rect 20085 31297 20119 31331
rect 20177 31297 20211 31331
rect 20361 31297 20395 31331
rect 20453 31297 20487 31331
rect 20545 31297 20579 31331
rect 20729 31297 20763 31331
rect 20821 31297 20855 31331
rect 20913 31297 20947 31331
rect 21097 31297 21131 31331
rect 21189 31297 21223 31331
rect 21373 31297 21407 31331
rect 22937 31297 22971 31331
rect 25211 31297 25245 31331
rect 25513 31297 25547 31331
rect 26157 31297 26191 31331
rect 26249 31297 26283 31331
rect 27445 31297 27479 31331
rect 27629 31297 27663 31331
rect 27905 31297 27939 31331
rect 28181 31319 28215 31353
rect 28549 31297 28583 31331
rect 28825 31297 28859 31331
rect 29101 31297 29135 31331
rect 29653 31297 29687 31331
rect 29837 31297 29871 31331
rect 30205 31297 30239 31331
rect 30389 31297 30423 31331
rect 30481 31297 30515 31331
rect 32597 31297 32631 31331
rect 32689 31297 32723 31331
rect 33241 31297 33275 31331
rect 5457 31229 5491 31263
rect 5549 31229 5583 31263
rect 7205 31229 7239 31263
rect 9045 31229 9079 31263
rect 10241 31229 10275 31263
rect 11805 31229 11839 31263
rect 12081 31229 12115 31263
rect 12541 31229 12575 31263
rect 13185 31229 13219 31263
rect 14657 31229 14691 31263
rect 16957 31229 16991 31263
rect 18705 31229 18739 31263
rect 23029 31229 23063 31263
rect 24961 31229 24995 31263
rect 25053 31229 25087 31263
rect 26525 31229 26559 31263
rect 30665 31229 30699 31263
rect 7297 31161 7331 31195
rect 7941 31161 7975 31195
rect 8125 31161 8159 31195
rect 8677 31161 8711 31195
rect 9413 31161 9447 31195
rect 21189 31161 21223 31195
rect 26801 31161 26835 31195
rect 27813 31161 27847 31195
rect 28089 31161 28123 31195
rect 28181 31161 28215 31195
rect 30297 31161 30331 31195
rect 31401 31161 31435 31195
rect 31585 31161 31619 31195
rect 32321 31161 32355 31195
rect 1869 31093 1903 31127
rect 6009 31093 6043 31127
rect 8033 31093 8067 31127
rect 8493 31093 8527 31127
rect 10149 31093 10183 31127
rect 12173 31093 12207 31127
rect 17325 31093 17359 31127
rect 20545 31093 20579 31127
rect 23213 31093 23247 31127
rect 26341 31093 26375 31127
rect 27209 31093 27243 31127
rect 27537 31093 27571 31127
rect 28917 31093 28951 31127
rect 31033 31093 31067 31127
rect 31809 31093 31843 31127
rect 32873 31093 32907 31127
rect 33425 31093 33459 31127
rect 4537 30889 4571 30923
rect 4813 30889 4847 30923
rect 5273 30889 5307 30923
rect 6837 30889 6871 30923
rect 7481 30889 7515 30923
rect 8401 30889 8435 30923
rect 11713 30889 11747 30923
rect 18061 30889 18095 30923
rect 21373 30889 21407 30923
rect 24593 30889 24627 30923
rect 27445 30889 27479 30923
rect 27721 30889 27755 30923
rect 30757 30889 30791 30923
rect 31217 30889 31251 30923
rect 6377 30821 6411 30855
rect 9781 30821 9815 30855
rect 10149 30821 10183 30855
rect 10977 30821 11011 30855
rect 14841 30821 14875 30855
rect 16497 30821 16531 30855
rect 19349 30821 19383 30855
rect 21189 30821 21223 30855
rect 23213 30821 23247 30855
rect 26893 30821 26927 30855
rect 28181 30821 28215 30855
rect 1501 30753 1535 30787
rect 6193 30753 6227 30787
rect 8033 30753 8067 30787
rect 9505 30753 9539 30787
rect 10701 30753 10735 30787
rect 11437 30753 11471 30787
rect 13829 30753 13863 30787
rect 3801 30685 3835 30719
rect 3985 30685 4019 30719
rect 4169 30685 4203 30719
rect 4261 30685 4295 30719
rect 4353 30685 4387 30719
rect 4537 30685 4571 30719
rect 6653 30685 6687 30719
rect 6745 30685 6779 30719
rect 6929 30685 6963 30719
rect 7113 30685 7147 30719
rect 7297 30685 7331 30719
rect 7573 30685 7607 30719
rect 7941 30685 7975 30719
rect 8125 30685 8159 30719
rect 8217 30685 8251 30719
rect 8401 30685 8435 30719
rect 9413 30685 9447 30719
rect 11345 30685 11379 30719
rect 11805 30685 11839 30719
rect 13553 30685 13587 30719
rect 14289 30685 14323 30719
rect 15853 30685 15887 30719
rect 15946 30685 15980 30719
rect 16129 30685 16163 30719
rect 16318 30685 16352 30719
rect 16589 30685 16623 30719
rect 16681 30685 16715 30719
rect 16865 30685 16899 30719
rect 16957 30685 16991 30719
rect 18981 30685 19015 30719
rect 19533 30685 19567 30719
rect 19625 30685 19659 30719
rect 19809 30685 19843 30719
rect 19901 30685 19935 30719
rect 21741 30685 21775 30719
rect 22017 30685 22051 30719
rect 22201 30685 22235 30719
rect 22477 30685 22511 30719
rect 22753 30685 22787 30719
rect 22845 30685 22879 30719
rect 23397 30685 23431 30719
rect 23581 30685 23615 30719
rect 23857 30685 23891 30719
rect 24409 30685 24443 30719
rect 24593 30685 24627 30719
rect 26617 30685 26651 30719
rect 27077 30685 27111 30719
rect 27261 30685 27295 30719
rect 27629 30685 27663 30719
rect 27813 30685 27847 30719
rect 27905 30685 27939 30719
rect 28089 30685 28123 30719
rect 28181 30685 28215 30719
rect 28365 30685 28399 30719
rect 28917 30685 28951 30719
rect 29101 30685 29135 30719
rect 29929 30685 29963 30719
rect 31125 30685 31159 30719
rect 31309 30685 31343 30719
rect 1777 30617 1811 30651
rect 3525 30617 3559 30651
rect 4997 30617 5031 30651
rect 5457 30617 5491 30651
rect 5917 30617 5951 30651
rect 6377 30617 6411 30651
rect 14105 30617 14139 30651
rect 14657 30617 14691 30651
rect 16221 30617 16255 30651
rect 17693 30617 17727 30651
rect 17877 30617 17911 30651
rect 24041 30617 24075 30651
rect 24225 30617 24259 30651
rect 26341 30617 26375 30651
rect 27537 30617 27571 30651
rect 28641 30617 28675 30651
rect 29745 30617 29779 30651
rect 30573 30617 30607 30651
rect 30757 30617 30791 30651
rect 4629 30549 4663 30583
rect 4797 30549 4831 30583
rect 5089 30549 5123 30583
rect 5257 30549 5291 30583
rect 5549 30549 5583 30583
rect 6009 30549 6043 30583
rect 6561 30549 6595 30583
rect 7757 30549 7791 30583
rect 10517 30549 10551 30583
rect 10609 30549 10643 30583
rect 13185 30549 13219 30583
rect 13645 30549 13679 30583
rect 14473 30549 14507 30583
rect 17141 30549 17175 30583
rect 18889 30549 18923 30583
rect 21373 30549 21407 30583
rect 23489 30549 23523 30583
rect 24869 30549 24903 30583
rect 27997 30549 28031 30583
rect 29561 30549 29595 30583
rect 30941 30549 30975 30583
rect 6101 30345 6135 30379
rect 10717 30345 10751 30379
rect 10885 30345 10919 30379
rect 11621 30345 11655 30379
rect 14105 30345 14139 30379
rect 22201 30345 22235 30379
rect 9137 30277 9171 30311
rect 10057 30277 10091 30311
rect 10517 30277 10551 30311
rect 18061 30277 18095 30311
rect 19165 30277 19199 30311
rect 27629 30277 27663 30311
rect 28181 30277 28215 30311
rect 28825 30277 28859 30311
rect 3617 30209 3651 30243
rect 3709 30209 3743 30243
rect 5733 30209 5767 30243
rect 7757 30209 7791 30243
rect 8861 30209 8895 30243
rect 9229 30209 9263 30243
rect 10149 30209 10183 30243
rect 11253 30209 11287 30243
rect 11529 30209 11563 30243
rect 11713 30209 11747 30243
rect 11805 30209 11839 30243
rect 13277 30209 13311 30243
rect 14013 30209 14047 30243
rect 14197 30209 14231 30243
rect 14841 30209 14875 30243
rect 14933 30209 14967 30243
rect 17877 30209 17911 30243
rect 18153 30209 18187 30243
rect 18521 30209 18555 30243
rect 18797 30209 18831 30243
rect 18889 30209 18923 30243
rect 19073 30209 19107 30243
rect 19257 30209 19291 30243
rect 19717 30209 19751 30243
rect 22017 30209 22051 30243
rect 22569 30209 22603 30243
rect 22661 30209 22695 30243
rect 22753 30209 22787 30243
rect 22871 30209 22905 30243
rect 23305 30209 23339 30243
rect 23489 30209 23523 30243
rect 23581 30209 23615 30243
rect 23765 30209 23799 30243
rect 26341 30209 26375 30243
rect 26433 30209 26467 30243
rect 26525 30209 26559 30243
rect 26709 30209 26743 30243
rect 27169 30209 27203 30243
rect 27261 30209 27295 30243
rect 27721 30209 27755 30243
rect 27905 30209 27939 30243
rect 28733 30209 28767 30243
rect 28917 30209 28951 30243
rect 29009 30209 29043 30243
rect 29561 30209 29595 30243
rect 29837 30209 29871 30243
rect 30297 30209 30331 30243
rect 30665 30209 30699 30243
rect 30849 30209 30883 30243
rect 33057 30209 33091 30243
rect 33150 30209 33184 30243
rect 33333 30209 33367 30243
rect 33425 30209 33459 30243
rect 33522 30209 33556 30243
rect 34253 30209 34287 30243
rect 34437 30209 34471 30243
rect 28641 30175 28675 30209
rect 1593 30141 1627 30175
rect 3341 30141 3375 30175
rect 3985 30141 4019 30175
rect 5825 30141 5859 30175
rect 7481 30141 7515 30175
rect 7665 30141 7699 30175
rect 8677 30141 8711 30175
rect 9781 30141 9815 30175
rect 10266 30141 10300 30175
rect 13185 30141 13219 30175
rect 17693 30141 17727 30175
rect 18337 30141 18371 30175
rect 19349 30141 19383 30175
rect 19441 30141 19475 30175
rect 23029 30141 23063 30175
rect 23949 30141 23983 30175
rect 24041 30141 24075 30175
rect 25789 30141 25823 30175
rect 26065 30141 26099 30175
rect 27537 30141 27571 30175
rect 28365 30141 28399 30175
rect 28549 30141 28583 30175
rect 29469 30141 29503 30175
rect 10425 30073 10459 30107
rect 13645 30073 13679 30107
rect 14565 30073 14599 30107
rect 18245 30073 18279 30107
rect 26157 30073 26191 30107
rect 30481 30073 30515 30107
rect 34069 30073 34103 30107
rect 5457 30005 5491 30039
rect 8125 30005 8159 30039
rect 10701 30005 10735 30039
rect 11069 30005 11103 30039
rect 11897 30005 11931 30039
rect 14933 30005 14967 30039
rect 19533 30005 19567 30039
rect 19625 30005 19659 30039
rect 22385 30005 22419 30039
rect 23121 30005 23155 30039
rect 26985 30005 27019 30039
rect 27721 30005 27755 30039
rect 29929 30005 29963 30039
rect 33701 30005 33735 30039
rect 3801 29801 3835 29835
rect 4813 29801 4847 29835
rect 10701 29801 10735 29835
rect 18429 29801 18463 29835
rect 18613 29801 18647 29835
rect 19257 29801 19291 29835
rect 26893 29801 26927 29835
rect 28181 29801 28215 29835
rect 11897 29733 11931 29767
rect 22109 29733 22143 29767
rect 22201 29733 22235 29767
rect 25421 29733 25455 29767
rect 25973 29733 26007 29767
rect 27905 29733 27939 29767
rect 1501 29665 1535 29699
rect 3249 29665 3283 29699
rect 3525 29665 3559 29699
rect 4261 29665 4295 29699
rect 4353 29665 4387 29699
rect 5457 29665 5491 29699
rect 9597 29665 9631 29699
rect 12173 29665 12207 29699
rect 13461 29665 13495 29699
rect 14105 29665 14139 29699
rect 15301 29665 15335 29699
rect 15853 29665 15887 29699
rect 16589 29665 16623 29699
rect 19533 29665 19567 29699
rect 19625 29665 19659 29699
rect 27537 29665 27571 29699
rect 31769 29665 31803 29699
rect 32045 29665 32079 29699
rect 5273 29597 5307 29631
rect 5641 29597 5675 29631
rect 7389 29597 7423 29631
rect 7757 29597 7791 29631
rect 8125 29597 8159 29631
rect 8309 29597 8343 29631
rect 10241 29597 10275 29631
rect 10517 29597 10551 29631
rect 10701 29597 10735 29631
rect 11805 29597 11839 29631
rect 12265 29597 12299 29631
rect 12633 29597 12667 29631
rect 12817 29597 12851 29631
rect 12909 29597 12943 29631
rect 13369 29597 13403 29631
rect 13737 29597 13771 29631
rect 13829 29597 13863 29631
rect 14381 29597 14415 29631
rect 14478 29597 14512 29631
rect 15669 29597 15703 29631
rect 16129 29597 16163 29631
rect 16957 29597 16991 29631
rect 17141 29597 17175 29631
rect 18153 29597 18187 29631
rect 18521 29597 18555 29631
rect 18889 29597 18923 29631
rect 19441 29597 19475 29631
rect 19717 29597 19751 29631
rect 20637 29597 20671 29631
rect 20821 29597 20855 29631
rect 20913 29597 20947 29631
rect 21005 29597 21039 29631
rect 21189 29597 21223 29631
rect 21649 29597 21683 29631
rect 22661 29597 22695 29631
rect 22845 29597 22879 29631
rect 23305 29597 23339 29631
rect 23765 29597 23799 29631
rect 25605 29597 25639 29631
rect 25789 29597 25823 29631
rect 26433 29597 26467 29631
rect 26893 29597 26927 29631
rect 27077 29597 27111 29631
rect 27169 29597 27203 29631
rect 28089 29597 28123 29631
rect 28273 29597 28307 29631
rect 31217 29597 31251 29631
rect 31401 29597 31435 29631
rect 31677 29597 31711 29631
rect 32137 29597 32171 29631
rect 4169 29529 4203 29563
rect 13001 29529 13035 29563
rect 14105 29529 14139 29563
rect 14289 29529 14323 29563
rect 16221 29529 16255 29563
rect 16313 29529 16347 29563
rect 16451 29529 16485 29563
rect 24593 29529 24627 29563
rect 25053 29529 25087 29563
rect 25237 29529 25271 29563
rect 26617 29529 26651 29563
rect 5181 29461 5215 29495
rect 5733 29461 5767 29495
rect 8953 29461 8987 29495
rect 9321 29461 9355 29495
rect 9413 29461 9447 29495
rect 10333 29461 10367 29495
rect 15669 29461 15703 29495
rect 15945 29461 15979 29495
rect 16773 29461 16807 29495
rect 18245 29461 18279 29495
rect 21373 29461 21407 29495
rect 21741 29461 21775 29495
rect 24869 29461 24903 29495
rect 26249 29461 26283 29495
rect 26709 29461 26743 29495
rect 27997 29461 28031 29495
rect 31585 29461 31619 29495
rect 31861 29461 31895 29495
rect 32321 29461 32355 29495
rect 4353 29257 4387 29291
rect 13277 29257 13311 29291
rect 18797 29257 18831 29291
rect 20177 29257 20211 29291
rect 22661 29257 22695 29291
rect 25559 29257 25593 29291
rect 29469 29257 29503 29291
rect 1777 29189 1811 29223
rect 4261 29189 4295 29223
rect 7113 29189 7147 29223
rect 7941 29189 7975 29223
rect 10241 29189 10275 29223
rect 20913 29189 20947 29223
rect 22293 29189 22327 29223
rect 30389 29189 30423 29223
rect 30757 29189 30791 29223
rect 17325 29155 17359 29189
rect 3801 29121 3835 29155
rect 6837 29121 6871 29155
rect 6929 29121 6963 29155
rect 7205 29121 7239 29155
rect 7370 29121 7404 29155
rect 7757 29121 7791 29155
rect 9597 29121 9631 29155
rect 9965 29121 9999 29155
rect 12081 29121 12115 29155
rect 12541 29121 12575 29155
rect 12909 29121 12943 29155
rect 13093 29121 13127 29155
rect 13645 29121 13679 29155
rect 14013 29121 14047 29155
rect 14473 29121 14507 29155
rect 15117 29121 15151 29155
rect 16865 29121 16899 29155
rect 17141 29121 17175 29155
rect 17601 29121 17635 29155
rect 17877 29121 17911 29155
rect 18429 29121 18463 29155
rect 18521 29121 18555 29155
rect 18613 29121 18647 29155
rect 20453 29121 20487 29155
rect 20545 29121 20579 29155
rect 20637 29121 20671 29155
rect 20821 29121 20855 29155
rect 21097 29121 21131 29155
rect 21189 29121 21223 29155
rect 21465 29121 21499 29155
rect 22017 29121 22051 29155
rect 22569 29121 22603 29155
rect 22845 29121 22879 29155
rect 23213 29121 23247 29155
rect 23765 29121 23799 29155
rect 26525 29121 26559 29155
rect 27537 29121 27571 29155
rect 28273 29121 28307 29155
rect 28549 29121 28583 29155
rect 28733 29121 28767 29155
rect 28917 29121 28951 29155
rect 29377 29121 29411 29155
rect 29561 29121 29595 29155
rect 29837 29121 29871 29155
rect 29929 29121 29963 29155
rect 30665 29121 30699 29155
rect 31217 29121 31251 29155
rect 31585 29121 31619 29155
rect 35817 29121 35851 29155
rect 3525 29053 3559 29087
rect 4445 29053 4479 29087
rect 7481 29053 7515 29087
rect 7573 29053 7607 29087
rect 9321 29053 9355 29087
rect 12633 29053 12667 29087
rect 13185 29053 13219 29087
rect 13461 29053 13495 29087
rect 13921 29053 13955 29087
rect 14749 29053 14783 29087
rect 15301 29053 15335 29087
rect 15577 29053 15611 29087
rect 15669 29053 15703 29087
rect 16037 29053 16071 29087
rect 17049 29053 17083 29087
rect 22201 29053 22235 29087
rect 24133 29053 24167 29087
rect 26249 29053 26283 29087
rect 27077 29053 27111 29087
rect 27169 29053 27203 29087
rect 30849 29053 30883 29087
rect 34713 29053 34747 29087
rect 34989 29053 35023 29087
rect 3893 28985 3927 29019
rect 12173 28985 12207 29019
rect 14289 28985 14323 29019
rect 14933 28985 14967 29019
rect 15393 28985 15427 29019
rect 16957 28985 16991 29019
rect 17417 28985 17451 29019
rect 17785 28985 17819 29019
rect 18245 28985 18279 29019
rect 21373 28985 21407 29019
rect 23581 28985 23615 29019
rect 28365 28985 28399 29019
rect 28457 28985 28491 29019
rect 30021 28985 30055 29019
rect 35633 28985 35667 29019
rect 14657 28917 14691 28951
rect 16681 28917 16715 28951
rect 21833 28917 21867 28951
rect 22017 28917 22051 28951
rect 28089 28917 28123 28951
rect 28733 28917 28767 28951
rect 31033 28917 31067 28951
rect 7941 28713 7975 28747
rect 8309 28713 8343 28747
rect 9505 28713 9539 28747
rect 15761 28713 15795 28747
rect 20821 28713 20855 28747
rect 21557 28713 21591 28747
rect 22293 28713 22327 28747
rect 25881 28713 25915 28747
rect 27629 28713 27663 28747
rect 28273 28713 28307 28747
rect 28457 28713 28491 28747
rect 34161 28713 34195 28747
rect 35357 28713 35391 28747
rect 5549 28645 5583 28679
rect 6285 28645 6319 28679
rect 8125 28645 8159 28679
rect 14105 28645 14139 28679
rect 16589 28645 16623 28679
rect 21695 28645 21729 28679
rect 22385 28645 22419 28679
rect 34345 28645 34379 28679
rect 1593 28577 1627 28611
rect 3617 28577 3651 28611
rect 4997 28577 5031 28611
rect 7573 28577 7607 28611
rect 7849 28577 7883 28611
rect 7941 28577 7975 28611
rect 9965 28577 9999 28611
rect 12909 28577 12943 28611
rect 20177 28577 20211 28611
rect 22477 28577 22511 28611
rect 22753 28577 22787 28611
rect 23397 28577 23431 28611
rect 27795 28577 27829 28611
rect 28549 28577 28583 28611
rect 28825 28577 28859 28611
rect 32229 28577 32263 28611
rect 34713 28577 34747 28611
rect 3985 28509 4019 28543
rect 4261 28509 4295 28543
rect 5641 28509 5675 28543
rect 5733 28509 5767 28543
rect 6043 28509 6077 28543
rect 6469 28509 6503 28543
rect 6561 28509 6595 28543
rect 7297 28509 7331 28543
rect 7389 28509 7423 28543
rect 7665 28509 7699 28543
rect 7757 28509 7791 28543
rect 8217 28509 8251 28543
rect 8493 28509 8527 28543
rect 8585 28509 8619 28543
rect 9229 28509 9263 28543
rect 9413 28509 9447 28543
rect 9689 28509 9723 28543
rect 9781 28509 9815 28543
rect 10057 28509 10091 28543
rect 10333 28509 10367 28543
rect 10425 28509 10459 28543
rect 10885 28509 10919 28543
rect 11069 28509 11103 28543
rect 12081 28509 12115 28543
rect 12357 28509 12391 28543
rect 13001 28509 13035 28543
rect 13369 28509 13403 28543
rect 13737 28509 13771 28543
rect 14565 28509 14599 28543
rect 14841 28509 14875 28543
rect 15209 28509 15243 28543
rect 15301 28509 15335 28543
rect 15393 28509 15427 28543
rect 15577 28509 15611 28543
rect 15945 28509 15979 28543
rect 16037 28509 16071 28543
rect 16221 28509 16255 28543
rect 16313 28509 16347 28543
rect 16405 28509 16439 28543
rect 16589 28509 16623 28543
rect 18797 28509 18831 28543
rect 18981 28509 19015 28543
rect 20545 28509 20579 28543
rect 20913 28509 20947 28543
rect 21097 28509 21131 28543
rect 21373 28509 21407 28543
rect 21833 28509 21867 28543
rect 22017 28509 22051 28543
rect 23213 28509 23247 28543
rect 24041 28509 24075 28543
rect 24409 28509 24443 28543
rect 24961 28509 24995 28543
rect 25237 28509 25271 28543
rect 26065 28509 26099 28543
rect 26249 28509 26283 28543
rect 26433 28509 26467 28543
rect 26525 28509 26559 28543
rect 26617 28509 26651 28543
rect 27077 28509 27111 28543
rect 27445 28509 27479 28543
rect 27905 28509 27939 28543
rect 28273 28509 28307 28543
rect 31769 28509 31803 28543
rect 32071 28509 32105 28543
rect 33793 28509 33827 28543
rect 35081 28509 35115 28543
rect 35173 28509 35207 28543
rect 3341 28441 3375 28475
rect 3801 28441 3835 28475
rect 5181 28441 5215 28475
rect 10149 28441 10183 28475
rect 11621 28441 11655 28475
rect 14289 28441 14323 28475
rect 14473 28441 14507 28475
rect 14933 28441 14967 28475
rect 15485 28441 15519 28475
rect 20453 28441 20487 28475
rect 20662 28441 20696 28475
rect 26157 28441 26191 28475
rect 27261 28441 27295 28475
rect 27353 28441 27387 28475
rect 31861 28441 31895 28475
rect 31953 28441 31987 28475
rect 34851 28441 34885 28475
rect 34989 28441 35023 28475
rect 4169 28373 4203 28407
rect 5089 28373 5123 28407
rect 6745 28373 6779 28407
rect 7113 28373 7147 28407
rect 8769 28373 8803 28407
rect 9321 28373 9355 28407
rect 10793 28373 10827 28407
rect 10977 28373 11011 28407
rect 11713 28373 11747 28407
rect 15025 28373 15059 28407
rect 18889 28373 18923 28407
rect 21005 28373 21039 28407
rect 21373 28373 21407 28407
rect 22661 28373 22695 28407
rect 23791 28373 23825 28407
rect 24593 28373 24627 28407
rect 26801 28373 26835 28407
rect 31585 28373 31619 28407
rect 34170 28373 34204 28407
rect 4353 28169 4387 28203
rect 7389 28169 7423 28203
rect 9229 28169 9263 28203
rect 13185 28169 13219 28203
rect 21005 28169 21039 28203
rect 25145 28169 25179 28203
rect 25513 28169 25547 28203
rect 25973 28169 26007 28203
rect 27169 28169 27203 28203
rect 27629 28169 27663 28203
rect 28825 28169 28859 28203
rect 6929 28101 6963 28135
rect 7113 28101 7147 28135
rect 7481 28101 7515 28135
rect 21189 28101 21223 28135
rect 22201 28101 22235 28135
rect 25605 28101 25639 28135
rect 26433 28101 26467 28135
rect 26985 28101 27019 28135
rect 29791 28101 29825 28135
rect 30021 28101 30055 28135
rect 31585 28101 31619 28135
rect 32597 28101 32631 28135
rect 3433 28033 3467 28067
rect 4350 28033 4384 28067
rect 4813 28033 4847 28067
rect 5825 28033 5859 28067
rect 6101 28033 6135 28067
rect 7389 28033 7423 28067
rect 7665 28033 7699 28067
rect 8308 28033 8342 28067
rect 8585 28033 8619 28067
rect 8769 28033 8803 28067
rect 8861 28033 8895 28067
rect 9137 28033 9171 28067
rect 9229 28033 9263 28067
rect 9413 28033 9447 28067
rect 9965 28033 9999 28067
rect 10057 28033 10091 28067
rect 10149 28033 10183 28067
rect 10241 28033 10275 28067
rect 10517 28033 10551 28067
rect 10609 28033 10643 28067
rect 11069 28033 11103 28067
rect 11253 28033 11287 28067
rect 11897 28033 11931 28067
rect 12357 28033 12391 28067
rect 12449 28033 12483 28067
rect 13369 28033 13403 28067
rect 13553 28033 13587 28067
rect 14105 28033 14139 28067
rect 14749 28033 14783 28067
rect 15485 28033 15519 28067
rect 16129 28033 16163 28067
rect 17141 28033 17175 28067
rect 17325 28033 17359 28067
rect 18521 28033 18555 28067
rect 18797 28033 18831 28067
rect 18981 28033 19015 28067
rect 19717 28033 19751 28067
rect 20729 28033 20763 28067
rect 22017 28033 22051 28067
rect 22293 28033 22327 28067
rect 22385 28033 22419 28067
rect 22937 28033 22971 28067
rect 23121 28033 23155 28067
rect 23397 28033 23431 28067
rect 27537 28033 27571 28067
rect 27721 28033 27755 28067
rect 28457 28033 28491 28067
rect 29653 28033 29687 28067
rect 29929 28033 29963 28067
rect 30113 28033 30147 28067
rect 30573 28033 30607 28067
rect 30665 28033 30699 28067
rect 30757 28033 30791 28067
rect 31493 28033 31527 28067
rect 31769 28033 31803 28067
rect 32413 28033 32447 28067
rect 32689 28033 32723 28067
rect 32781 28033 32815 28067
rect 1409 27965 1443 27999
rect 3157 27965 3191 27999
rect 4721 27965 4755 27999
rect 4951 27965 4985 27999
rect 7205 27965 7239 27999
rect 7849 27965 7883 27999
rect 7941 27965 7975 27999
rect 8493 27965 8527 27999
rect 10977 27965 11011 27999
rect 11161 27965 11195 27999
rect 12081 27965 12115 27999
rect 14933 27965 14967 27999
rect 16773 27965 16807 27999
rect 19073 27965 19107 27999
rect 19533 27965 19567 27999
rect 22845 27965 22879 27999
rect 23029 27965 23063 27999
rect 23673 27965 23707 27999
rect 25421 27965 25455 27999
rect 28733 27965 28767 27999
rect 28942 27965 28976 27999
rect 30389 27965 30423 27999
rect 30849 27965 30883 27999
rect 5365 27897 5399 27931
rect 11529 27897 11563 27931
rect 19165 27897 19199 27931
rect 19901 27897 19935 27931
rect 26065 27897 26099 27931
rect 30297 27897 30331 27931
rect 4169 27829 4203 27863
rect 6653 27829 6687 27863
rect 9045 27829 9079 27863
rect 9781 27829 9815 27863
rect 10793 27829 10827 27863
rect 18337 27829 18371 27863
rect 21005 27829 21039 27863
rect 22569 27829 22603 27863
rect 22661 27829 22695 27863
rect 26433 27829 26467 27863
rect 26617 27829 26651 27863
rect 27169 27829 27203 27863
rect 27353 27829 27387 27863
rect 29101 27829 29135 27863
rect 31953 27829 31987 27863
rect 32965 27829 32999 27863
rect 4721 27625 4755 27659
rect 4905 27625 4939 27659
rect 6285 27625 6319 27659
rect 7389 27625 7423 27659
rect 10333 27625 10367 27659
rect 11529 27625 11563 27659
rect 15412 27625 15446 27659
rect 23397 27625 23431 27659
rect 26065 27625 26099 27659
rect 26617 27625 26651 27659
rect 26893 27625 26927 27659
rect 30757 27625 30791 27659
rect 31677 27625 31711 27659
rect 2237 27557 2271 27591
rect 12265 27557 12299 27591
rect 13645 27557 13679 27591
rect 15301 27557 15335 27591
rect 17141 27557 17175 27591
rect 31401 27557 31435 27591
rect 4537 27489 4571 27523
rect 5457 27489 5491 27523
rect 7573 27489 7607 27523
rect 8769 27489 8803 27523
rect 9321 27489 9355 27523
rect 11621 27489 11655 27523
rect 13277 27489 13311 27523
rect 14841 27489 14875 27523
rect 15209 27489 15243 27523
rect 19533 27489 19567 27523
rect 25145 27489 25179 27523
rect 26249 27489 26283 27523
rect 29837 27489 29871 27523
rect 30021 27489 30055 27523
rect 30389 27489 30423 27523
rect 2421 27421 2455 27455
rect 2697 27421 2731 27455
rect 4445 27421 4479 27455
rect 5273 27421 5307 27455
rect 5914 27421 5948 27455
rect 6377 27421 6411 27455
rect 7665 27421 7699 27455
rect 8585 27421 8619 27455
rect 9137 27421 9171 27455
rect 9505 27421 9539 27455
rect 10241 27421 10275 27455
rect 10425 27421 10459 27455
rect 11102 27421 11136 27455
rect 11713 27421 11747 27455
rect 11806 27421 11840 27455
rect 12173 27421 12207 27455
rect 12449 27421 12483 27455
rect 12633 27421 12667 27455
rect 13001 27421 13035 27455
rect 13185 27421 13219 27455
rect 13461 27421 13495 27455
rect 13553 27421 13587 27455
rect 13737 27421 13771 27455
rect 14657 27421 14691 27455
rect 14749 27421 14783 27455
rect 18889 27421 18923 27455
rect 19257 27421 19291 27455
rect 20729 27421 20763 27455
rect 21281 27421 21315 27455
rect 23581 27421 23615 27455
rect 23765 27421 23799 27455
rect 23949 27421 23983 27455
rect 25973 27421 26007 27455
rect 26893 27421 26927 27455
rect 27169 27421 27203 27455
rect 29745 27421 29779 27455
rect 29929 27421 29963 27455
rect 31033 27421 31067 27455
rect 31217 27421 31251 27455
rect 31677 27421 31711 27455
rect 31861 27421 31895 27455
rect 2605 27353 2639 27387
rect 4813 27353 4847 27387
rect 7941 27353 7975 27387
rect 8033 27353 8067 27387
rect 9413 27353 9447 27387
rect 12081 27353 12115 27387
rect 14197 27353 14231 27387
rect 15577 27353 15611 27387
rect 18613 27353 18647 27387
rect 21557 27353 21591 27387
rect 23305 27353 23339 27387
rect 23673 27353 23707 27387
rect 26249 27353 26283 27387
rect 26801 27353 26835 27387
rect 5365 27285 5399 27319
rect 5733 27285 5767 27319
rect 5917 27285 5951 27319
rect 10977 27285 11011 27319
rect 11161 27285 11195 27319
rect 20177 27285 20211 27319
rect 24501 27285 24535 27319
rect 26433 27285 26467 27319
rect 26617 27285 26651 27319
rect 27077 27285 27111 27319
rect 29561 27285 29595 27319
rect 30757 27285 30791 27319
rect 30941 27285 30975 27319
rect 32045 27285 32079 27319
rect 9321 27081 9355 27115
rect 17785 27081 17819 27115
rect 21189 27081 21223 27115
rect 24485 27081 24519 27115
rect 5181 27013 5215 27047
rect 12265 27013 12299 27047
rect 22477 27013 22511 27047
rect 24685 27013 24719 27047
rect 26157 27013 26191 27047
rect 2237 26945 2271 26979
rect 4813 26945 4847 26979
rect 7113 26945 7147 26979
rect 7297 26945 7331 26979
rect 7757 26945 7791 26979
rect 8953 26945 8987 26979
rect 10977 26945 11011 26979
rect 11345 26945 11379 26979
rect 12173 26945 12207 26979
rect 12633 26945 12667 26979
rect 13001 26945 13035 26979
rect 13185 26945 13219 26979
rect 14657 26945 14691 26979
rect 14749 26945 14783 26979
rect 14933 26945 14967 26979
rect 16681 26945 16715 26979
rect 16957 26945 16991 26979
rect 17233 26945 17267 26979
rect 17417 26945 17451 26979
rect 17693 26945 17727 26979
rect 17877 26945 17911 26979
rect 18061 26945 18095 26979
rect 18245 26945 18279 26979
rect 18337 26945 18371 26979
rect 18429 26945 18463 26979
rect 18705 26945 18739 26979
rect 20637 26945 20671 26979
rect 20821 26945 20855 26979
rect 20913 26945 20947 26979
rect 21005 26945 21039 26979
rect 21281 26945 21315 26979
rect 26065 26945 26099 26979
rect 26249 26945 26283 26979
rect 26387 26945 26421 26979
rect 27445 26945 27479 26979
rect 27537 26945 27571 26979
rect 34529 26945 34563 26979
rect 34622 26945 34656 26979
rect 34805 26945 34839 26979
rect 34897 26945 34931 26979
rect 34994 26945 35028 26979
rect 2513 26877 2547 26911
rect 4997 26877 5031 26911
rect 9045 26877 9079 26911
rect 10793 26877 10827 26911
rect 12725 26877 12759 26911
rect 14381 26877 14415 26911
rect 14841 26877 14875 26911
rect 17049 26877 17083 26911
rect 18981 26877 19015 26911
rect 21557 26877 21591 26911
rect 22201 26877 22235 26911
rect 24225 26877 24259 26911
rect 26525 26877 26559 26911
rect 3985 26809 4019 26843
rect 7757 26809 7791 26843
rect 11161 26809 11195 26843
rect 18613 26809 18647 26843
rect 21281 26809 21315 26843
rect 21373 26809 21407 26843
rect 5089 26741 5123 26775
rect 8953 26741 8987 26775
rect 20453 26741 20487 26775
rect 24317 26741 24351 26775
rect 24501 26741 24535 26775
rect 25881 26741 25915 26775
rect 27445 26741 27479 26775
rect 27813 26741 27847 26775
rect 35173 26741 35207 26775
rect 1672 26537 1706 26571
rect 3801 26537 3835 26571
rect 5273 26537 5307 26571
rect 5733 26537 5767 26571
rect 6285 26537 6319 26571
rect 7389 26537 7423 26571
rect 7757 26537 7791 26571
rect 11161 26537 11195 26571
rect 11529 26537 11563 26571
rect 16129 26537 16163 26571
rect 17693 26537 17727 26571
rect 18153 26537 18187 26571
rect 22201 26537 22235 26571
rect 26525 26537 26559 26571
rect 31677 26537 31711 26571
rect 31953 26537 31987 26571
rect 32229 26537 32263 26571
rect 5917 26469 5951 26503
rect 13277 26469 13311 26503
rect 20269 26469 20303 26503
rect 23489 26469 23523 26503
rect 1409 26401 1443 26435
rect 3157 26401 3191 26435
rect 4261 26401 4295 26435
rect 4353 26401 4387 26435
rect 5549 26401 5583 26435
rect 7481 26401 7515 26435
rect 13369 26401 13403 26435
rect 16497 26401 16531 26435
rect 20821 26401 20855 26435
rect 25513 26401 25547 26435
rect 31677 26401 31711 26435
rect 4169 26333 4203 26367
rect 4721 26333 4755 26367
rect 5825 26333 5859 26367
rect 6193 26333 6227 26367
rect 6285 26333 6319 26367
rect 7389 26333 7423 26367
rect 11069 26333 11103 26367
rect 11253 26333 11287 26367
rect 11437 26333 11471 26367
rect 11621 26333 11655 26367
rect 12633 26333 12667 26367
rect 12726 26333 12760 26367
rect 13098 26333 13132 26367
rect 13553 26333 13587 26367
rect 13737 26333 13771 26367
rect 14289 26333 14323 26367
rect 14473 26333 14507 26367
rect 15025 26333 15059 26367
rect 15209 26333 15243 26367
rect 15853 26333 15887 26367
rect 16037 26333 16071 26367
rect 16405 26333 16439 26367
rect 16957 26333 16991 26367
rect 18061 26333 18095 26367
rect 18245 26333 18279 26367
rect 20361 26333 20395 26367
rect 20637 26333 20671 26367
rect 23305 26333 23339 26367
rect 25421 26333 25455 26367
rect 25605 26333 25639 26367
rect 25697 26333 25731 26367
rect 25881 26333 25915 26367
rect 25973 26333 26007 26367
rect 26249 26333 26283 26367
rect 26709 26333 26743 26367
rect 27077 26333 27111 26367
rect 27261 26333 27295 26367
rect 27353 26333 27387 26367
rect 27445 26333 27479 26367
rect 27537 26333 27571 26367
rect 27721 26333 27755 26367
rect 27869 26333 27903 26367
rect 27997 26333 28031 26367
rect 28089 26333 28123 26367
rect 28227 26333 28261 26367
rect 29561 26333 29595 26367
rect 29653 26333 29687 26367
rect 29837 26333 29871 26367
rect 29929 26333 29963 26367
rect 30113 26333 30147 26367
rect 31769 26333 31803 26367
rect 34069 26333 34103 26367
rect 34161 26333 34195 26367
rect 5089 26265 5123 26299
rect 12909 26265 12943 26299
rect 13001 26265 13035 26299
rect 14841 26265 14875 26299
rect 17325 26265 17359 26299
rect 17509 26265 17543 26299
rect 19993 26265 20027 26299
rect 21925 26265 21959 26299
rect 25789 26265 25823 26299
rect 27169 26265 27203 26299
rect 31493 26265 31527 26299
rect 32045 26265 32079 26299
rect 32245 26265 32279 26299
rect 14197 26197 14231 26231
rect 16037 26197 16071 26231
rect 26249 26197 26283 26231
rect 28365 26197 28399 26231
rect 32413 26197 32447 26231
rect 33885 26197 33919 26231
rect 2145 25993 2179 26027
rect 4445 25993 4479 26027
rect 4813 25993 4847 26027
rect 6101 25993 6135 26027
rect 14096 25993 14130 26027
rect 18889 25993 18923 26027
rect 19349 25993 19383 26027
rect 20085 25993 20119 26027
rect 23029 25993 23063 26027
rect 24225 25993 24259 26027
rect 29745 25993 29779 26027
rect 29913 25993 29947 26027
rect 32137 25993 32171 26027
rect 7297 25925 7331 25959
rect 7481 25925 7515 25959
rect 9137 25925 9171 25959
rect 9781 25925 9815 25959
rect 9873 25925 9907 25959
rect 10885 25925 10919 25959
rect 10977 25925 11011 25959
rect 12725 25925 12759 25959
rect 16313 25925 16347 25959
rect 17969 25925 18003 25959
rect 20269 25925 20303 25959
rect 21097 25925 21131 25959
rect 22753 25925 22787 25959
rect 23489 25925 23523 25959
rect 30113 25925 30147 25959
rect 32413 25925 32447 25959
rect 6009 25857 6043 25891
rect 6193 25857 6227 25891
rect 7573 25857 7607 25891
rect 7941 25857 7975 25891
rect 8769 25857 8803 25891
rect 8862 25857 8896 25891
rect 9045 25857 9079 25891
rect 9275 25857 9309 25891
rect 9505 25857 9539 25891
rect 9598 25857 9632 25891
rect 9970 25857 10004 25891
rect 10609 25857 10643 25891
rect 10701 25857 10735 25891
rect 11069 25857 11103 25891
rect 11897 25857 11931 25891
rect 12357 25857 12391 25891
rect 12450 25857 12484 25891
rect 12633 25857 12667 25891
rect 12822 25857 12856 25891
rect 13829 25857 13863 25891
rect 14473 25857 14507 25891
rect 14840 25857 14874 25891
rect 14933 25857 14967 25891
rect 15025 25857 15059 25891
rect 15209 25857 15243 25891
rect 15945 25857 15979 25891
rect 17601 25857 17635 25891
rect 18153 25857 18187 25891
rect 18429 25857 18463 25891
rect 18613 25857 18647 25891
rect 19073 25857 19107 25891
rect 20637 25857 20671 25891
rect 22017 25857 22051 25891
rect 22109 25857 22143 25891
rect 22293 25857 22327 25891
rect 22385 25857 22419 25891
rect 22569 25857 22603 25891
rect 23213 25857 23247 25891
rect 23581 25857 23615 25891
rect 23674 25857 23708 25891
rect 23857 25857 23891 25891
rect 23949 25857 23983 25891
rect 24087 25857 24121 25891
rect 24501 25857 24535 25891
rect 24593 25857 24627 25891
rect 24869 25857 24903 25891
rect 25329 25857 25363 25891
rect 26065 25857 26099 25891
rect 27537 25857 27571 25891
rect 27721 25857 27755 25891
rect 28917 25857 28951 25891
rect 29101 25857 29135 25891
rect 29469 25857 29503 25891
rect 29561 25857 29595 25891
rect 32289 25857 32323 25891
rect 32505 25857 32539 25891
rect 32689 25857 32723 25891
rect 32781 25857 32815 25891
rect 33517 25857 33551 25891
rect 33793 25857 33827 25891
rect 34069 25857 34103 25891
rect 2237 25789 2271 25823
rect 2421 25789 2455 25823
rect 2605 25789 2639 25823
rect 2881 25789 2915 25823
rect 4905 25789 4939 25823
rect 5089 25789 5123 25823
rect 5825 25789 5859 25823
rect 11161 25789 11195 25823
rect 11714 25789 11748 25823
rect 11805 25789 11839 25823
rect 11989 25789 12023 25823
rect 14565 25789 14599 25823
rect 15669 25789 15703 25823
rect 15853 25789 15887 25823
rect 17417 25789 17451 25823
rect 17877 25789 17911 25823
rect 18337 25789 18371 25823
rect 18521 25789 18555 25823
rect 19165 25789 19199 25823
rect 19441 25789 19475 25823
rect 19533 25789 19567 25823
rect 21189 25789 21223 25823
rect 21373 25789 21407 25823
rect 23397 25789 23431 25823
rect 24317 25789 24351 25823
rect 29009 25789 29043 25823
rect 33701 25789 33735 25823
rect 34345 25789 34379 25823
rect 36093 25789 36127 25823
rect 22937 25721 22971 25755
rect 25973 25721 26007 25755
rect 27721 25721 27755 25755
rect 33977 25721 34011 25755
rect 1777 25653 1811 25687
rect 4353 25653 4387 25687
rect 5273 25653 5307 25687
rect 7021 25653 7055 25687
rect 7849 25653 7883 25687
rect 9413 25653 9447 25687
rect 10149 25653 10183 25687
rect 11529 25653 11563 25687
rect 13001 25653 13035 25687
rect 14105 25653 14139 25687
rect 17785 25653 17819 25687
rect 20269 25653 20303 25687
rect 20729 25653 20763 25687
rect 21833 25653 21867 25687
rect 23397 25653 23431 25687
rect 24777 25653 24811 25687
rect 29285 25653 29319 25687
rect 29929 25653 29963 25687
rect 33517 25653 33551 25687
rect 3157 25449 3191 25483
rect 4813 25449 4847 25483
rect 6653 25449 6687 25483
rect 9781 25449 9815 25483
rect 18153 25449 18187 25483
rect 19625 25449 19659 25483
rect 23305 25449 23339 25483
rect 24869 25449 24903 25483
rect 33333 25449 33367 25483
rect 33793 25449 33827 25483
rect 35909 25449 35943 25483
rect 8493 25381 8527 25415
rect 16589 25381 16623 25415
rect 20361 25381 20395 25415
rect 23489 25381 23523 25415
rect 25053 25381 25087 25415
rect 32781 25381 32815 25415
rect 33701 25381 33735 25415
rect 1409 25313 1443 25347
rect 4537 25313 4571 25347
rect 5273 25313 5307 25347
rect 5457 25313 5491 25347
rect 7297 25313 7331 25347
rect 8125 25313 8159 25347
rect 8309 25313 8343 25347
rect 9965 25313 9999 25347
rect 14933 25313 14967 25347
rect 16405 25313 16439 25347
rect 23213 25313 23247 25347
rect 5917 25245 5951 25279
rect 6561 25245 6595 25279
rect 7205 25245 7239 25279
rect 7389 25245 7423 25279
rect 8033 25245 8067 25279
rect 8217 25245 8251 25279
rect 9229 25245 9263 25279
rect 9413 25245 9447 25279
rect 9597 25245 9631 25279
rect 9873 25245 9907 25279
rect 10057 25245 10091 25279
rect 11529 25245 11563 25279
rect 11621 25245 11655 25279
rect 11713 25245 11747 25279
rect 14473 25245 14507 25279
rect 14565 25245 14599 25279
rect 14657 25245 14691 25279
rect 15117 25245 15151 25279
rect 15393 25245 15427 25279
rect 16221 25245 16255 25279
rect 16773 25245 16807 25279
rect 17601 25245 17635 25279
rect 17877 25245 17911 25279
rect 17969 25245 18003 25279
rect 18981 25245 19015 25279
rect 20729 25245 20763 25279
rect 20913 25245 20947 25279
rect 21465 25245 21499 25279
rect 21557 25245 21591 25279
rect 21741 25245 21775 25279
rect 21833 25245 21867 25279
rect 23121 25245 23155 25279
rect 32137 25255 32171 25289
rect 32275 25245 32309 25279
rect 32629 25245 32663 25279
rect 33609 25245 33643 25279
rect 34069 25245 34103 25279
rect 35725 25245 35759 25279
rect 32505 25211 32539 25245
rect 1685 25177 1719 25211
rect 3801 25177 3835 25211
rect 6469 25177 6503 25211
rect 6837 25177 6871 25211
rect 6929 25177 6963 25211
rect 9505 25177 9539 25211
rect 11437 25177 11471 25211
rect 11897 25177 11931 25211
rect 14749 25177 14783 25211
rect 16037 25177 16071 25211
rect 17785 25177 17819 25211
rect 18613 25177 18647 25211
rect 19809 25177 19843 25211
rect 20361 25177 20395 25211
rect 21925 25177 21959 25211
rect 22109 25177 22143 25211
rect 22293 25177 22327 25211
rect 25329 25177 25363 25211
rect 32413 25177 32447 25211
rect 5181 25109 5215 25143
rect 5733 25109 5767 25143
rect 15117 25109 15151 25143
rect 15853 25109 15887 25143
rect 16129 25109 16163 25143
rect 19901 25109 19935 25143
rect 20545 25109 20579 25143
rect 21281 25109 21315 25143
rect 33977 25109 34011 25143
rect 12173 24905 12207 24939
rect 16313 24905 16347 24939
rect 22753 24905 22787 24939
rect 28733 24905 28767 24939
rect 35909 24905 35943 24939
rect 2605 24837 2639 24871
rect 2697 24837 2731 24871
rect 6377 24837 6411 24871
rect 8401 24837 8435 24871
rect 3709 24769 3743 24803
rect 6561 24769 6595 24803
rect 6929 24769 6963 24803
rect 7021 24769 7055 24803
rect 7113 24769 7147 24803
rect 8585 24769 8619 24803
rect 8677 24769 8711 24803
rect 9137 24769 9171 24803
rect 9230 24769 9264 24803
rect 9413 24769 9447 24803
rect 9505 24769 9539 24803
rect 9602 24769 9636 24803
rect 11161 24769 11195 24803
rect 11345 24769 11379 24803
rect 11529 24769 11563 24803
rect 11622 24769 11656 24803
rect 11805 24769 11839 24803
rect 11897 24769 11931 24803
rect 12035 24769 12069 24803
rect 12265 24769 12299 24803
rect 12449 24769 12483 24803
rect 12541 24769 12575 24803
rect 12653 24769 12687 24803
rect 12817 24769 12851 24803
rect 13001 24769 13035 24803
rect 13093 24769 13127 24803
rect 16313 24769 16347 24803
rect 16497 24769 16531 24803
rect 17141 24769 17175 24803
rect 17233 24769 17267 24803
rect 17417 24769 17451 24803
rect 17969 24769 18003 24803
rect 18797 24769 18831 24803
rect 18981 24769 19015 24803
rect 19257 24769 19291 24803
rect 19625 24769 19659 24803
rect 22937 24769 22971 24803
rect 23397 24769 23431 24803
rect 23673 24769 23707 24803
rect 25697 24769 25731 24803
rect 25790 24769 25824 24803
rect 25973 24769 26007 24803
rect 26065 24769 26099 24803
rect 26162 24769 26196 24803
rect 27261 24769 27295 24803
rect 27445 24769 27479 24803
rect 27537 24769 27571 24803
rect 28273 24769 28307 24803
rect 29009 24769 29043 24803
rect 29147 24769 29181 24803
rect 33885 24769 33919 24803
rect 34069 24769 34103 24803
rect 35173 24769 35207 24803
rect 35357 24769 35391 24803
rect 36001 24769 36035 24803
rect 28181 24735 28215 24769
rect 2789 24701 2823 24735
rect 3985 24701 4019 24735
rect 6193 24701 6227 24735
rect 18889 24701 18923 24735
rect 23121 24701 23155 24735
rect 23489 24701 23523 24735
rect 23949 24701 23983 24735
rect 28365 24701 28399 24735
rect 28457 24701 28491 24735
rect 28917 24701 28951 24735
rect 29285 24701 29319 24735
rect 29377 24701 29411 24735
rect 5457 24633 5491 24667
rect 8401 24633 8435 24667
rect 12265 24633 12299 24667
rect 16681 24633 16715 24667
rect 26341 24633 26375 24667
rect 27721 24633 27755 24667
rect 28641 24633 28675 24667
rect 2237 24565 2271 24599
rect 5549 24565 5583 24599
rect 6653 24565 6687 24599
rect 9781 24565 9815 24599
rect 11345 24565 11379 24599
rect 12817 24565 12851 24599
rect 16957 24565 16991 24599
rect 17049 24565 17083 24599
rect 17877 24565 17911 24599
rect 23305 24565 23339 24599
rect 23857 24565 23891 24599
rect 27537 24565 27571 24599
rect 33885 24565 33919 24599
rect 34253 24565 34287 24599
rect 35541 24565 35575 24599
rect 3157 24361 3191 24395
rect 4813 24361 4847 24395
rect 5733 24361 5767 24395
rect 11621 24361 11655 24395
rect 14289 24361 14323 24395
rect 14933 24361 14967 24395
rect 17141 24361 17175 24395
rect 18981 24361 19015 24395
rect 20085 24361 20119 24395
rect 20637 24361 20671 24395
rect 21097 24361 21131 24395
rect 21373 24361 21407 24395
rect 25329 24361 25363 24395
rect 26617 24361 26651 24395
rect 27905 24361 27939 24395
rect 31585 24361 31619 24395
rect 31769 24361 31803 24395
rect 35909 24361 35943 24395
rect 6653 24293 6687 24327
rect 7297 24293 7331 24327
rect 9321 24293 9355 24327
rect 12173 24293 12207 24327
rect 12357 24293 12391 24327
rect 17601 24293 17635 24327
rect 21189 24293 21223 24327
rect 27261 24293 27295 24327
rect 1685 24225 1719 24259
rect 5273 24225 5307 24259
rect 5457 24225 5491 24259
rect 8217 24225 8251 24259
rect 15025 24225 15059 24259
rect 15117 24225 15151 24259
rect 17233 24225 17267 24259
rect 17325 24225 17359 24259
rect 19809 24225 19843 24259
rect 19901 24225 19935 24259
rect 24593 24225 24627 24259
rect 31493 24225 31527 24259
rect 1409 24157 1443 24191
rect 6837 24157 6871 24191
rect 6929 24157 6963 24191
rect 7021 24157 7055 24191
rect 7297 24157 7331 24191
rect 7389 24157 7423 24191
rect 9500 24157 9534 24191
rect 9817 24157 9851 24191
rect 9965 24157 9999 24191
rect 10236 24157 10270 24191
rect 10333 24157 10367 24191
rect 10553 24157 10587 24191
rect 10701 24157 10735 24191
rect 11069 24157 11103 24191
rect 11253 24157 11287 24191
rect 11437 24157 11471 24191
rect 13001 24157 13035 24191
rect 13094 24157 13128 24191
rect 13277 24157 13311 24191
rect 13466 24157 13500 24191
rect 14473 24157 14507 24191
rect 14565 24157 14599 24191
rect 14841 24157 14875 24191
rect 16865 24157 16899 24191
rect 18797 24157 18831 24191
rect 18981 24157 19015 24191
rect 19441 24157 19475 24191
rect 19533 24157 19567 24191
rect 20269 24157 20303 24191
rect 20361 24157 20395 24191
rect 20821 24157 20855 24191
rect 20913 24157 20947 24191
rect 24465 24157 24499 24191
rect 25053 24157 25087 24191
rect 25145 24157 25179 24191
rect 26065 24157 26099 24191
rect 26341 24157 26375 24191
rect 26433 24157 26467 24191
rect 26709 24157 26743 24191
rect 26985 24157 27019 24191
rect 27077 24157 27111 24191
rect 27353 24157 27387 24191
rect 27537 24157 27571 24191
rect 27721 24157 27755 24191
rect 30665 24157 30699 24191
rect 30849 24157 30883 24191
rect 31033 24157 31067 24191
rect 31585 24157 31619 24191
rect 36093 24157 36127 24191
rect 5181 24089 5215 24123
rect 5825 24089 5859 24123
rect 6009 24089 6043 24123
rect 6653 24089 6687 24123
rect 9597 24089 9631 24123
rect 9689 24089 9723 24123
rect 10425 24089 10459 24123
rect 11345 24089 11379 24123
rect 12633 24089 12667 24123
rect 13389 24089 13423 24123
rect 14657 24089 14691 24123
rect 15393 24089 15427 24123
rect 20085 24089 20119 24123
rect 20637 24089 20671 24123
rect 21557 24089 21591 24123
rect 24593 24089 24627 24123
rect 24685 24089 24719 24123
rect 24869 24089 24903 24123
rect 26249 24089 26283 24123
rect 26893 24089 26927 24123
rect 27629 24089 27663 24123
rect 30941 24089 30975 24123
rect 31309 24089 31343 24123
rect 7113 24021 7147 24055
rect 10057 24021 10091 24055
rect 13645 24021 13679 24055
rect 15301 24021 15335 24055
rect 16957 24021 16991 24055
rect 19257 24021 19291 24055
rect 20545 24021 20579 24055
rect 21357 24021 21391 24055
rect 31217 24021 31251 24055
rect 7021 23817 7055 23851
rect 8861 23817 8895 23851
rect 13001 23817 13035 23851
rect 15669 23817 15703 23851
rect 20177 23817 20211 23851
rect 20821 23817 20855 23851
rect 26249 23817 26283 23851
rect 29101 23817 29135 23851
rect 4353 23749 4387 23783
rect 5365 23749 5399 23783
rect 6745 23749 6779 23783
rect 9045 23749 9079 23783
rect 11697 23749 11731 23783
rect 11897 23749 11931 23783
rect 17877 23749 17911 23783
rect 18061 23749 18095 23783
rect 19809 23749 19843 23783
rect 20009 23749 20043 23783
rect 20269 23749 20303 23783
rect 22293 23749 22327 23783
rect 25973 23749 26007 23783
rect 28733 23749 28767 23783
rect 30849 23749 30883 23783
rect 5181 23681 5215 23715
rect 5457 23681 5491 23715
rect 5549 23681 5583 23715
rect 6009 23681 6043 23715
rect 6193 23681 6227 23715
rect 6377 23681 6411 23715
rect 6470 23681 6504 23715
rect 6653 23681 6687 23715
rect 6883 23681 6917 23715
rect 7941 23681 7975 23715
rect 8309 23681 8343 23715
rect 8769 23681 8803 23715
rect 13180 23681 13214 23715
rect 13277 23681 13311 23715
rect 13369 23681 13403 23715
rect 13552 23681 13586 23715
rect 13645 23681 13679 23715
rect 15485 23681 15519 23715
rect 15761 23681 15795 23715
rect 18613 23681 18647 23715
rect 18889 23681 18923 23715
rect 19165 23681 19199 23715
rect 20453 23681 20487 23715
rect 20545 23681 20579 23715
rect 22477 23681 22511 23715
rect 25329 23681 25363 23715
rect 25697 23681 25731 23715
rect 25881 23681 25915 23715
rect 26065 23681 26099 23715
rect 28549 23681 28583 23715
rect 28825 23681 28859 23715
rect 28917 23681 28951 23715
rect 29193 23681 29227 23715
rect 29285 23681 29319 23715
rect 30711 23681 30745 23715
rect 30941 23681 30975 23715
rect 31033 23681 31067 23715
rect 33333 23681 33367 23715
rect 34437 23681 34471 23715
rect 34621 23681 34655 23715
rect 34713 23681 34747 23715
rect 1593 23613 1627 23647
rect 1869 23613 1903 23647
rect 3525 23613 3559 23647
rect 5089 23613 5123 23647
rect 18521 23613 18555 23647
rect 18981 23613 19015 23647
rect 21005 23613 21039 23647
rect 21097 23613 21131 23647
rect 21465 23613 21499 23647
rect 25145 23613 25179 23647
rect 30573 23613 30607 23647
rect 33057 23613 33091 23647
rect 3341 23545 3375 23579
rect 20269 23545 20303 23579
rect 25513 23545 25547 23579
rect 29561 23545 29595 23579
rect 33517 23545 33551 23579
rect 4445 23477 4479 23511
rect 5733 23477 5767 23511
rect 5917 23477 5951 23511
rect 9045 23477 9079 23511
rect 11529 23477 11563 23511
rect 11713 23477 11747 23511
rect 17693 23477 17727 23511
rect 17877 23477 17911 23511
rect 18245 23477 18279 23511
rect 18429 23477 18463 23511
rect 18705 23477 18739 23511
rect 18981 23477 19015 23511
rect 19993 23477 20027 23511
rect 22661 23477 22695 23511
rect 29377 23477 29411 23511
rect 31217 23477 31251 23511
rect 33149 23477 33183 23511
rect 34529 23477 34563 23511
rect 34897 23477 34931 23511
rect 6285 23273 6319 23307
rect 6745 23273 6779 23307
rect 13093 23273 13127 23307
rect 17049 23273 17083 23307
rect 17233 23273 17267 23307
rect 17601 23273 17635 23307
rect 21649 23273 21683 23307
rect 22293 23273 22327 23307
rect 25605 23273 25639 23307
rect 28457 23273 28491 23307
rect 13369 23205 13403 23239
rect 14381 23205 14415 23239
rect 17417 23205 17451 23239
rect 4353 23137 4387 23171
rect 11161 23137 11195 23171
rect 13737 23137 13771 23171
rect 18337 23137 18371 23171
rect 18521 23137 18555 23171
rect 18613 23137 18647 23171
rect 21557 23137 21591 23171
rect 1409 23069 1443 23103
rect 3249 23069 3283 23103
rect 4905 23069 4939 23103
rect 4998 23069 5032 23103
rect 5181 23069 5215 23103
rect 5411 23069 5445 23103
rect 5641 23069 5675 23103
rect 5779 23069 5813 23103
rect 5917 23069 5951 23103
rect 6106 23069 6140 23103
rect 7113 23069 7147 23103
rect 7206 23069 7240 23103
rect 7578 23069 7612 23103
rect 8401 23069 8435 23103
rect 8585 23069 8619 23103
rect 8769 23069 8803 23103
rect 11352 23069 11386 23103
rect 11493 23069 11527 23103
rect 11810 23069 11844 23103
rect 12081 23069 12115 23103
rect 12265 23069 12299 23103
rect 12633 23069 12667 23103
rect 12725 23069 12759 23103
rect 13093 23069 13127 23103
rect 13277 23069 13311 23103
rect 13553 23069 13587 23103
rect 14657 23069 14691 23103
rect 15025 23069 15059 23103
rect 15485 23069 15519 23103
rect 15761 23069 15795 23103
rect 15945 23069 15979 23103
rect 16129 23069 16163 23103
rect 16865 23069 16899 23103
rect 16957 23069 16991 23103
rect 18429 23069 18463 23103
rect 21833 23069 21867 23103
rect 22845 23069 22879 23103
rect 23029 23069 23063 23103
rect 23121 23069 23155 23103
rect 25789 23069 25823 23103
rect 25881 23069 25915 23103
rect 27905 23069 27939 23103
rect 28273 23069 28307 23103
rect 1685 23001 1719 23035
rect 4169 23001 4203 23035
rect 5273 23001 5307 23035
rect 6009 23001 6043 23035
rect 6837 23001 6871 23035
rect 7021 23001 7055 23035
rect 7389 23001 7423 23035
rect 7481 23001 7515 23035
rect 8493 23001 8527 23035
rect 11621 23001 11655 23035
rect 11713 23001 11747 23035
rect 12449 23001 12483 23035
rect 17785 23001 17819 23035
rect 22017 23001 22051 23035
rect 22109 23001 22143 23035
rect 22309 23001 22343 23035
rect 28089 23001 28123 23035
rect 28181 23001 28215 23035
rect 3157 22933 3191 22967
rect 3801 22933 3835 22967
rect 4261 22933 4295 22967
rect 5549 22933 5583 22967
rect 7757 22933 7791 22967
rect 8217 22933 8251 22967
rect 10609 22933 10643 22967
rect 11989 22933 12023 22967
rect 12173 22933 12207 22967
rect 12909 22933 12943 22967
rect 16037 22933 16071 22967
rect 17585 22933 17619 22967
rect 18153 22933 18187 22967
rect 22477 22933 22511 22967
rect 22661 22933 22695 22967
rect 1777 22729 1811 22763
rect 2145 22729 2179 22763
rect 5181 22729 5215 22763
rect 6929 22729 6963 22763
rect 8493 22729 8527 22763
rect 9873 22729 9907 22763
rect 10241 22729 10275 22763
rect 10333 22729 10367 22763
rect 14013 22729 14047 22763
rect 14933 22729 14967 22763
rect 15301 22729 15335 22763
rect 19901 22729 19935 22763
rect 20637 22729 20671 22763
rect 23397 22729 23431 22763
rect 25421 22729 25455 22763
rect 32781 22729 32815 22763
rect 35909 22729 35943 22763
rect 4077 22661 4111 22695
rect 5457 22661 5491 22695
rect 6561 22661 6595 22695
rect 6653 22661 6687 22695
rect 8125 22661 8159 22695
rect 8953 22661 8987 22695
rect 9413 22661 9447 22695
rect 9781 22661 9815 22695
rect 10977 22661 11011 22695
rect 11069 22661 11103 22695
rect 11897 22661 11931 22695
rect 11989 22661 12023 22695
rect 12909 22661 12943 22695
rect 13185 22661 13219 22695
rect 14381 22661 14415 22695
rect 14565 22661 14599 22695
rect 22569 22661 22603 22695
rect 32413 22661 32447 22695
rect 32505 22661 32539 22695
rect 2237 22593 2271 22627
rect 4353 22593 4387 22627
rect 5365 22593 5399 22627
rect 5549 22593 5583 22627
rect 5733 22593 5767 22627
rect 5825 22593 5859 22627
rect 6009 22593 6043 22627
rect 6377 22593 6411 22627
rect 6745 22593 6779 22627
rect 7849 22593 7883 22627
rect 7997 22593 8031 22627
rect 8217 22593 8251 22627
rect 8314 22593 8348 22627
rect 8585 22593 8619 22627
rect 8678 22593 8712 22627
rect 8861 22593 8895 22627
rect 9050 22593 9084 22627
rect 9597 22593 9631 22627
rect 10839 22593 10873 22627
rect 11161 22593 11195 22627
rect 11759 22593 11793 22627
rect 12172 22593 12206 22627
rect 12265 22593 12299 22627
rect 13460 22593 13494 22627
rect 13553 22593 13587 22627
rect 13645 22593 13679 22627
rect 13829 22593 13863 22627
rect 14013 22593 14047 22627
rect 14289 22593 14323 22627
rect 14657 22593 14691 22627
rect 15117 22593 15151 22627
rect 15577 22593 15611 22627
rect 15945 22593 15979 22627
rect 16129 22593 16163 22627
rect 18245 22593 18279 22627
rect 18429 22593 18463 22627
rect 18521 22593 18555 22627
rect 20085 22593 20119 22627
rect 20545 22593 20579 22627
rect 22109 22593 22143 22627
rect 22293 22593 22327 22627
rect 23581 22593 23615 22627
rect 23765 22593 23799 22627
rect 23995 22593 24029 22627
rect 24133 22593 24167 22627
rect 24225 22593 24259 22627
rect 24408 22593 24442 22627
rect 24501 22593 24535 22627
rect 25605 22593 25639 22627
rect 27537 22593 27571 22627
rect 28457 22593 28491 22627
rect 28641 22593 28675 22627
rect 32137 22593 32171 22627
rect 32230 22593 32264 22627
rect 32641 22593 32675 22627
rect 33333 22593 33367 22627
rect 33425 22593 33459 22627
rect 34529 22593 34563 22627
rect 34805 22593 34839 22627
rect 36093 22593 36127 22627
rect 2421 22525 2455 22559
rect 5089 22525 5123 22559
rect 7113 22525 7147 22559
rect 7665 22525 7699 22559
rect 10425 22525 10459 22559
rect 10701 22525 10735 22559
rect 15209 22525 15243 22559
rect 15485 22525 15519 22559
rect 18061 22525 18095 22559
rect 20361 22525 20395 22559
rect 25789 22525 25823 22559
rect 27813 22525 27847 22559
rect 34621 22525 34655 22559
rect 9229 22457 9263 22491
rect 12449 22457 12483 22491
rect 12541 22457 12575 22491
rect 14381 22457 14415 22491
rect 21925 22457 21959 22491
rect 2605 22389 2639 22423
rect 4445 22389 4479 22423
rect 6101 22389 6135 22423
rect 11345 22389 11379 22423
rect 11621 22389 11655 22423
rect 15761 22389 15795 22423
rect 20269 22389 20303 22423
rect 22477 22389 22511 22423
rect 23765 22389 23799 22423
rect 23857 22389 23891 22423
rect 28457 22389 28491 22423
rect 33517 22389 33551 22423
rect 33701 22389 33735 22423
rect 34529 22389 34563 22423
rect 34989 22389 35023 22423
rect 2329 22185 2363 22219
rect 4445 22185 4479 22219
rect 5457 22185 5491 22219
rect 9308 22185 9342 22219
rect 13369 22185 13403 22219
rect 13829 22185 13863 22219
rect 17233 22185 17267 22219
rect 23121 22185 23155 22219
rect 35265 22185 35299 22219
rect 11069 22117 11103 22151
rect 13001 22117 13035 22151
rect 14841 22117 14875 22151
rect 17417 22117 17451 22151
rect 23029 22117 23063 22151
rect 2789 22049 2823 22083
rect 2973 22049 3007 22083
rect 3893 22049 3927 22083
rect 6929 22049 6963 22083
rect 8217 22049 8251 22083
rect 12081 22049 12115 22083
rect 15209 22049 15243 22083
rect 15393 22049 15427 22083
rect 15761 22049 15795 22083
rect 16865 22049 16899 22083
rect 19349 22049 19383 22083
rect 19533 22049 19567 22083
rect 21465 22049 21499 22083
rect 23213 22049 23247 22083
rect 26065 22049 26099 22083
rect 27261 22049 27295 22083
rect 27905 22049 27939 22083
rect 35817 22049 35851 22083
rect 4905 21981 4939 22015
rect 5273 21981 5307 22015
rect 6653 21981 6687 22015
rect 7481 21981 7515 22015
rect 9045 21981 9079 22015
rect 11253 21981 11287 22015
rect 11345 21981 11379 22015
rect 11529 21981 11563 22015
rect 11621 21981 11655 22015
rect 11805 21981 11839 22015
rect 11989 21981 12023 22015
rect 12449 21981 12483 22015
rect 12633 21981 12667 22015
rect 12725 21981 12759 22015
rect 13185 21981 13219 22015
rect 13461 21981 13495 22015
rect 13553 21981 13587 22015
rect 13737 21981 13771 22015
rect 13829 21981 13863 22015
rect 15025 21981 15059 22015
rect 15301 21981 15335 22015
rect 15577 21981 15611 22015
rect 15853 21981 15887 22015
rect 16129 21981 16163 22015
rect 19625 21981 19659 22015
rect 19717 21981 19751 22015
rect 19901 21981 19935 22015
rect 20085 21981 20119 22015
rect 21741 21981 21775 22015
rect 23305 21981 23339 22015
rect 23489 21981 23523 22015
rect 26249 21981 26283 22015
rect 27537 21981 27571 22015
rect 27721 21981 27755 22015
rect 28273 21981 28307 22015
rect 30205 21981 30239 22015
rect 30573 21981 30607 22015
rect 35173 21981 35207 22015
rect 35357 21981 35391 22015
rect 36093 21981 36127 22015
rect 2697 21913 2731 21947
rect 5089 21913 5123 21947
rect 5181 21913 5215 21947
rect 6745 21913 6779 21947
rect 11897 21913 11931 21947
rect 12265 21913 12299 21947
rect 21256 21913 21290 21947
rect 22845 21913 22879 21947
rect 27399 21913 27433 21947
rect 27629 21913 27663 21947
rect 30297 21913 30331 21947
rect 30389 21913 30423 21947
rect 6285 21845 6319 21879
rect 10793 21845 10827 21879
rect 16037 21845 16071 21879
rect 17233 21845 17267 21879
rect 19993 21845 20027 21879
rect 21097 21845 21131 21879
rect 21373 21845 21407 21879
rect 26433 21845 26467 21879
rect 28089 21845 28123 21879
rect 30021 21845 30055 21879
rect 35541 21845 35575 21879
rect 12449 21641 12483 21675
rect 12617 21641 12651 21675
rect 13645 21641 13679 21675
rect 17509 21641 17543 21675
rect 18889 21641 18923 21675
rect 20177 21641 20211 21675
rect 20361 21641 20395 21675
rect 35909 21641 35943 21675
rect 4261 21573 4295 21607
rect 6653 21573 6687 21607
rect 10977 21573 11011 21607
rect 11069 21573 11103 21607
rect 11897 21573 11931 21607
rect 12817 21573 12851 21607
rect 18613 21573 18647 21607
rect 23841 21573 23875 21607
rect 24041 21573 24075 21607
rect 29101 21573 29135 21607
rect 4077 21505 4111 21539
rect 4353 21505 4387 21539
rect 4445 21505 4479 21539
rect 6377 21505 6411 21539
rect 8396 21505 8430 21539
rect 8493 21505 8527 21539
rect 8585 21505 8619 21539
rect 8768 21505 8802 21539
rect 8861 21505 8895 21539
rect 8953 21505 8987 21539
rect 10793 21505 10827 21539
rect 11161 21505 11195 21539
rect 11713 21505 11747 21539
rect 11805 21505 11839 21539
rect 12081 21505 12115 21539
rect 14197 21505 14231 21539
rect 17233 21505 17267 21539
rect 18245 21505 18279 21539
rect 18393 21505 18427 21539
rect 18521 21505 18555 21539
rect 18710 21505 18744 21539
rect 19441 21505 19475 21539
rect 19717 21505 19751 21539
rect 19809 21505 19843 21539
rect 20269 21505 20303 21539
rect 20453 21505 20487 21539
rect 28825 21505 28859 21539
rect 28918 21505 28952 21539
rect 29193 21505 29227 21539
rect 29290 21505 29324 21539
rect 29561 21505 29595 21539
rect 36093 21505 36127 21539
rect 1409 21437 1443 21471
rect 1685 21437 1719 21471
rect 3157 21437 3191 21471
rect 3893 21437 3927 21471
rect 9229 21437 9263 21471
rect 10701 21437 10735 21471
rect 13921 21437 13955 21471
rect 17509 21437 17543 21471
rect 19901 21437 19935 21471
rect 8217 21369 8251 21403
rect 19257 21369 19291 21403
rect 29469 21369 29503 21403
rect 3249 21301 3283 21335
rect 4629 21301 4663 21335
rect 8125 21301 8159 21335
rect 11345 21301 11379 21335
rect 11529 21301 11563 21335
rect 12633 21301 12667 21335
rect 13829 21301 13863 21335
rect 17325 21301 17359 21335
rect 19625 21301 19659 21335
rect 19809 21301 19843 21335
rect 23673 21301 23707 21335
rect 23857 21301 23891 21335
rect 29745 21301 29779 21335
rect 2145 21097 2179 21131
rect 9781 21097 9815 21131
rect 11897 21097 11931 21131
rect 12173 21097 12207 21131
rect 14105 21097 14139 21131
rect 17233 21097 17267 21131
rect 21649 21097 21683 21131
rect 22937 21097 22971 21131
rect 23581 21097 23615 21131
rect 23949 21097 23983 21131
rect 25053 21097 25087 21131
rect 26893 21097 26927 21131
rect 32781 21097 32815 21131
rect 7481 21029 7515 21063
rect 11529 21029 11563 21063
rect 11621 21029 11655 21063
rect 12449 21029 12483 21063
rect 22661 21029 22695 21063
rect 23765 21029 23799 21063
rect 2605 20961 2639 20995
rect 2697 20961 2731 20995
rect 7389 20961 7423 20995
rect 8769 20961 8803 20995
rect 9413 20961 9447 20995
rect 9505 20961 9539 20995
rect 10425 20961 10459 20995
rect 11161 20961 11195 20995
rect 15117 20961 15151 20995
rect 15393 20961 15427 20995
rect 23029 20961 23063 20995
rect 32873 20961 32907 20995
rect 2513 20893 2547 20927
rect 2973 20893 3007 20927
rect 3249 20893 3283 20927
rect 3341 20893 3375 20927
rect 4629 20893 4663 20927
rect 4905 20893 4939 20927
rect 4997 20893 5031 20927
rect 6745 20893 6779 20927
rect 7021 20893 7055 20927
rect 7113 20893 7147 20927
rect 7665 20893 7699 20927
rect 7756 20893 7790 20927
rect 10241 20893 10275 20927
rect 11437 20893 11471 20927
rect 11713 20893 11747 20927
rect 12633 20893 12667 20927
rect 12725 20893 12759 20927
rect 13185 20893 13219 20927
rect 13461 20893 13495 20927
rect 13553 20893 13587 20927
rect 14105 20893 14139 20927
rect 14289 20893 14323 20927
rect 15209 20893 15243 20927
rect 15301 20893 15335 20927
rect 16313 20893 16347 20927
rect 16957 20893 16991 20927
rect 17049 20893 17083 20927
rect 21373 20893 21407 20927
rect 21465 20893 21499 20927
rect 21557 20893 21591 20927
rect 22845 20893 22879 20927
rect 23397 20893 23431 20927
rect 23489 20893 23523 20927
rect 23673 20893 23707 20927
rect 23949 20893 23983 20927
rect 24041 20893 24075 20927
rect 24409 20893 24443 20927
rect 24501 20893 24535 20927
rect 24685 20893 24719 20927
rect 24777 20893 24811 20927
rect 25237 20893 25271 20927
rect 25513 20893 25547 20927
rect 26249 20893 26283 20927
rect 27997 20893 28031 20927
rect 28365 20893 28399 20927
rect 28457 20893 28491 20927
rect 31493 20893 31527 20927
rect 31677 20893 31711 20927
rect 31769 20893 31803 20927
rect 33057 20893 33091 20927
rect 3157 20825 3191 20859
rect 4813 20825 4847 20859
rect 6929 20825 6963 20859
rect 9321 20825 9355 20859
rect 10149 20825 10183 20859
rect 10609 20825 10643 20859
rect 11989 20825 12023 20859
rect 13001 20825 13035 20859
rect 13093 20825 13127 20859
rect 13369 20825 13403 20859
rect 19349 20825 19383 20859
rect 21189 20825 21223 20859
rect 22201 20825 22235 20859
rect 22385 20825 22419 20859
rect 23121 20825 23155 20859
rect 24225 20825 24259 20859
rect 24961 20825 24995 20859
rect 25421 20825 25455 20859
rect 26709 20825 26743 20859
rect 26925 20825 26959 20859
rect 28155 20825 28189 20859
rect 28273 20825 28307 20859
rect 32781 20825 32815 20859
rect 3525 20757 3559 20791
rect 5181 20757 5215 20791
rect 7297 20757 7331 20791
rect 7941 20757 7975 20791
rect 8125 20757 8159 20791
rect 8953 20757 8987 20791
rect 12189 20757 12223 20791
rect 12357 20757 12391 20791
rect 13737 20757 13771 20791
rect 15577 20757 15611 20791
rect 15761 20757 15795 20791
rect 19441 20757 19475 20791
rect 22569 20757 22603 20791
rect 23213 20757 23247 20791
rect 26341 20757 26375 20791
rect 27077 20757 27111 20791
rect 28641 20757 28675 20791
rect 31309 20757 31343 20791
rect 33241 20757 33275 20791
rect 7757 20553 7791 20587
rect 10241 20553 10275 20587
rect 11713 20553 11747 20587
rect 13093 20553 13127 20587
rect 22293 20553 22327 20587
rect 24225 20553 24259 20587
rect 24961 20553 24995 20587
rect 34989 20553 35023 20587
rect 7849 20485 7883 20519
rect 8677 20485 8711 20519
rect 11897 20485 11931 20519
rect 15485 20485 15519 20519
rect 15945 20485 15979 20519
rect 16145 20485 16179 20519
rect 17509 20485 17543 20519
rect 17693 20485 17727 20519
rect 19993 20485 20027 20519
rect 20361 20485 20395 20519
rect 20913 20485 20947 20519
rect 21129 20485 21163 20519
rect 21833 20485 21867 20519
rect 23857 20485 23891 20519
rect 27169 20485 27203 20519
rect 27813 20485 27847 20519
rect 28273 20485 28307 20519
rect 4445 20417 4479 20451
rect 4537 20417 4571 20451
rect 4905 20417 4939 20451
rect 5549 20417 5583 20451
rect 6929 20417 6963 20451
rect 7021 20417 7055 20451
rect 8401 20417 8435 20451
rect 10793 20417 10827 20451
rect 15577 20417 15611 20451
rect 16681 20417 16715 20451
rect 19917 20407 19951 20441
rect 20177 20417 20211 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 22845 20417 22879 20451
rect 23029 20417 23063 20451
rect 24041 20417 24075 20451
rect 25145 20417 25179 20451
rect 25513 20417 25547 20451
rect 25697 20417 25731 20451
rect 25789 20417 25823 20451
rect 25881 20417 25915 20451
rect 26157 20417 26191 20451
rect 26315 20417 26349 20451
rect 26433 20417 26467 20451
rect 26525 20417 26559 20451
rect 26617 20417 26651 20451
rect 26985 20417 27019 20451
rect 27261 20417 27295 20451
rect 27353 20417 27387 20451
rect 27629 20417 27663 20451
rect 28089 20417 28123 20451
rect 30297 20417 30331 20451
rect 30573 20417 30607 20451
rect 30941 20417 30975 20451
rect 31125 20417 31159 20451
rect 31309 20417 31343 20451
rect 34529 20417 34563 20451
rect 34805 20417 34839 20451
rect 5641 20349 5675 20383
rect 7297 20349 7331 20383
rect 8033 20349 8067 20383
rect 10149 20349 10183 20383
rect 11621 20349 11655 20383
rect 12541 20349 12575 20383
rect 14749 20349 14783 20383
rect 15025 20349 15059 20383
rect 15669 20349 15703 20383
rect 16773 20349 16807 20383
rect 25329 20349 25363 20383
rect 26801 20349 26835 20383
rect 27997 20349 28031 20383
rect 30389 20349 30423 20383
rect 31217 20349 31251 20383
rect 34621 20349 34655 20383
rect 21281 20281 21315 20315
rect 22845 20281 22879 20315
rect 27537 20281 27571 20315
rect 30757 20281 30791 20315
rect 6745 20213 6779 20247
rect 7205 20213 7239 20247
rect 7389 20213 7423 20247
rect 12173 20213 12207 20247
rect 13277 20213 13311 20247
rect 15117 20213 15151 20247
rect 16129 20213 16163 20247
rect 16313 20213 16347 20247
rect 16865 20213 16899 20247
rect 17049 20213 17083 20247
rect 17325 20213 17359 20247
rect 17509 20213 17543 20247
rect 21097 20213 21131 20247
rect 21833 20213 21867 20247
rect 26065 20213 26099 20247
rect 28457 20213 28491 20247
rect 30481 20213 30515 20247
rect 31401 20213 31435 20247
rect 31677 20213 31711 20247
rect 34529 20213 34563 20247
rect 4353 20009 4387 20043
rect 5181 20009 5215 20043
rect 6916 20009 6950 20043
rect 8401 20009 8435 20043
rect 8585 20009 8619 20043
rect 11437 20009 11471 20043
rect 13645 20009 13679 20043
rect 15945 20009 15979 20043
rect 16589 20009 16623 20043
rect 20545 20009 20579 20043
rect 26065 20009 26099 20043
rect 28365 20009 28399 20043
rect 29561 20009 29595 20043
rect 30021 20009 30055 20043
rect 33885 20009 33919 20043
rect 21741 19941 21775 19975
rect 5089 19873 5123 19907
rect 5917 19873 5951 19907
rect 6331 19873 6365 19907
rect 6653 19873 6687 19907
rect 9413 19873 9447 19907
rect 9689 19873 9723 19907
rect 11897 19873 11931 19907
rect 12173 19873 12207 19907
rect 14197 19873 14231 19907
rect 16129 19873 16163 19907
rect 16221 19873 16255 19907
rect 25697 19873 25731 19907
rect 29745 19873 29779 19907
rect 33977 19873 34011 19907
rect 1409 19805 1443 19839
rect 3801 19805 3835 19839
rect 3985 19805 4019 19839
rect 4169 19805 4203 19839
rect 5608 19805 5642 19839
rect 6193 19805 6227 19839
rect 8493 19805 8527 19839
rect 8677 19805 8711 19839
rect 9137 19805 9171 19839
rect 9229 19805 9263 19839
rect 9505 19805 9539 19839
rect 16313 19805 16347 19839
rect 16405 19805 16439 19839
rect 17233 19805 17267 19839
rect 18245 19805 18279 19839
rect 21097 19805 21131 19839
rect 21281 19805 21315 19839
rect 21373 19805 21407 19839
rect 21465 19805 21499 19839
rect 25881 19805 25915 19839
rect 27813 19805 27847 19839
rect 27997 19805 28031 19839
rect 28181 19805 28215 19839
rect 29837 19805 29871 19839
rect 34161 19805 34195 19839
rect 1685 19737 1719 19771
rect 4077 19737 4111 19771
rect 5825 19737 5859 19771
rect 9965 19737 9999 19771
rect 14473 19737 14507 19771
rect 16865 19737 16899 19771
rect 17049 19737 17083 19771
rect 18429 19737 18463 19771
rect 19257 19737 19291 19771
rect 28089 19737 28123 19771
rect 29561 19737 29595 19771
rect 33885 19737 33919 19771
rect 3157 19669 3191 19703
rect 5549 19669 5583 19703
rect 5733 19669 5767 19703
rect 6469 19669 6503 19703
rect 8953 19669 8987 19703
rect 18613 19669 18647 19703
rect 34345 19669 34379 19703
rect 2053 19465 2087 19499
rect 2513 19465 2547 19499
rect 10241 19465 10275 19499
rect 15878 19465 15912 19499
rect 18521 19465 18555 19499
rect 19165 19465 19199 19499
rect 19809 19465 19843 19499
rect 22477 19465 22511 19499
rect 23121 19465 23155 19499
rect 24409 19465 24443 19499
rect 33149 19465 33183 19499
rect 3801 19397 3835 19431
rect 5825 19397 5859 19431
rect 8585 19397 8619 19431
rect 9321 19397 9355 19431
rect 10701 19397 10735 19431
rect 12357 19397 12391 19431
rect 13645 19397 13679 19431
rect 19533 19397 19567 19431
rect 20177 19397 20211 19431
rect 23029 19397 23063 19431
rect 23489 19397 23523 19431
rect 25421 19397 25455 19431
rect 2421 19329 2455 19363
rect 2881 19329 2915 19363
rect 3433 19329 3467 19363
rect 3617 19329 3651 19363
rect 3893 19329 3927 19363
rect 3985 19329 4019 19363
rect 5457 19329 5491 19363
rect 6377 19329 6411 19363
rect 8217 19329 8251 19363
rect 8310 19329 8344 19363
rect 8493 19329 8527 19363
rect 8723 19329 8757 19363
rect 9224 19351 9258 19385
rect 9413 19329 9447 19363
rect 9551 19329 9585 19363
rect 10057 19329 10091 19363
rect 10609 19329 10643 19363
rect 11529 19329 11563 19363
rect 12081 19329 12115 19363
rect 12541 19329 12575 19363
rect 12725 19329 12759 19363
rect 13185 19329 13219 19363
rect 13461 19329 13495 19363
rect 14105 19329 14139 19363
rect 14381 19329 14415 19363
rect 14657 19329 14691 19363
rect 15485 19329 15519 19363
rect 15761 19329 15795 19363
rect 16313 19329 16347 19363
rect 17141 19329 17175 19363
rect 18521 19329 18555 19363
rect 18705 19329 18739 19363
rect 18981 19329 19015 19363
rect 19165 19329 19199 19363
rect 19257 19329 19291 19363
rect 19441 19329 19475 19363
rect 19625 19329 19659 19363
rect 19901 19329 19935 19363
rect 20085 19329 20119 19363
rect 20269 19329 20303 19363
rect 22661 19329 22695 19363
rect 22753 19329 22787 19363
rect 22937 19329 22971 19363
rect 24041 19329 24075 19363
rect 24133 19329 24167 19363
rect 24501 19329 24535 19363
rect 25237 19329 25271 19363
rect 25513 19329 25547 19363
rect 27905 19329 27939 19363
rect 28053 19329 28087 19363
rect 28181 19329 28215 19363
rect 28273 19329 28307 19363
rect 28411 19329 28445 19363
rect 32781 19329 32815 19363
rect 2605 19261 2639 19295
rect 5641 19261 5675 19295
rect 6653 19261 6687 19295
rect 8125 19261 8159 19295
rect 9321 19261 9355 19295
rect 9781 19261 9815 19295
rect 10885 19261 10919 19295
rect 13093 19261 13127 19295
rect 13921 19261 13955 19295
rect 14289 19261 14323 19295
rect 14473 19261 14507 19295
rect 16865 19261 16899 19295
rect 23305 19261 23339 19295
rect 23397 19261 23431 19295
rect 25053 19261 25087 19295
rect 32873 19261 32907 19295
rect 14381 19193 14415 19227
rect 4169 19125 4203 19159
rect 5733 19125 5767 19159
rect 8861 19125 8895 19159
rect 12817 19125 12851 19159
rect 13001 19125 13035 19159
rect 13737 19125 13771 19159
rect 20453 19125 20487 19159
rect 22661 19125 22695 19159
rect 24225 19125 24259 19159
rect 28549 19125 28583 19159
rect 32781 19125 32815 19159
rect 3157 18921 3191 18955
rect 4905 18921 4939 18955
rect 6745 18921 6779 18955
rect 10701 18921 10735 18955
rect 17049 18921 17083 18955
rect 21741 18921 21775 18955
rect 23121 18921 23155 18955
rect 24409 18921 24443 18955
rect 26525 18921 26559 18955
rect 30205 18921 30239 18955
rect 30665 18921 30699 18955
rect 34713 18921 34747 18955
rect 13277 18853 13311 18887
rect 18153 18853 18187 18887
rect 26157 18853 26191 18887
rect 7297 18785 7331 18819
rect 8309 18785 8343 18819
rect 8953 18785 8987 18819
rect 11437 18785 11471 18819
rect 16221 18785 16255 18819
rect 22845 18785 22879 18819
rect 26617 18785 26651 18819
rect 34805 18785 34839 18819
rect 1409 18717 1443 18751
rect 4353 18717 4387 18751
rect 4445 18717 4479 18751
rect 4629 18717 4663 18751
rect 4721 18717 4755 18751
rect 7205 18717 7239 18751
rect 8585 18717 8619 18751
rect 11713 18717 11747 18751
rect 11805 18717 11839 18751
rect 11989 18717 12023 18751
rect 12081 18717 12115 18751
rect 12357 18717 12391 18751
rect 12541 18717 12575 18751
rect 12817 18717 12851 18751
rect 13093 18717 13127 18751
rect 13277 18717 13311 18751
rect 13461 18717 13495 18751
rect 13553 18717 13587 18751
rect 14473 18717 14507 18751
rect 14749 18717 14783 18751
rect 15758 18717 15792 18751
rect 16129 18717 16163 18751
rect 17049 18717 17083 18751
rect 17417 18717 17451 18751
rect 17785 18717 17819 18751
rect 17969 18717 18003 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 21557 18717 21591 18751
rect 21925 18717 21959 18751
rect 22109 18717 22143 18751
rect 23305 18717 23339 18751
rect 23397 18717 23431 18751
rect 23489 18717 23523 18751
rect 23581 18717 23615 18751
rect 23949 18717 23983 18751
rect 24593 18717 24627 18751
rect 24685 18717 24719 18751
rect 24777 18717 24811 18751
rect 24869 18717 24903 18751
rect 25697 18717 25731 18751
rect 25789 18717 25823 18751
rect 25881 18717 25915 18751
rect 25973 18717 26007 18751
rect 26341 18717 26375 18751
rect 26709 18717 26743 18751
rect 26893 18717 26927 18751
rect 27537 18717 27571 18751
rect 27630 18717 27664 18751
rect 27813 18717 27847 18751
rect 28002 18717 28036 18751
rect 29561 18717 29595 18751
rect 29654 18717 29688 18751
rect 29837 18717 29871 18751
rect 30067 18717 30101 18751
rect 30849 18717 30883 18751
rect 31217 18717 31251 18751
rect 34713 18717 34747 18751
rect 34989 18717 35023 18751
rect 1685 18649 1719 18683
rect 7113 18649 7147 18683
rect 7665 18649 7699 18683
rect 9229 18649 9263 18683
rect 10793 18649 10827 18683
rect 12265 18649 12299 18683
rect 12725 18649 12759 18683
rect 14381 18649 14415 18683
rect 23765 18649 23799 18683
rect 24133 18649 24167 18683
rect 27905 18649 27939 18683
rect 29929 18649 29963 18683
rect 30941 18649 30975 18683
rect 31033 18649 31067 18683
rect 8677 18581 8711 18615
rect 12909 18581 12943 18615
rect 15577 18581 15611 18615
rect 15761 18581 15795 18615
rect 16865 18581 16899 18615
rect 21373 18581 21407 18615
rect 25513 18581 25547 18615
rect 27077 18581 27111 18615
rect 28181 18581 28215 18615
rect 35173 18581 35207 18615
rect 2053 18377 2087 18411
rect 7757 18377 7791 18411
rect 7849 18377 7883 18411
rect 8217 18377 8251 18411
rect 9045 18377 9079 18411
rect 9413 18377 9447 18411
rect 11253 18377 11287 18411
rect 13277 18377 13311 18411
rect 13829 18377 13863 18411
rect 20821 18377 20855 18411
rect 23029 18377 23063 18411
rect 24317 18377 24351 18411
rect 26065 18377 26099 18411
rect 27813 18377 27847 18411
rect 34069 18377 34103 18411
rect 35265 18377 35299 18411
rect 6837 18309 6871 18343
rect 9505 18309 9539 18343
rect 10057 18309 10091 18343
rect 10241 18309 10275 18343
rect 10609 18309 10643 18343
rect 10793 18309 10827 18343
rect 21005 18309 21039 18343
rect 23181 18309 23215 18343
rect 23397 18309 23431 18343
rect 24869 18309 24903 18343
rect 27445 18309 27479 18343
rect 32505 18309 32539 18343
rect 33701 18309 33735 18343
rect 35081 18309 35115 18343
rect 35357 18309 35391 18343
rect 2421 18241 2455 18275
rect 2881 18241 2915 18275
rect 3525 18241 3559 18275
rect 6745 18241 6779 18275
rect 7021 18241 7055 18275
rect 8401 18241 8435 18275
rect 8493 18241 8527 18275
rect 8677 18241 8711 18275
rect 8769 18241 8803 18275
rect 10333 18241 10367 18275
rect 11069 18241 11103 18275
rect 11345 18241 11379 18275
rect 12173 18241 12207 18275
rect 12541 18241 12575 18275
rect 12725 18241 12759 18275
rect 13001 18241 13035 18275
rect 13277 18241 13311 18275
rect 13461 18241 13495 18275
rect 13737 18241 13771 18275
rect 14013 18241 14047 18275
rect 21097 18241 21131 18275
rect 21281 18241 21315 18275
rect 21373 18241 21407 18275
rect 22201 18241 22235 18275
rect 23673 18241 23707 18275
rect 23857 18241 23891 18275
rect 23949 18241 23983 18275
rect 24041 18241 24075 18275
rect 24501 18241 24535 18275
rect 25421 18241 25455 18275
rect 25513 18241 25547 18275
rect 25697 18241 25731 18275
rect 25789 18241 25823 18275
rect 26157 18241 26191 18275
rect 27261 18241 27295 18275
rect 27537 18241 27571 18275
rect 27629 18241 27663 18275
rect 32275 18241 32309 18275
rect 32413 18241 32447 18275
rect 32688 18241 32722 18275
rect 32781 18241 32815 18275
rect 32965 18241 32999 18275
rect 33517 18241 33551 18275
rect 33793 18241 33827 18275
rect 33885 18241 33919 18275
rect 34897 18241 34931 18275
rect 35541 18241 35575 18275
rect 2513 18173 2547 18207
rect 2605 18173 2639 18207
rect 8033 18173 8067 18207
rect 9689 18173 9723 18207
rect 10885 18173 10919 18207
rect 11529 18173 11563 18207
rect 12265 18173 12299 18207
rect 13185 18173 13219 18207
rect 33241 18173 33275 18207
rect 7205 18105 7239 18139
rect 14013 18105 14047 18139
rect 21097 18105 21131 18139
rect 32137 18105 32171 18139
rect 7389 18037 7423 18071
rect 9873 18037 9907 18071
rect 10609 18037 10643 18071
rect 12817 18037 12851 18071
rect 20637 18037 20671 18071
rect 20821 18037 20855 18071
rect 23213 18037 23247 18071
rect 25237 18037 25271 18071
rect 35725 18037 35759 18071
rect 4445 17833 4479 17867
rect 7113 17833 7147 17867
rect 10149 17833 10183 17867
rect 11345 17833 11379 17867
rect 11713 17833 11747 17867
rect 12449 17833 12483 17867
rect 14105 17833 14139 17867
rect 14381 17833 14415 17867
rect 18705 17833 18739 17867
rect 22017 17833 22051 17867
rect 23673 17833 23707 17867
rect 30389 17833 30423 17867
rect 34345 17833 34379 17867
rect 34529 17833 34563 17867
rect 9229 17765 9263 17799
rect 20269 17765 20303 17799
rect 22753 17765 22787 17799
rect 23489 17765 23523 17799
rect 7757 17697 7791 17731
rect 8493 17697 8527 17731
rect 9321 17697 9355 17731
rect 14565 17697 14599 17731
rect 17233 17697 17267 17731
rect 30481 17697 30515 17731
rect 2605 17629 2639 17663
rect 2789 17629 2823 17663
rect 2973 17629 3007 17663
rect 3893 17629 3927 17663
rect 4261 17629 4295 17663
rect 4629 17629 4663 17663
rect 4721 17629 4755 17663
rect 4813 17629 4847 17663
rect 4905 17629 4939 17663
rect 5365 17629 5399 17663
rect 8953 17629 8987 17663
rect 9137 17629 9171 17663
rect 9413 17629 9447 17663
rect 9873 17629 9907 17663
rect 10057 17629 10091 17663
rect 10232 17623 10266 17657
rect 10333 17629 10367 17663
rect 10517 17629 10551 17663
rect 10885 17629 10919 17663
rect 11069 17629 11103 17663
rect 11892 17629 11926 17663
rect 12209 17629 12243 17663
rect 12357 17629 12391 17663
rect 12633 17629 12667 17663
rect 12817 17629 12851 17663
rect 14473 17629 14507 17663
rect 14841 17629 14875 17663
rect 15669 17629 15703 17663
rect 15761 17629 15795 17663
rect 15945 17629 15979 17663
rect 16037 17629 16071 17663
rect 17417 17629 17451 17663
rect 17509 17629 17543 17663
rect 17693 17629 17727 17663
rect 17785 17629 17819 17663
rect 18521 17629 18555 17663
rect 18797 17629 18831 17663
rect 20269 17629 20303 17663
rect 21005 17629 21039 17663
rect 21373 17629 21407 17663
rect 21465 17629 21499 17663
rect 22661 17629 22695 17663
rect 22845 17629 22879 17663
rect 22937 17629 22971 17663
rect 28825 17629 28859 17663
rect 29745 17629 29779 17663
rect 30113 17629 30147 17663
rect 30389 17629 30423 17663
rect 30665 17629 30699 17663
rect 34161 17629 34195 17663
rect 34253 17629 34287 17663
rect 21971 17595 22005 17629
rect 2881 17561 2915 17595
rect 4077 17561 4111 17595
rect 4169 17561 4203 17595
rect 5089 17561 5123 17595
rect 5641 17561 5675 17595
rect 8309 17561 8343 17595
rect 11161 17561 11195 17595
rect 11345 17561 11379 17595
rect 11989 17561 12023 17595
rect 12081 17561 12115 17595
rect 18061 17561 18095 17595
rect 18245 17561 18279 17595
rect 18337 17561 18371 17595
rect 22201 17561 22235 17595
rect 23857 17561 23891 17595
rect 29837 17561 29871 17595
rect 29929 17561 29963 17595
rect 3157 17493 3191 17527
rect 7205 17493 7239 17527
rect 7941 17493 7975 17527
rect 8401 17493 8435 17527
rect 9689 17493 9723 17527
rect 10517 17493 10551 17527
rect 10793 17493 10827 17527
rect 11529 17493 11563 17527
rect 14749 17493 14783 17527
rect 15485 17493 15519 17527
rect 17877 17493 17911 17527
rect 21833 17493 21867 17527
rect 23121 17493 23155 17527
rect 23657 17493 23691 17527
rect 29561 17493 29595 17527
rect 30205 17493 30239 17527
rect 3157 17289 3191 17323
rect 4537 17289 4571 17323
rect 6377 17289 6411 17323
rect 6745 17289 6779 17323
rect 9045 17289 9079 17323
rect 9965 17289 9999 17323
rect 11621 17289 11655 17323
rect 11989 17289 12023 17323
rect 12173 17289 12207 17323
rect 12633 17289 12667 17323
rect 15301 17289 15335 17323
rect 24961 17289 24995 17323
rect 27905 17289 27939 17323
rect 30757 17289 30791 17323
rect 31953 17289 31987 17323
rect 4169 17221 4203 17255
rect 7573 17221 7607 17255
rect 9505 17221 9539 17255
rect 17693 17221 17727 17255
rect 17877 17221 17911 17255
rect 27537 17221 27571 17255
rect 30297 17221 30331 17255
rect 3801 17153 3835 17187
rect 3985 17153 4019 17187
rect 4261 17153 4295 17187
rect 4353 17153 4387 17187
rect 4905 17153 4939 17187
rect 4997 17153 5031 17187
rect 5181 17153 5215 17187
rect 5457 17153 5491 17187
rect 5641 17153 5675 17187
rect 5825 17153 5859 17187
rect 5917 17153 5951 17187
rect 7297 17153 7331 17187
rect 9229 17153 9263 17187
rect 9321 17153 9355 17187
rect 9595 17153 9629 17187
rect 9721 17153 9755 17187
rect 10149 17153 10183 17187
rect 10333 17153 10367 17187
rect 11529 17153 11563 17187
rect 11805 17153 11839 17187
rect 12449 17153 12483 17187
rect 12725 17153 12759 17187
rect 15117 17153 15151 17187
rect 15393 17153 15427 17187
rect 16221 17153 16255 17187
rect 16313 17153 16347 17187
rect 19533 17153 19567 17187
rect 19809 17153 19843 17187
rect 20177 17153 20211 17187
rect 22109 17153 22143 17187
rect 22201 17153 22235 17187
rect 22293 17153 22327 17187
rect 22471 17153 22505 17187
rect 23397 17153 23431 17187
rect 25145 17153 25179 17187
rect 25237 17153 25271 17187
rect 25421 17153 25455 17187
rect 27353 17153 27387 17187
rect 27629 17153 27663 17187
rect 27721 17153 27755 17187
rect 27997 17153 28031 17187
rect 30573 17153 30607 17187
rect 31309 17153 31343 17187
rect 31457 17153 31491 17187
rect 31585 17153 31619 17187
rect 31677 17153 31711 17187
rect 31815 17153 31849 17187
rect 32137 17153 32171 17187
rect 32229 17153 32263 17187
rect 1409 17085 1443 17119
rect 1685 17085 1719 17119
rect 5089 17085 5123 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 10241 17085 10275 17119
rect 10425 17085 10459 17119
rect 12173 17085 12207 17119
rect 15853 17085 15887 17119
rect 16037 17085 16071 17119
rect 16129 17085 16163 17119
rect 19717 17085 19751 17119
rect 19993 17085 20027 17119
rect 20453 17085 20487 17119
rect 21833 17085 21867 17119
rect 28825 17085 28859 17119
rect 30481 17085 30515 17119
rect 3249 17017 3283 17051
rect 5365 17017 5399 17051
rect 12357 17017 12391 17051
rect 19625 17017 19659 17051
rect 20361 17017 20395 17051
rect 25329 17017 25363 17051
rect 9873 16949 9907 16983
rect 15117 16949 15151 16983
rect 19349 16949 19383 16983
rect 30389 16949 30423 16983
rect 32229 16949 32263 16983
rect 32505 16949 32539 16983
rect 1961 16745 1995 16779
rect 3157 16745 3191 16779
rect 6101 16745 6135 16779
rect 9781 16745 9815 16779
rect 10333 16745 10367 16779
rect 10701 16745 10735 16779
rect 12817 16745 12851 16779
rect 24409 16745 24443 16779
rect 25881 16745 25915 16779
rect 26985 16745 27019 16779
rect 2421 16609 2455 16643
rect 2513 16609 2547 16643
rect 4353 16609 4387 16643
rect 6561 16609 6595 16643
rect 6745 16609 6779 16643
rect 9505 16609 9539 16643
rect 10793 16609 10827 16643
rect 22661 16609 22695 16643
rect 26341 16609 26375 16643
rect 32045 16609 32079 16643
rect 32321 16609 32355 16643
rect 35173 16609 35207 16643
rect 35265 16609 35299 16643
rect 2329 16541 2363 16575
rect 3341 16541 3375 16575
rect 3617 16541 3651 16575
rect 4721 16541 4755 16575
rect 4997 16541 5031 16575
rect 5457 16541 5491 16575
rect 5825 16541 5859 16575
rect 7481 16541 7515 16575
rect 8493 16541 8527 16575
rect 8953 16541 8987 16575
rect 9045 16541 9079 16575
rect 9413 16541 9447 16575
rect 10517 16541 10551 16575
rect 11069 16541 11103 16575
rect 11621 16541 11655 16575
rect 11805 16541 11839 16575
rect 12633 16541 12667 16575
rect 12817 16541 12851 16575
rect 23489 16541 23523 16575
rect 24547 16541 24581 16575
rect 24905 16541 24939 16575
rect 25053 16541 25087 16575
rect 25513 16541 25547 16575
rect 25697 16541 25731 16575
rect 25973 16541 26007 16575
rect 26525 16541 26559 16575
rect 26617 16541 26651 16575
rect 26801 16541 26835 16575
rect 26893 16541 26927 16575
rect 27169 16541 27203 16575
rect 27261 16541 27295 16575
rect 27537 16541 27571 16575
rect 34069 16541 34103 16575
rect 35541 16541 35575 16575
rect 3525 16473 3559 16507
rect 4537 16473 4571 16507
rect 5641 16473 5675 16507
rect 5733 16473 5767 16507
rect 6469 16473 6503 16507
rect 6929 16473 6963 16507
rect 9229 16473 9263 16507
rect 9321 16473 9355 16507
rect 9689 16473 9723 16507
rect 10885 16473 10919 16507
rect 24685 16473 24719 16507
rect 24777 16473 24811 16507
rect 27353 16473 27387 16507
rect 28181 16473 28215 16507
rect 28917 16473 28951 16507
rect 3801 16405 3835 16439
rect 4905 16405 4939 16439
rect 6009 16405 6043 16439
rect 7941 16405 7975 16439
rect 3157 16201 3191 16235
rect 3617 16201 3651 16235
rect 3709 16201 3743 16235
rect 4905 16201 4939 16235
rect 5365 16201 5399 16235
rect 8217 16201 8251 16235
rect 9045 16201 9079 16235
rect 11345 16201 11379 16235
rect 17141 16201 17175 16235
rect 24593 16201 24627 16235
rect 29561 16201 29595 16235
rect 12265 16133 12299 16167
rect 14841 16133 14875 16167
rect 24225 16133 24259 16167
rect 24317 16133 24351 16167
rect 25881 16133 25915 16167
rect 27997 16133 28031 16167
rect 29193 16133 29227 16167
rect 34897 16133 34931 16167
rect 1409 16065 1443 16099
rect 6469 16065 6503 16099
rect 8953 16065 8987 16099
rect 11713 16065 11747 16099
rect 12081 16065 12115 16099
rect 12725 16065 12759 16099
rect 12909 16065 12943 16099
rect 13001 16065 13035 16099
rect 13185 16065 13219 16099
rect 13369 16065 13403 16099
rect 14019 16065 14053 16099
rect 14197 16065 14231 16099
rect 14473 16065 14507 16099
rect 14657 16065 14691 16099
rect 14749 16065 14783 16099
rect 14933 16065 14967 16099
rect 15209 16065 15243 16099
rect 17325 16065 17359 16099
rect 17601 16065 17635 16099
rect 22017 16065 22051 16099
rect 22293 16065 22327 16099
rect 22523 16065 22557 16099
rect 22707 16065 22741 16099
rect 23949 16065 23983 16099
rect 24042 16065 24076 16099
rect 24455 16065 24489 16099
rect 24869 16065 24903 16099
rect 24961 16065 24995 16099
rect 25145 16065 25179 16099
rect 25237 16065 25271 16099
rect 26065 16065 26099 16099
rect 27905 16065 27939 16099
rect 28089 16065 28123 16099
rect 28273 16065 28307 16099
rect 29009 16065 29043 16099
rect 29285 16065 29319 16099
rect 29377 16065 29411 16099
rect 31217 16065 31251 16099
rect 31401 16065 31435 16099
rect 34621 16065 34655 16099
rect 34805 16065 34839 16099
rect 34989 16065 35023 16099
rect 1685 15997 1719 16031
rect 3893 15997 3927 16031
rect 4997 15997 5031 16031
rect 5181 15997 5215 16031
rect 5917 15997 5951 16031
rect 6745 15997 6779 16031
rect 9229 15997 9263 16031
rect 9597 15997 9631 16031
rect 9873 15997 9907 16031
rect 13277 15997 13311 16031
rect 22201 15997 22235 16031
rect 22845 15997 22879 16031
rect 23397 15997 23431 16031
rect 3249 15929 3283 15963
rect 12817 15929 12851 15963
rect 17417 15929 17451 15963
rect 17509 15929 17543 15963
rect 4537 15861 4571 15895
rect 8585 15861 8619 15895
rect 12541 15861 12575 15895
rect 14105 15861 14139 15895
rect 14289 15861 14323 15895
rect 21833 15861 21867 15895
rect 22017 15861 22051 15895
rect 24685 15861 24719 15895
rect 25697 15861 25731 15895
rect 30941 15861 30975 15895
rect 31585 15861 31619 15895
rect 35173 15861 35207 15895
rect 3617 15657 3651 15691
rect 7113 15657 7147 15691
rect 7205 15657 7239 15691
rect 8033 15657 8067 15691
rect 9321 15657 9355 15691
rect 10609 15657 10643 15691
rect 16497 15657 16531 15691
rect 19349 15657 19383 15691
rect 19901 15657 19935 15691
rect 20269 15657 20303 15691
rect 20637 15657 20671 15691
rect 21373 15657 21407 15691
rect 31125 15657 31159 15691
rect 33149 15657 33183 15691
rect 33977 15657 34011 15691
rect 34713 15657 34747 15691
rect 34897 15657 34931 15691
rect 3801 15589 3835 15623
rect 12449 15589 12483 15623
rect 18613 15589 18647 15623
rect 18889 15589 18923 15623
rect 21189 15589 21223 15623
rect 23121 15589 23155 15623
rect 31861 15589 31895 15623
rect 1869 15521 1903 15555
rect 2145 15521 2179 15555
rect 4445 15521 4479 15555
rect 5181 15521 5215 15555
rect 5365 15521 5399 15555
rect 5641 15521 5675 15555
rect 7849 15521 7883 15555
rect 9873 15521 9907 15555
rect 11253 15521 11287 15555
rect 11989 15521 12023 15555
rect 12909 15521 12943 15555
rect 19533 15521 19567 15555
rect 19809 15521 19843 15555
rect 23581 15521 23615 15555
rect 30481 15521 30515 15555
rect 33057 15521 33091 15555
rect 33241 15521 33275 15555
rect 34161 15521 34195 15555
rect 34989 15521 35023 15555
rect 7573 15453 7607 15487
rect 7665 15453 7699 15487
rect 8217 15453 8251 15487
rect 8309 15453 8343 15487
rect 8585 15453 8619 15487
rect 9137 15453 9171 15487
rect 10057 15453 10091 15487
rect 10149 15453 10183 15487
rect 10517 15453 10551 15487
rect 12633 15453 12667 15487
rect 12817 15453 12851 15487
rect 14749 15453 14783 15487
rect 14842 15453 14876 15487
rect 15025 15453 15059 15487
rect 15255 15453 15289 15487
rect 15853 15453 15887 15487
rect 15946 15453 15980 15487
rect 16359 15453 16393 15487
rect 18889 15453 18923 15487
rect 19073 15453 19107 15487
rect 19257 15453 19291 15487
rect 19993 15453 20027 15487
rect 20085 15453 20119 15487
rect 20177 15453 20211 15487
rect 20453 15453 20487 15487
rect 21097 15453 21131 15487
rect 23029 15453 23063 15487
rect 23397 15453 23431 15487
rect 30639 15453 30673 15487
rect 30757 15453 30791 15487
rect 30941 15453 30975 15487
rect 31217 15453 31251 15487
rect 31310 15453 31344 15487
rect 31493 15453 31527 15487
rect 31682 15453 31716 15487
rect 32781 15453 32815 15487
rect 33425 15453 33459 15487
rect 34253 15453 34287 15487
rect 34897 15453 34931 15487
rect 35173 15453 35207 15487
rect 4169 15385 4203 15419
rect 4629 15385 4663 15419
rect 8401 15385 8435 15419
rect 10977 15385 11011 15419
rect 11437 15385 11471 15419
rect 15117 15385 15151 15419
rect 16129 15385 16163 15419
rect 16221 15385 16255 15419
rect 19533 15385 19567 15419
rect 20729 15385 20763 15419
rect 20913 15385 20947 15419
rect 21341 15385 21375 15419
rect 21557 15385 21591 15419
rect 30849 15385 30883 15419
rect 31585 15385 31619 15419
rect 33149 15385 33183 15419
rect 33977 15385 34011 15419
rect 4261 15317 4295 15351
rect 9045 15317 9079 15351
rect 10241 15317 10275 15351
rect 11069 15317 11103 15351
rect 15393 15317 15427 15351
rect 33609 15317 33643 15351
rect 34437 15317 34471 15351
rect 5549 15113 5583 15147
rect 15577 15113 15611 15147
rect 17785 15113 17819 15147
rect 19257 15113 19291 15147
rect 23765 15113 23799 15147
rect 24961 15113 24995 15147
rect 32781 15113 32815 15147
rect 4077 15045 4111 15079
rect 8125 15045 8159 15079
rect 15025 15045 15059 15079
rect 20269 15045 20303 15079
rect 20453 15045 20487 15079
rect 32413 15045 32447 15079
rect 32505 15045 32539 15079
rect 1961 14977 1995 15011
rect 3801 14977 3835 15011
rect 5825 14977 5859 15011
rect 6377 14977 6411 15011
rect 6561 14977 6595 15011
rect 6653 14977 6687 15011
rect 6837 14977 6871 15011
rect 7481 14977 7515 15011
rect 7665 14977 7699 15011
rect 7849 14977 7883 15011
rect 9873 14977 9907 15011
rect 10149 14977 10183 15011
rect 10333 14977 10367 15011
rect 10517 14977 10551 15011
rect 10701 14977 10735 15011
rect 10793 14977 10827 15011
rect 10977 14977 11011 15011
rect 15301 14977 15335 15011
rect 15393 14977 15427 15011
rect 15669 14977 15703 15011
rect 19349 14977 19383 15011
rect 20545 14977 20579 15011
rect 23949 14977 23983 15011
rect 25053 14977 25087 15011
rect 27537 14977 27571 15011
rect 27721 14977 27755 15011
rect 32137 14977 32171 15011
rect 32295 14977 32329 15011
rect 32597 14977 32631 15011
rect 2237 14909 2271 14943
rect 5641 14909 5675 14943
rect 9597 14909 9631 14943
rect 9689 14909 9723 14943
rect 10057 14909 10091 14943
rect 17969 14909 18003 14943
rect 18061 14909 18095 14943
rect 18153 14909 18187 14943
rect 18245 14909 18279 14943
rect 24225 14909 24259 14943
rect 24777 14909 24811 14943
rect 3709 14841 3743 14875
rect 9965 14841 9999 14875
rect 20269 14841 20303 14875
rect 24133 14841 24167 14875
rect 6009 14773 6043 14807
rect 6561 14773 6595 14807
rect 6653 14773 6687 14807
rect 7573 14773 7607 14807
rect 11161 14773 11195 14807
rect 15393 14773 15427 14807
rect 24317 14773 24351 14807
rect 24593 14773 24627 14807
rect 24685 14773 24719 14807
rect 27537 14773 27571 14807
rect 27905 14773 27939 14807
rect 3801 14569 3835 14603
rect 9229 14569 9263 14603
rect 9413 14569 9447 14603
rect 23305 14569 23339 14603
rect 25053 14569 25087 14603
rect 26249 14569 26283 14603
rect 27445 14569 27479 14603
rect 30297 14569 30331 14603
rect 33793 14569 33827 14603
rect 3617 14501 3651 14535
rect 7849 14501 7883 14535
rect 25421 14501 25455 14535
rect 25973 14501 26007 14535
rect 1869 14433 1903 14467
rect 4261 14433 4295 14467
rect 4445 14433 4479 14467
rect 6561 14433 6595 14467
rect 7389 14433 7423 14467
rect 8677 14433 8711 14467
rect 9965 14433 9999 14467
rect 10057 14433 10091 14467
rect 10793 14433 10827 14467
rect 10977 14433 11011 14467
rect 20545 14433 20579 14467
rect 23489 14433 23523 14467
rect 25329 14433 25363 14467
rect 27813 14433 27847 14467
rect 28181 14433 28215 14467
rect 33885 14433 33919 14467
rect 5181 14365 5215 14399
rect 5733 14365 5767 14399
rect 7757 14365 7791 14399
rect 8401 14365 8435 14399
rect 11161 14365 11195 14399
rect 11253 14365 11287 14399
rect 11529 14365 11563 14399
rect 13093 14365 13127 14399
rect 13277 14365 13311 14399
rect 13369 14365 13403 14399
rect 13553 14365 13587 14399
rect 13645 14365 13679 14399
rect 17785 14365 17819 14399
rect 17969 14365 18003 14399
rect 18061 14365 18095 14399
rect 19901 14365 19935 14399
rect 19993 14365 20027 14399
rect 20269 14365 20303 14399
rect 20453 14365 20487 14399
rect 20729 14365 20763 14399
rect 20821 14365 20855 14399
rect 21005 14365 21039 14399
rect 21097 14365 21131 14399
rect 23397 14365 23431 14399
rect 23581 14365 23615 14399
rect 23765 14365 23799 14399
rect 25237 14365 25271 14399
rect 25513 14365 25547 14399
rect 25789 14365 25823 14399
rect 25881 14365 25915 14399
rect 26065 14365 26099 14399
rect 26525 14365 26559 14399
rect 26709 14365 26743 14399
rect 26985 14365 27019 14399
rect 27353 14365 27387 14399
rect 27629 14365 27663 14399
rect 27721 14365 27755 14399
rect 27905 14365 27939 14399
rect 29653 14365 29687 14399
rect 29801 14365 29835 14399
rect 30159 14365 30193 14399
rect 34069 14365 34103 14399
rect 2145 14297 2179 14331
rect 4169 14297 4203 14331
rect 4629 14297 4663 14331
rect 5549 14297 5583 14331
rect 6285 14297 6319 14331
rect 7205 14297 7239 14331
rect 9045 14297 9079 14331
rect 9873 14297 9907 14331
rect 19257 14297 19291 14331
rect 23029 14297 23063 14331
rect 28457 14297 28491 14331
rect 29929 14297 29963 14331
rect 30021 14297 30055 14331
rect 33793 14297 33827 14331
rect 5365 14229 5399 14263
rect 5917 14229 5951 14263
rect 6377 14229 6411 14263
rect 6837 14229 6871 14263
rect 7297 14229 7331 14263
rect 8033 14229 8067 14263
rect 8493 14229 8527 14263
rect 9250 14229 9284 14263
rect 9505 14229 9539 14263
rect 10333 14229 10367 14263
rect 10701 14229 10735 14263
rect 17601 14229 17635 14263
rect 26893 14229 26927 14263
rect 27169 14229 27203 14263
rect 34253 14229 34287 14263
rect 3249 14025 3283 14059
rect 3709 14025 3743 14059
rect 5917 14025 5951 14059
rect 6745 14025 6779 14059
rect 6929 14025 6963 14059
rect 7389 14025 7423 14059
rect 7941 14025 7975 14059
rect 8309 14025 8343 14059
rect 8401 14025 8435 14059
rect 11345 14025 11379 14059
rect 13921 14025 13955 14059
rect 15853 14025 15887 14059
rect 21373 14025 21407 14059
rect 25605 14025 25639 14059
rect 26157 14025 26191 14059
rect 27629 14025 27663 14059
rect 28365 14025 28399 14059
rect 31677 14025 31711 14059
rect 32873 14025 32907 14059
rect 33609 14025 33643 14059
rect 35357 14025 35391 14059
rect 35817 14025 35851 14059
rect 12265 13957 12299 13991
rect 14381 13957 14415 13991
rect 16681 13957 16715 13991
rect 22109 13957 22143 13991
rect 25145 13957 25179 13991
rect 26341 13957 26375 13991
rect 27261 13957 27295 13991
rect 27477 13957 27511 13991
rect 28733 13957 28767 13991
rect 31309 13957 31343 13991
rect 34897 13957 34931 13991
rect 1409 13889 1443 13923
rect 3617 13889 3651 13923
rect 4077 13889 4111 13923
rect 4721 13889 4755 13923
rect 4813 13889 4847 13923
rect 4997 13889 5031 13923
rect 5181 13889 5215 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 6561 13889 6595 13923
rect 6837 13889 6871 13923
rect 7297 13889 7331 13923
rect 8769 13889 8803 13923
rect 8953 13889 8987 13923
rect 9229 13889 9263 13923
rect 9505 13889 9539 13923
rect 9597 13889 9631 13923
rect 12081 13889 12115 13923
rect 12449 13889 12483 13923
rect 14105 13889 14139 13923
rect 16037 13889 16071 13923
rect 16313 13889 16347 13923
rect 16865 13889 16899 13923
rect 16957 13889 16991 13923
rect 17141 13889 17175 13923
rect 17233 13889 17267 13923
rect 21189 13889 21223 13923
rect 21465 13889 21499 13923
rect 22569 13889 22603 13923
rect 22753 13889 22787 13923
rect 22845 13889 22879 13923
rect 23029 13889 23063 13923
rect 24225 13889 24259 13923
rect 24409 13889 24443 13923
rect 24501 13889 24535 13923
rect 25421 13889 25455 13923
rect 26525 13889 26559 13923
rect 28549 13889 28583 13923
rect 28641 13889 28675 13923
rect 28917 13889 28951 13923
rect 29009 13889 29043 13923
rect 31033 13889 31067 13923
rect 31126 13889 31160 13923
rect 31401 13889 31435 13923
rect 31539 13889 31573 13923
rect 32413 13889 32447 13923
rect 32689 13889 32723 13923
rect 33793 13889 33827 13923
rect 34069 13889 34103 13923
rect 35081 13889 35115 13923
rect 35173 13889 35207 13923
rect 35449 13889 35483 13923
rect 1685 13821 1719 13855
rect 3893 13821 3927 13855
rect 6377 13821 6411 13855
rect 7481 13821 7515 13855
rect 8493 13821 8527 13855
rect 9873 13821 9907 13855
rect 12633 13821 12667 13855
rect 14197 13821 14231 13855
rect 16129 13821 16163 13855
rect 21005 13821 21039 13855
rect 25237 13821 25271 13855
rect 32505 13821 32539 13855
rect 33885 13821 33919 13855
rect 35541 13821 35575 13855
rect 3157 13753 3191 13787
rect 5457 13753 5491 13787
rect 24041 13753 24075 13787
rect 5825 13685 5859 13719
rect 8861 13685 8895 13719
rect 9413 13685 9447 13719
rect 11529 13685 11563 13719
rect 14381 13685 14415 13719
rect 16313 13685 16347 13719
rect 25421 13685 25455 13719
rect 27445 13685 27479 13719
rect 32689 13685 32723 13719
rect 33793 13685 33827 13719
rect 34897 13685 34931 13719
rect 35449 13685 35483 13719
rect 2421 13481 2455 13515
rect 4445 13481 4479 13515
rect 4997 13481 5031 13515
rect 5549 13481 5583 13515
rect 9965 13481 9999 13515
rect 12725 13481 12759 13515
rect 14749 13481 14783 13515
rect 16589 13481 16623 13515
rect 20269 13481 20303 13515
rect 26433 13481 26467 13515
rect 29561 13481 29595 13515
rect 30297 13481 30331 13515
rect 33149 13481 33183 13515
rect 4813 13413 4847 13447
rect 6837 13413 6871 13447
rect 16957 13413 16991 13447
rect 19533 13413 19567 13447
rect 19625 13413 19659 13447
rect 20085 13413 20119 13447
rect 26249 13413 26283 13447
rect 2881 13345 2915 13379
rect 3065 13345 3099 13379
rect 5365 13345 5399 13379
rect 7389 13345 7423 13379
rect 9321 13345 9355 13379
rect 9597 13345 9631 13379
rect 14657 13345 14691 13379
rect 16037 13345 16071 13379
rect 17785 13345 17819 13379
rect 19717 13345 19751 13379
rect 29745 13345 29779 13379
rect 29837 13345 29871 13379
rect 30021 13345 30055 13379
rect 32505 13345 32539 13379
rect 4445 13277 4479 13311
rect 4721 13277 4755 13311
rect 5641 13277 5675 13311
rect 5917 13277 5951 13311
rect 6101 13277 6135 13311
rect 6285 13277 6319 13311
rect 6377 13277 6411 13311
rect 6561 13277 6595 13311
rect 7297 13277 7331 13311
rect 8033 13277 8067 13311
rect 8309 13277 8343 13311
rect 8493 13277 8527 13311
rect 9229 13277 9263 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 10517 13277 10551 13311
rect 10609 13277 10643 13311
rect 10793 13277 10827 13311
rect 12725 13277 12759 13311
rect 12817 13277 12851 13311
rect 14473 13277 14507 13311
rect 14749 13277 14783 13311
rect 16221 13277 16255 13311
rect 16497 13277 16531 13311
rect 16773 13277 16807 13311
rect 17049 13277 17083 13311
rect 17601 13277 17635 13311
rect 17693 13277 17727 13311
rect 17877 13277 17911 13311
rect 19993 13277 20027 13311
rect 20269 13277 20303 13311
rect 20361 13277 20395 13311
rect 29929 13277 29963 13311
rect 30481 13277 30515 13311
rect 30849 13277 30883 13311
rect 32643 13277 32677 13311
rect 32965 13277 32999 13311
rect 2789 13209 2823 13243
rect 3985 13209 4019 13243
rect 4169 13209 4203 13243
rect 5181 13209 5215 13243
rect 7849 13209 7883 13243
rect 8401 13209 8435 13243
rect 10333 13209 10367 13243
rect 13001 13209 13035 13243
rect 16405 13209 16439 13243
rect 20545 13209 20579 13243
rect 26617 13209 26651 13243
rect 30573 13209 30607 13243
rect 30665 13209 30699 13243
rect 32781 13209 32815 13243
rect 32873 13209 32907 13243
rect 3801 13141 3835 13175
rect 4629 13141 4663 13175
rect 4981 13141 5015 13175
rect 5365 13141 5399 13175
rect 6469 13141 6503 13175
rect 7205 13141 7239 13175
rect 8217 13141 8251 13175
rect 10609 13141 10643 13175
rect 12541 13141 12575 13175
rect 14933 13141 14967 13175
rect 17417 13141 17451 13175
rect 19257 13141 19291 13175
rect 19901 13141 19935 13175
rect 26433 13141 26467 13175
rect 3157 12937 3191 12971
rect 3249 12937 3283 12971
rect 5825 12937 5859 12971
rect 7021 12937 7055 12971
rect 8861 12937 8895 12971
rect 9689 12937 9723 12971
rect 14289 12937 14323 12971
rect 19533 12937 19567 12971
rect 22293 12937 22327 12971
rect 4353 12869 4387 12903
rect 4537 12869 4571 12903
rect 9045 12869 9079 12903
rect 10149 12869 10183 12903
rect 14749 12869 14783 12903
rect 22845 12869 22879 12903
rect 23045 12869 23079 12903
rect 3617 12801 3651 12835
rect 4169 12801 4203 12835
rect 4808 12801 4842 12835
rect 4905 12801 4939 12835
rect 4997 12801 5031 12835
rect 5180 12801 5214 12835
rect 5273 12801 5307 12835
rect 5435 12801 5469 12835
rect 5733 12801 5767 12835
rect 5825 12801 5859 12835
rect 6009 12801 6043 12835
rect 6929 12801 6963 12835
rect 7573 12801 7607 12835
rect 8217 12801 8251 12835
rect 8309 12801 8343 12835
rect 8401 12801 8435 12835
rect 8585 12801 8619 12835
rect 8677 12801 8711 12835
rect 9321 12801 9355 12835
rect 9965 12801 9999 12835
rect 10241 12801 10275 12835
rect 14473 12801 14507 12835
rect 15025 12801 15059 12835
rect 15577 12801 15611 12835
rect 19717 12801 19751 12835
rect 19901 12801 19935 12835
rect 21833 12801 21867 12835
rect 22017 12801 22051 12835
rect 22109 12801 22143 12835
rect 24041 12801 24075 12835
rect 1409 12733 1443 12767
rect 1685 12733 1719 12767
rect 3709 12733 3743 12767
rect 3893 12733 3927 12767
rect 5549 12733 5583 12767
rect 7113 12733 7147 12767
rect 7849 12733 7883 12767
rect 7941 12733 7975 12767
rect 9229 12733 9263 12767
rect 10333 12733 10367 12767
rect 10609 12733 10643 12767
rect 14565 12733 14599 12767
rect 15761 12733 15795 12767
rect 5365 12665 5399 12699
rect 15025 12665 15059 12699
rect 4629 12597 4663 12631
rect 5641 12597 5675 12631
rect 6561 12597 6595 12631
rect 7389 12597 7423 12631
rect 7757 12597 7791 12631
rect 9781 12597 9815 12631
rect 14657 12597 14691 12631
rect 19901 12597 19935 12631
rect 21833 12597 21867 12631
rect 23029 12597 23063 12631
rect 23213 12597 23247 12631
rect 23949 12597 23983 12631
rect 2513 12393 2547 12427
rect 3801 12393 3835 12427
rect 8585 12393 8619 12427
rect 8769 12393 8803 12427
rect 10333 12393 10367 12427
rect 10609 12393 10643 12427
rect 13093 12393 13127 12427
rect 15393 12393 15427 12427
rect 17509 12393 17543 12427
rect 18613 12393 18647 12427
rect 18797 12393 18831 12427
rect 21649 12393 21683 12427
rect 23857 12393 23891 12427
rect 24041 12393 24075 12427
rect 24777 12393 24811 12427
rect 25789 12393 25823 12427
rect 27629 12393 27663 12427
rect 28089 12393 28123 12427
rect 30205 12393 30239 12427
rect 31217 12393 31251 12427
rect 32781 12393 32815 12427
rect 34529 12393 34563 12427
rect 35357 12393 35391 12427
rect 4721 12325 4755 12359
rect 7389 12325 7423 12359
rect 8217 12325 8251 12359
rect 10517 12325 10551 12359
rect 14105 12325 14139 12359
rect 17693 12325 17727 12359
rect 18153 12325 18187 12359
rect 22753 12325 22787 12359
rect 23305 12325 23339 12359
rect 25145 12325 25179 12359
rect 2145 12257 2179 12291
rect 3985 12257 4019 12291
rect 4169 12257 4203 12291
rect 4261 12257 4295 12291
rect 5181 12257 5215 12291
rect 5733 12257 5767 12291
rect 5917 12257 5951 12291
rect 6009 12257 6043 12291
rect 6193 12257 6227 12291
rect 6469 12257 6503 12291
rect 7205 12257 7239 12291
rect 10977 12257 11011 12291
rect 15301 12257 15335 12291
rect 18337 12257 18371 12291
rect 21189 12257 21223 12291
rect 21281 12257 21315 12291
rect 26985 12257 27019 12291
rect 29561 12257 29595 12291
rect 2053 12189 2087 12223
rect 2692 12189 2726 12223
rect 2789 12189 2823 12223
rect 3064 12189 3098 12223
rect 3157 12189 3191 12223
rect 3433 12189 3467 12223
rect 3617 12189 3651 12223
rect 4077 12189 4111 12223
rect 4445 12189 4479 12223
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 5273 12189 5307 12223
rect 5365 12189 5399 12223
rect 5825 12189 5859 12223
rect 6561 12189 6595 12223
rect 7481 12189 7515 12223
rect 7757 12189 7791 12223
rect 7849 12189 7883 12223
rect 7941 12189 7975 12223
rect 8033 12189 8067 12223
rect 9137 12189 9171 12223
rect 9321 12189 9355 12223
rect 9413 12189 9447 12223
rect 9505 12189 9539 12223
rect 9689 12189 9723 12223
rect 9873 12189 9907 12223
rect 9965 12189 9999 12223
rect 10333 12189 10367 12223
rect 10793 12189 10827 12223
rect 11621 12189 11655 12223
rect 11815 12189 11849 12223
rect 13001 12189 13035 12223
rect 13093 12189 13127 12223
rect 14657 12189 14691 12223
rect 15209 12189 15243 12223
rect 15485 12189 15519 12223
rect 17785 12189 17819 12223
rect 18061 12189 18095 12223
rect 18245 12189 18279 12223
rect 18521 12189 18555 12223
rect 21465 12189 21499 12223
rect 22109 12189 22143 12223
rect 22385 12189 22419 12223
rect 22937 12189 22971 12223
rect 24409 12189 24443 12223
rect 24961 12189 24995 12223
rect 25053 12189 25087 12223
rect 25237 12189 25271 12223
rect 25421 12189 25455 12223
rect 26801 12189 26835 12223
rect 27169 12189 27203 12223
rect 27537 12189 27571 12223
rect 27813 12189 27847 12223
rect 27905 12189 27939 12223
rect 28273 12189 28307 12223
rect 28457 12189 28491 12223
rect 29929 12189 29963 12223
rect 30021 12189 30055 12223
rect 30573 12189 30607 12223
rect 30721 12189 30755 12223
rect 30941 12189 30975 12223
rect 31038 12189 31072 12223
rect 32413 12189 32447 12223
rect 32597 12189 32631 12223
rect 33977 12189 34011 12223
rect 34253 12189 34287 12223
rect 34345 12189 34379 12223
rect 34713 12189 34747 12223
rect 34851 12189 34885 12223
rect 35173 12189 35207 12223
rect 23903 12155 23937 12189
rect 2881 12121 2915 12155
rect 3525 12121 3559 12155
rect 6837 12121 6871 12155
rect 6929 12121 6963 12155
rect 8585 12121 8619 12155
rect 11713 12121 11747 12155
rect 14289 12121 14323 12155
rect 17325 12121 17359 12155
rect 18981 12121 19015 12155
rect 23673 12121 23707 12155
rect 25605 12121 25639 12155
rect 29699 12121 29733 12155
rect 29837 12121 29871 12155
rect 30849 12121 30883 12155
rect 34161 12121 34195 12155
rect 34989 12121 35023 12155
rect 35081 12121 35115 12155
rect 2421 12053 2455 12087
rect 4997 12053 5031 12087
rect 6285 12053 6319 12087
rect 7481 12053 7515 12087
rect 7573 12053 7607 12087
rect 12725 12053 12759 12087
rect 14381 12053 14415 12087
rect 14473 12053 14507 12087
rect 15025 12053 15059 12087
rect 17535 12053 17569 12087
rect 18781 12053 18815 12087
rect 21925 12053 21959 12087
rect 22293 12053 22327 12087
rect 23029 12053 23063 12087
rect 23121 12053 23155 12087
rect 24593 12053 24627 12087
rect 2421 11849 2455 11883
rect 2973 11849 3007 11883
rect 4445 11849 4479 11883
rect 5917 11849 5951 11883
rect 6009 11849 6043 11883
rect 6469 11849 6503 11883
rect 9137 11849 9171 11883
rect 9873 11849 9907 11883
rect 10057 11849 10091 11883
rect 10977 11849 11011 11883
rect 16681 11849 16715 11883
rect 23121 11849 23155 11883
rect 26709 11849 26743 11883
rect 30757 11849 30791 11883
rect 31493 11849 31527 11883
rect 31861 11849 31895 11883
rect 17417 11781 17451 11815
rect 28273 11781 28307 11815
rect 30481 11781 30515 11815
rect 32965 11781 32999 11815
rect 2635 11713 2669 11747
rect 2789 11713 2823 11747
rect 2881 11713 2915 11747
rect 3065 11713 3099 11747
rect 4537 11713 4571 11747
rect 4905 11713 4939 11747
rect 4997 11713 5031 11747
rect 5273 11713 5307 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 6009 11713 6043 11747
rect 6193 11713 6227 11747
rect 6648 11713 6682 11747
rect 6745 11713 6779 11747
rect 6837 11713 6871 11747
rect 6965 11713 6999 11747
rect 7113 11713 7147 11747
rect 7205 11713 7239 11747
rect 7389 11713 7423 11747
rect 7481 11713 7515 11747
rect 7665 11713 7699 11747
rect 7757 11713 7791 11747
rect 7941 11713 7975 11747
rect 8309 11713 8343 11747
rect 8401 11713 8435 11747
rect 8493 11713 8527 11747
rect 8677 11713 8711 11747
rect 8769 11713 8803 11747
rect 8923 11713 8957 11747
rect 9689 11713 9723 11747
rect 9968 11713 10002 11747
rect 10241 11713 10275 11747
rect 10701 11713 10735 11747
rect 11161 11713 11195 11747
rect 11253 11713 11287 11747
rect 11713 11713 11747 11747
rect 12265 11713 12299 11747
rect 13001 11713 13035 11747
rect 13277 11713 13311 11747
rect 15393 11713 15427 11747
rect 15577 11713 15611 11747
rect 16865 11713 16899 11747
rect 17325 11713 17359 11747
rect 17601 11713 17635 11747
rect 17693 11713 17727 11747
rect 17877 11713 17911 11747
rect 17969 11713 18003 11747
rect 20361 11713 20395 11747
rect 20545 11713 20579 11747
rect 20637 11713 20671 11747
rect 20729 11713 20763 11747
rect 23305 11713 23339 11747
rect 26617 11713 26651 11747
rect 26801 11713 26835 11747
rect 27261 11713 27295 11747
rect 27445 11713 27479 11747
rect 27721 11713 27755 11747
rect 29193 11713 29227 11747
rect 30113 11713 30147 11747
rect 30271 11713 30305 11747
rect 30389 11713 30423 11747
rect 30573 11713 30607 11747
rect 31309 11713 31343 11747
rect 31677 11713 31711 11747
rect 32321 11713 32355 11747
rect 32689 11713 32723 11747
rect 4721 11645 4755 11679
rect 4813 11645 4847 11679
rect 9229 11645 9263 11679
rect 10425 11645 10459 11679
rect 11529 11645 11563 11679
rect 12541 11645 12575 11679
rect 17049 11645 17083 11679
rect 27353 11645 27387 11679
rect 35817 11645 35851 11679
rect 36093 11645 36127 11679
rect 7205 11577 7239 11611
rect 7481 11577 7515 11611
rect 7757 11577 7791 11611
rect 9597 11577 9631 11611
rect 12725 11577 12759 11611
rect 26985 11577 27019 11611
rect 28089 11577 28123 11611
rect 5181 11509 5215 11543
rect 8033 11509 8067 11543
rect 9505 11509 9539 11543
rect 10609 11509 10643 11543
rect 12909 11509 12943 11543
rect 15209 11509 15243 11543
rect 16865 11509 16899 11543
rect 21005 11509 21039 11543
rect 27537 11509 27571 11543
rect 28917 11509 28951 11543
rect 33057 11509 33091 11543
rect 34345 11509 34379 11543
rect 2329 11305 2363 11339
rect 3065 11305 3099 11339
rect 11805 11305 11839 11339
rect 12357 11305 12391 11339
rect 12541 11305 12575 11339
rect 12909 11305 12943 11339
rect 17141 11305 17175 11339
rect 19441 11305 19475 11339
rect 19625 11305 19659 11339
rect 23213 11305 23247 11339
rect 23489 11305 23523 11339
rect 27629 11305 27663 11339
rect 31585 11305 31619 11339
rect 32597 11305 32631 11339
rect 33241 11305 33275 11339
rect 34897 11305 34931 11339
rect 4721 11237 4755 11271
rect 5733 11237 5767 11271
rect 17233 11237 17267 11271
rect 29929 11237 29963 11271
rect 31401 11237 31435 11271
rect 32689 11237 32723 11271
rect 2053 11169 2087 11203
rect 3801 11169 3835 11203
rect 5917 11169 5951 11203
rect 7389 11169 7423 11203
rect 8585 11169 8619 11203
rect 8953 11169 8987 11203
rect 16773 11169 16807 11203
rect 27905 11169 27939 11203
rect 31953 11169 31987 11203
rect 35081 11169 35115 11203
rect 1961 11101 1995 11135
rect 2421 11101 2455 11135
rect 2605 11101 2639 11135
rect 2697 11101 2731 11135
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 3065 11101 3099 11135
rect 3249 11101 3283 11135
rect 3985 11101 4019 11135
rect 4169 11101 4203 11135
rect 4261 11101 4295 11135
rect 4905 11101 4939 11135
rect 4998 11101 5032 11135
rect 5273 11101 5307 11135
rect 5411 11101 5445 11135
rect 5825 11101 5859 11135
rect 6101 11101 6135 11135
rect 6377 11101 6411 11135
rect 6469 11101 6503 11135
rect 7113 11101 7147 11135
rect 8493 11101 8527 11135
rect 9965 11101 9999 11135
rect 10149 11101 10183 11135
rect 10333 11101 10367 11135
rect 10609 11101 10643 11135
rect 10885 11101 10919 11135
rect 10977 11101 11011 11135
rect 11989 11101 12023 11135
rect 12173 11101 12207 11135
rect 12817 11101 12851 11135
rect 13093 11101 13127 11135
rect 14381 11101 14415 11135
rect 14565 11101 14599 11135
rect 14657 11101 14691 11135
rect 14841 11101 14875 11135
rect 14933 11101 14967 11135
rect 16957 11101 16991 11135
rect 17509 11101 17543 11135
rect 18429 11101 18463 11135
rect 19257 11101 19291 11135
rect 19441 11101 19475 11135
rect 22661 11101 22695 11135
rect 22753 11101 22787 11135
rect 22937 11101 22971 11135
rect 23029 11101 23063 11135
rect 27445 11101 27479 11135
rect 27629 11101 27663 11135
rect 27997 11101 28031 11135
rect 28181 11101 28215 11135
rect 28365 11101 28399 11135
rect 28917 11101 28951 11135
rect 29009 11101 29043 11135
rect 29101 11101 29135 11135
rect 29193 11101 29227 11135
rect 29561 11101 29595 11135
rect 30113 11101 30147 11135
rect 32091 11101 32125 11135
rect 32229 11101 32263 11135
rect 32321 11101 32355 11135
rect 32413 11101 32447 11135
rect 34805 11101 34839 11135
rect 35357 11101 35391 11135
rect 4353 11033 4387 11067
rect 5181 11033 5215 11067
rect 6285 11033 6319 11067
rect 7665 11033 7699 11067
rect 12449 11033 12483 11067
rect 17233 11033 17267 11067
rect 23673 11033 23707 11067
rect 24409 11033 24443 11067
rect 24593 11033 24627 11067
rect 28273 11033 28307 11067
rect 28641 11033 28675 11067
rect 31569 11033 31603 11067
rect 31769 11033 31803 11067
rect 32965 11033 32999 11067
rect 33057 11033 33091 11067
rect 3433 10965 3467 10999
rect 4813 10965 4847 10999
rect 5549 10965 5583 10999
rect 10241 10965 10275 10999
rect 17417 10965 17451 10999
rect 18245 10965 18279 10999
rect 23305 10965 23339 10999
rect 23473 10965 23507 10999
rect 28733 10965 28767 10999
rect 29745 10965 29779 10999
rect 32873 10965 32907 10999
rect 3157 10761 3191 10795
rect 7941 10761 7975 10795
rect 10517 10761 10551 10795
rect 15025 10761 15059 10795
rect 21649 10761 21683 10795
rect 24041 10761 24075 10795
rect 24225 10761 24259 10795
rect 25237 10761 25271 10795
rect 27905 10761 27939 10795
rect 29377 10761 29411 10795
rect 29469 10761 29503 10795
rect 29653 10761 29687 10795
rect 30205 10761 30239 10795
rect 32413 10761 32447 10795
rect 3709 10693 3743 10727
rect 9965 10693 9999 10727
rect 10149 10693 10183 10727
rect 18705 10693 18739 10727
rect 22937 10693 22971 10727
rect 24409 10693 24443 10727
rect 28273 10693 28307 10727
rect 29101 10693 29135 10727
rect 29929 10693 29963 10727
rect 34529 10693 34563 10727
rect 1409 10625 1443 10659
rect 3249 10625 3283 10659
rect 3403 10625 3437 10659
rect 3985 10625 4019 10659
rect 4169 10625 4203 10659
rect 4813 10625 4847 10659
rect 5273 10625 5307 10659
rect 5457 10625 5491 10659
rect 5549 10625 5583 10659
rect 8125 10625 8159 10659
rect 8309 10625 8343 10659
rect 8401 10625 8435 10659
rect 8493 10625 8527 10659
rect 8861 10625 8895 10659
rect 8953 10625 8987 10659
rect 9229 10625 9263 10659
rect 9413 10625 9447 10659
rect 9505 10625 9539 10659
rect 9597 10625 9631 10659
rect 10333 10625 10367 10659
rect 10701 10625 10735 10659
rect 15209 10625 15243 10659
rect 15301 10625 15335 10659
rect 15485 10625 15519 10659
rect 17601 10625 17635 10659
rect 17877 10625 17911 10659
rect 18061 10625 18095 10659
rect 18337 10625 18371 10659
rect 19165 10625 19199 10659
rect 19625 10625 19659 10659
rect 20729 10625 20763 10659
rect 20913 10625 20947 10659
rect 21097 10625 21131 10659
rect 21189 10625 21223 10659
rect 21465 10625 21499 10659
rect 23121 10625 23155 10659
rect 27997 10625 28031 10659
rect 28733 10625 28767 10659
rect 29009 10625 29043 10659
rect 29285 10625 29319 10659
rect 30389 10625 30423 10659
rect 31677 10625 31711 10659
rect 31861 10625 31895 10659
rect 32321 10625 32355 10659
rect 32505 10625 32539 10659
rect 32689 10625 32723 10659
rect 32873 10625 32907 10659
rect 33057 10625 33091 10659
rect 1685 10557 1719 10591
rect 4721 10557 4755 10591
rect 8585 10557 8619 10591
rect 17693 10557 17727 10591
rect 18613 10557 18647 10591
rect 19073 10557 19107 10591
rect 19441 10557 19475 10591
rect 19901 10557 19935 10591
rect 21373 10557 21407 10591
rect 23305 10557 23339 10591
rect 25697 10557 25731 10591
rect 34253 10557 34287 10591
rect 5089 10489 5123 10523
rect 17785 10489 17819 10523
rect 18153 10489 18187 10523
rect 19349 10489 19383 10523
rect 20637 10489 20671 10523
rect 25421 10489 25455 10523
rect 28917 10489 28951 10523
rect 31861 10489 31895 10523
rect 3433 10421 3467 10455
rect 3893 10421 3927 10455
rect 4353 10421 4387 10455
rect 4445 10421 4479 10455
rect 9137 10421 9171 10455
rect 9873 10421 9907 10455
rect 15209 10421 15243 10455
rect 17417 10421 17451 10455
rect 18521 10421 18555 10455
rect 19073 10421 19107 10455
rect 19809 10421 19843 10455
rect 20361 10421 20395 10455
rect 20821 10421 20855 10455
rect 21189 10421 21223 10455
rect 24225 10421 24259 10455
rect 30021 10421 30055 10455
rect 33241 10421 33275 10455
rect 36001 10421 36035 10455
rect 1777 10217 1811 10251
rect 3801 10217 3835 10251
rect 4721 10217 4755 10251
rect 11713 10217 11747 10251
rect 12357 10217 12391 10251
rect 12541 10217 12575 10251
rect 14749 10217 14783 10251
rect 17417 10217 17451 10251
rect 20821 10217 20855 10251
rect 21005 10217 21039 10251
rect 23029 10217 23063 10251
rect 23213 10217 23247 10251
rect 24501 10217 24535 10251
rect 25053 10217 25087 10251
rect 25513 10217 25547 10251
rect 26893 10217 26927 10251
rect 31217 10217 31251 10251
rect 34437 10217 34471 10251
rect 6469 10149 6503 10183
rect 10793 10149 10827 10183
rect 17785 10149 17819 10183
rect 26709 10149 26743 10183
rect 28825 10149 28859 10183
rect 32597 10149 32631 10183
rect 33517 10149 33551 10183
rect 2053 10081 2087 10115
rect 2329 10081 2363 10115
rect 6193 10081 6227 10115
rect 9045 10081 9079 10115
rect 11253 10081 11287 10115
rect 12081 10081 12115 10115
rect 25605 10081 25639 10115
rect 27169 10081 27203 10115
rect 27445 10081 27479 10115
rect 29745 10081 29779 10115
rect 31401 10081 31435 10115
rect 34989 10081 35023 10115
rect 1685 10013 1719 10047
rect 1869 10013 1903 10047
rect 1961 10013 1995 10047
rect 2145 10013 2179 10047
rect 2421 10013 2455 10047
rect 3340 10013 3374 10047
rect 3433 10013 3467 10047
rect 3985 10013 4019 10047
rect 4077 10013 4111 10047
rect 4169 10013 4203 10047
rect 4287 10013 4321 10047
rect 4445 10013 4479 10047
rect 4721 10013 4755 10047
rect 5089 10013 5123 10047
rect 5457 10013 5491 10047
rect 5550 10013 5584 10047
rect 5825 10013 5859 10047
rect 5922 10013 5956 10047
rect 6745 10013 6779 10047
rect 6838 10013 6872 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 7941 10013 7975 10047
rect 8125 10013 8159 10047
rect 8218 10013 8252 10047
rect 8401 10013 8435 10047
rect 8629 10013 8663 10047
rect 10885 10013 10919 10047
rect 11069 10013 11103 10047
rect 11897 10013 11931 10047
rect 14933 10013 14967 10047
rect 15025 10013 15059 10047
rect 15209 10013 15243 10047
rect 15301 10013 15335 10047
rect 17601 10013 17635 10047
rect 17877 10013 17911 10047
rect 18153 10013 18187 10047
rect 21097 10013 21131 10047
rect 21189 10013 21223 10047
rect 24685 10013 24719 10047
rect 24869 10013 24903 10047
rect 25329 10013 25363 10047
rect 25421 10013 25455 10047
rect 25789 10013 25823 10047
rect 25881 10013 25915 10047
rect 26249 10013 26283 10047
rect 26985 10013 27019 10047
rect 27077 10013 27111 10047
rect 27537 10013 27571 10047
rect 27997 10013 28031 10047
rect 28089 10013 28123 10047
rect 28365 10013 28399 10047
rect 28457 10013 28491 10047
rect 28641 10013 28675 10047
rect 28917 10013 28951 10047
rect 29009 10013 29043 10047
rect 29561 10013 29595 10047
rect 30297 10013 30331 10047
rect 30573 10013 30607 10047
rect 31033 10013 31067 10047
rect 31217 10013 31251 10047
rect 31677 10013 31711 10047
rect 33701 10013 33735 10047
rect 33793 10013 33827 10047
rect 34713 10013 34747 10047
rect 3065 9945 3099 9979
rect 5733 9945 5767 9979
rect 8493 9945 8527 9979
rect 9321 9945 9355 9979
rect 12725 9945 12759 9979
rect 23397 9945 23431 9979
rect 27629 9945 27663 9979
rect 30113 9945 30147 9979
rect 32413 9945 32447 9979
rect 34069 9945 34103 9979
rect 34253 9945 34287 9979
rect 35633 9945 35667 9979
rect 36001 9945 36035 9979
rect 2789 9877 2823 9911
rect 4537 9877 4571 9911
rect 6101 9877 6135 9911
rect 6653 9877 6687 9911
rect 7113 9877 7147 9911
rect 7481 9877 7515 9911
rect 7849 9877 7883 9911
rect 8769 9877 8803 9911
rect 12525 9877 12559 9911
rect 18337 9877 18371 9911
rect 23213 9877 23247 9911
rect 27813 9877 27847 9911
rect 28549 9877 28583 9911
rect 29193 9877 29227 9911
rect 30205 9877 30239 9911
rect 30665 9877 30699 9911
rect 34161 9877 34195 9911
rect 3157 9673 3191 9707
rect 5457 9673 5491 9707
rect 8953 9673 8987 9707
rect 13277 9673 13311 9707
rect 22569 9673 22603 9707
rect 32229 9673 32263 9707
rect 35265 9673 35299 9707
rect 2329 9605 2363 9639
rect 2697 9605 2731 9639
rect 7021 9605 7055 9639
rect 11989 9605 12023 9639
rect 12617 9605 12651 9639
rect 12817 9605 12851 9639
rect 12909 9605 12943 9639
rect 16681 9605 16715 9639
rect 17049 9605 17083 9639
rect 19349 9605 19383 9639
rect 19533 9605 19567 9639
rect 22737 9605 22771 9639
rect 22937 9605 22971 9639
rect 26433 9605 26467 9639
rect 33333 9605 33367 9639
rect 33793 9605 33827 9639
rect 35725 9605 35759 9639
rect 2513 9537 2547 9571
rect 2973 9537 3007 9571
rect 3985 9537 4019 9571
rect 4169 9537 4203 9571
rect 4997 9537 5031 9571
rect 5181 9537 5215 9571
rect 5454 9537 5488 9571
rect 6009 9537 6043 9571
rect 6193 9537 6227 9571
rect 6377 9537 6411 9571
rect 6561 9537 6595 9571
rect 6924 9537 6958 9571
rect 7113 9537 7147 9571
rect 7296 9537 7330 9571
rect 7389 9537 7423 9571
rect 7665 9537 7699 9571
rect 7849 9537 7883 9571
rect 8217 9537 8251 9571
rect 8401 9537 8435 9571
rect 8677 9537 8711 9571
rect 8861 9537 8895 9571
rect 9137 9537 9171 9571
rect 9229 9537 9263 9571
rect 9413 9537 9447 9571
rect 9505 9537 9539 9571
rect 10425 9537 10459 9571
rect 10701 9537 10735 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 11069 9537 11103 9571
rect 11161 9537 11195 9571
rect 13093 9537 13127 9571
rect 13369 9537 13403 9571
rect 13829 9537 13863 9571
rect 14105 9537 14139 9571
rect 14749 9537 14783 9571
rect 14841 9537 14875 9571
rect 15209 9537 15243 9571
rect 16865 9537 16899 9571
rect 17141 9537 17175 9571
rect 19165 9537 19199 9571
rect 20821 9537 20855 9571
rect 20913 9537 20947 9571
rect 21005 9537 21039 9571
rect 21189 9537 21223 9571
rect 22089 9537 22123 9571
rect 22201 9537 22235 9571
rect 22293 9537 22327 9571
rect 22477 9537 22511 9571
rect 25605 9537 25639 9571
rect 26065 9537 26099 9571
rect 26341 9537 26375 9571
rect 26525 9537 26559 9571
rect 26709 9537 26743 9571
rect 26985 9537 27019 9571
rect 27169 9537 27203 9571
rect 27261 9537 27295 9571
rect 29837 9537 29871 9571
rect 30481 9537 30515 9571
rect 30665 9537 30699 9571
rect 31401 9537 31435 9571
rect 31585 9537 31619 9571
rect 32321 9537 32355 9571
rect 32413 9537 32447 9571
rect 33241 9537 33275 9571
rect 33425 9537 33459 9571
rect 33517 9537 33551 9571
rect 35541 9537 35575 9571
rect 2789 9469 2823 9503
rect 5089 9469 5123 9503
rect 5917 9469 5951 9503
rect 6101 9469 6135 9503
rect 8033 9469 8067 9503
rect 10333 9469 10367 9503
rect 11529 9469 11563 9503
rect 14013 9469 14047 9503
rect 15025 9469 15059 9503
rect 25789 9469 25823 9503
rect 29653 9469 29687 9503
rect 31769 9469 31803 9503
rect 8769 9401 8803 9435
rect 11713 9401 11747 9435
rect 13645 9401 13679 9435
rect 20637 9401 20671 9435
rect 25697 9401 25731 9435
rect 26157 9401 26191 9435
rect 26985 9401 27019 9435
rect 30021 9401 30055 9435
rect 30389 9401 30423 9435
rect 35909 9401 35943 9435
rect 4077 9333 4111 9367
rect 5273 9333 5307 9367
rect 5825 9333 5859 9367
rect 6561 9333 6595 9367
rect 6745 9333 6779 9367
rect 8585 9333 8619 9367
rect 10057 9333 10091 9367
rect 10425 9333 10459 9367
rect 10517 9333 10551 9367
rect 12449 9333 12483 9367
rect 12633 9333 12667 9367
rect 14105 9333 14139 9367
rect 14473 9333 14507 9367
rect 14933 9333 14967 9367
rect 21833 9333 21867 9367
rect 22753 9333 22787 9367
rect 25329 9333 25363 9367
rect 25881 9333 25915 9367
rect 35357 9333 35391 9367
rect 3617 9129 3651 9163
rect 7021 9129 7055 9163
rect 8677 9129 8711 9163
rect 11345 9129 11379 9163
rect 11713 9129 11747 9163
rect 16405 9129 16439 9163
rect 16865 9129 16899 9163
rect 18337 9129 18371 9163
rect 28457 9129 28491 9163
rect 30757 9129 30791 9163
rect 31401 9129 31435 9163
rect 32873 9129 32907 9163
rect 17601 9061 17635 9095
rect 23581 9061 23615 9095
rect 27353 9061 27387 9095
rect 30941 9061 30975 9095
rect 34069 9061 34103 9095
rect 34253 9061 34287 9095
rect 4997 8993 5031 9027
rect 9873 8993 9907 9027
rect 12817 8993 12851 9027
rect 16681 8993 16715 9027
rect 20085 8993 20119 9027
rect 20269 8993 20303 9027
rect 31769 8993 31803 9027
rect 33793 8993 33827 9027
rect 3341 8925 3375 8959
rect 3617 8925 3651 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 4537 8925 4571 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 5457 8925 5491 8959
rect 5733 8925 5767 8959
rect 6193 8925 6227 8959
rect 6377 8925 6411 8959
rect 6469 8925 6503 8959
rect 6653 8925 6687 8959
rect 6745 8925 6779 8959
rect 7112 8925 7146 8959
rect 7205 8925 7239 8959
rect 7481 8925 7515 8959
rect 7849 8925 7883 8959
rect 8769 8925 8803 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 9597 8925 9631 8959
rect 11529 8925 11563 8959
rect 11713 8925 11747 8959
rect 12725 8925 12759 8959
rect 16957 8925 16991 8959
rect 17049 8925 17083 8959
rect 17785 8925 17819 8959
rect 17877 8925 17911 8959
rect 18061 8925 18095 8959
rect 18153 8925 18187 8959
rect 18593 8925 18627 8959
rect 18705 8925 18739 8959
rect 18797 8925 18831 8959
rect 18981 8925 19015 8959
rect 20453 8925 20487 8959
rect 20637 8925 20671 8959
rect 23397 8925 23431 8959
rect 23489 8925 23523 8959
rect 23673 8925 23707 8959
rect 27169 8925 27203 8959
rect 27445 8925 27479 8959
rect 28457 8925 28491 8959
rect 28733 8925 28767 8959
rect 29193 8925 29227 8959
rect 29377 8925 29411 8959
rect 30113 8925 30147 8959
rect 31585 8925 31619 8959
rect 31861 8925 31895 8959
rect 32321 8925 32355 8959
rect 32505 8925 32539 8959
rect 32873 8925 32907 8959
rect 33057 8925 33091 8959
rect 34897 8925 34931 8959
rect 35265 8925 35299 8959
rect 3525 8857 3559 8891
rect 4353 8857 4387 8891
rect 7297 8857 7331 8891
rect 9229 8857 9263 8891
rect 17417 8857 17451 8891
rect 23213 8857 23247 8891
rect 26709 8857 26743 8891
rect 28641 8857 28675 8891
rect 30297 8857 30331 8891
rect 31217 8857 31251 8891
rect 3893 8789 3927 8823
rect 4261 8789 4295 8823
rect 4721 8789 4755 8823
rect 4905 8789 4939 8823
rect 5089 8789 5123 8823
rect 5273 8789 5307 8823
rect 5641 8789 5675 8823
rect 7665 8789 7699 8823
rect 9505 8789 9539 8823
rect 12265 8789 12299 8823
rect 12633 8789 12667 8823
rect 29101 8789 29135 8823
rect 30021 8789 30055 8823
rect 35081 8789 35115 8823
rect 35449 8789 35483 8823
rect 4261 8585 4295 8619
rect 6025 8585 6059 8619
rect 6377 8585 6411 8619
rect 9689 8585 9723 8619
rect 12725 8585 12759 8619
rect 16037 8585 16071 8619
rect 20269 8585 20303 8619
rect 23213 8585 23247 8619
rect 25329 8585 25363 8619
rect 4905 8517 4939 8551
rect 4997 8517 5031 8551
rect 5825 8517 5859 8551
rect 7757 8517 7791 8551
rect 8493 8517 8527 8551
rect 12541 8517 12575 8551
rect 16497 8517 16531 8551
rect 18337 8517 18371 8551
rect 30021 8517 30055 8551
rect 30849 8517 30883 8551
rect 31033 8517 31067 8551
rect 2513 8449 2547 8483
rect 4813 8449 4847 8483
rect 5181 8449 5215 8483
rect 5273 8449 5307 8483
rect 5365 8449 5399 8483
rect 5549 8449 5583 8483
rect 6653 8449 6687 8483
rect 6929 8449 6963 8483
rect 7113 8449 7147 8483
rect 7389 8449 7423 8483
rect 7573 8449 7607 8483
rect 7665 8449 7699 8483
rect 9229 8449 9263 8483
rect 9505 8449 9539 8483
rect 9689 8449 9723 8483
rect 10241 8449 10275 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 10793 8449 10827 8483
rect 11161 8449 11195 8483
rect 11345 8449 11379 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 11989 8449 12023 8483
rect 12081 8449 12115 8483
rect 12173 8449 12207 8483
rect 16221 8449 16255 8483
rect 16865 8449 16899 8483
rect 16957 8449 16991 8483
rect 17141 8449 17175 8483
rect 17233 8449 17267 8483
rect 18245 8449 18279 8483
rect 18613 8449 18647 8483
rect 20545 8449 20579 8483
rect 20637 8449 20671 8483
rect 23397 8449 23431 8483
rect 23673 8449 23707 8483
rect 25513 8449 25547 8483
rect 26157 8449 26191 8483
rect 29285 8449 29319 8483
rect 29837 8449 29871 8483
rect 30389 8449 30423 8483
rect 30665 8449 30699 8483
rect 31125 8449 31159 8483
rect 32873 8449 32907 8483
rect 33057 8449 33091 8483
rect 33517 8449 33551 8483
rect 34161 8449 34195 8483
rect 36093 8449 36127 8483
rect 2789 8381 2823 8415
rect 6377 8381 6411 8415
rect 8953 8381 8987 8415
rect 9045 8381 9079 8415
rect 9137 8381 9171 8415
rect 9781 8381 9815 8415
rect 11253 8381 11287 8415
rect 16313 8381 16347 8415
rect 18797 8381 18831 8415
rect 23581 8381 23615 8415
rect 25789 8381 25823 8415
rect 30481 8381 30515 8415
rect 33425 8381 33459 8415
rect 34345 8381 34379 8415
rect 35817 8381 35851 8415
rect 4629 8313 4663 8347
rect 6193 8313 6227 8347
rect 6561 8313 6595 8347
rect 6837 8313 6871 8347
rect 30849 8313 30883 8347
rect 32873 8313 32907 8347
rect 5733 8245 5767 8279
rect 6009 8245 6043 8279
rect 7205 8245 7239 8279
rect 8769 8245 8803 8279
rect 10793 8245 10827 8279
rect 11529 8245 11563 8279
rect 12541 8245 12575 8279
rect 16497 8245 16531 8279
rect 16681 8245 16715 8279
rect 20453 8245 20487 8279
rect 23673 8245 23707 8279
rect 25697 8245 25731 8279
rect 25973 8245 26007 8279
rect 30205 8245 30239 8279
rect 6377 8041 6411 8075
rect 7573 8041 7607 8075
rect 10057 8041 10091 8075
rect 15301 8041 15335 8075
rect 15853 8041 15887 8075
rect 23121 8041 23155 8075
rect 23305 8041 23339 8075
rect 25881 8041 25915 8075
rect 26985 8041 27019 8075
rect 29837 8041 29871 8075
rect 30113 8041 30147 8075
rect 35081 8041 35115 8075
rect 35357 8041 35391 8075
rect 5641 7973 5675 8007
rect 10425 7973 10459 8007
rect 13553 7973 13587 8007
rect 26801 7973 26835 8007
rect 30021 7973 30055 8007
rect 30481 7973 30515 8007
rect 35173 7973 35207 8007
rect 7389 7905 7423 7939
rect 9045 7905 9079 7939
rect 11161 7905 11195 7939
rect 11437 7905 11471 7939
rect 23213 7905 23247 7939
rect 24593 7905 24627 7939
rect 24777 7905 24811 7939
rect 26893 7905 26927 7939
rect 27813 7905 27847 7939
rect 28549 7905 28583 7939
rect 29929 7905 29963 7939
rect 35265 7905 35299 7939
rect 4353 7837 4387 7871
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 4813 7837 4847 7871
rect 5365 7837 5399 7871
rect 5733 7837 5767 7871
rect 6009 7837 6043 7871
rect 6561 7837 6595 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 7297 7837 7331 7871
rect 7665 7837 7699 7871
rect 10333 7837 10367 7871
rect 10517 7837 10551 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 13645 7837 13679 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 14565 7837 14599 7871
rect 14928 7837 14962 7871
rect 15117 7837 15151 7871
rect 15301 7837 15335 7871
rect 20821 7837 20855 7871
rect 21097 7837 21131 7871
rect 23029 7837 23063 7871
rect 23489 7837 23523 7871
rect 24501 7837 24535 7871
rect 24685 7837 24719 7871
rect 25329 7837 25363 7871
rect 25513 7837 25547 7871
rect 25697 7837 25731 7871
rect 25789 7837 25823 7871
rect 25881 7837 25915 7871
rect 26065 7837 26099 7871
rect 26341 7837 26375 7871
rect 26433 7837 26467 7871
rect 27445 7837 27479 7871
rect 27721 7837 27755 7871
rect 27905 7837 27939 7871
rect 28089 7837 28123 7871
rect 28641 7837 28675 7871
rect 28733 7837 28767 7871
rect 30573 7837 30607 7871
rect 30941 7837 30975 7871
rect 31125 7837 31159 7871
rect 34713 7837 34747 7871
rect 5641 7769 5675 7803
rect 5917 7769 5951 7803
rect 7021 7769 7055 7803
rect 8401 7769 8435 7803
rect 9229 7769 9263 7803
rect 9873 7769 9907 7803
rect 15025 7769 15059 7803
rect 15577 7769 15611 7803
rect 15761 7769 15795 7803
rect 25421 7769 25455 7803
rect 27353 7769 27387 7803
rect 4169 7701 4203 7735
rect 4721 7701 4755 7735
rect 5457 7701 5491 7735
rect 6009 7701 6043 7735
rect 6745 7701 6779 7735
rect 9321 7701 9355 7735
rect 9689 7701 9723 7735
rect 10073 7701 10107 7735
rect 10241 7701 10275 7735
rect 14749 7701 14783 7735
rect 20637 7701 20671 7735
rect 21005 7701 21039 7735
rect 22753 7701 22787 7735
rect 24961 7701 24995 7735
rect 25145 7701 25179 7735
rect 30665 7701 30699 7735
rect 2237 7497 2271 7531
rect 4445 7497 4479 7531
rect 5181 7497 5215 7531
rect 6009 7497 6043 7531
rect 8493 7497 8527 7531
rect 9137 7497 9171 7531
rect 10609 7497 10643 7531
rect 14105 7497 14139 7531
rect 15669 7497 15703 7531
rect 16681 7497 16715 7531
rect 18153 7497 18187 7531
rect 20269 7497 20303 7531
rect 27813 7497 27847 7531
rect 30849 7497 30883 7531
rect 31769 7497 31803 7531
rect 8769 7429 8803 7463
rect 8861 7429 8895 7463
rect 9505 7429 9539 7463
rect 11897 7429 11931 7463
rect 11989 7429 12023 7463
rect 14381 7429 14415 7463
rect 14749 7429 14783 7463
rect 19717 7429 19751 7463
rect 19917 7429 19951 7463
rect 21833 7429 21867 7463
rect 33057 7429 33091 7463
rect 3985 7361 4019 7395
rect 4537 7361 4571 7395
rect 5365 7361 5399 7395
rect 5457 7361 5491 7395
rect 5549 7361 5583 7395
rect 5733 7361 5767 7395
rect 5825 7361 5859 7395
rect 5917 7361 5951 7395
rect 6193 7361 6227 7395
rect 7205 7361 7239 7395
rect 7757 7361 7791 7395
rect 8677 7361 8711 7395
rect 9045 7361 9079 7395
rect 9321 7361 9355 7395
rect 9873 7361 9907 7395
rect 10149 7361 10183 7395
rect 10241 7361 10275 7395
rect 10425 7361 10459 7395
rect 10517 7361 10551 7395
rect 10885 7361 10919 7395
rect 11621 7361 11655 7395
rect 11713 7361 11747 7395
rect 12113 7361 12147 7395
rect 15485 7361 15519 7395
rect 15761 7361 15795 7395
rect 16865 7361 16899 7395
rect 17141 7361 17175 7395
rect 18613 7361 18647 7395
rect 18705 7361 18739 7395
rect 18889 7361 18923 7395
rect 20453 7361 20487 7395
rect 21649 7361 21683 7395
rect 22017 7361 22051 7395
rect 22293 7361 22327 7395
rect 22477 7361 22511 7395
rect 22845 7361 22879 7395
rect 22937 7361 22971 7395
rect 23029 7361 23063 7395
rect 23121 7361 23155 7395
rect 24961 7361 24995 7395
rect 25145 7361 25179 7395
rect 25513 7361 25547 7395
rect 25789 7361 25823 7395
rect 27721 7361 27755 7395
rect 27905 7361 27939 7395
rect 31033 7361 31067 7395
rect 31401 7361 31435 7395
rect 31677 7361 31711 7395
rect 31861 7361 31895 7395
rect 32321 7361 32355 7395
rect 32873 7361 32907 7395
rect 3709 7293 3743 7327
rect 4721 7293 4755 7327
rect 6377 7293 6411 7327
rect 6929 7293 6963 7327
rect 10793 7293 10827 7327
rect 10977 7293 11011 7327
rect 11069 7293 11103 7327
rect 12357 7293 12391 7327
rect 12633 7293 12667 7327
rect 17049 7293 17083 7327
rect 25697 7293 25731 7327
rect 31493 7293 31527 7327
rect 4077 7225 4111 7259
rect 6193 7225 6227 7259
rect 6653 7225 6687 7259
rect 7021 7225 7055 7259
rect 18429 7225 18463 7259
rect 18521 7225 18555 7259
rect 22109 7225 22143 7259
rect 22201 7225 22235 7259
rect 24961 7225 24995 7259
rect 25329 7225 25363 7259
rect 6837 7157 6871 7191
rect 7389 7157 7423 7191
rect 9781 7157 9815 7191
rect 9965 7157 9999 7191
rect 12265 7157 12299 7191
rect 15485 7157 15519 7191
rect 17141 7157 17175 7191
rect 19901 7157 19935 7191
rect 20085 7157 20119 7191
rect 21465 7157 21499 7191
rect 22661 7157 22695 7191
rect 25789 7157 25823 7191
rect 31033 7157 31067 7191
rect 4537 6953 4571 6987
rect 8585 6953 8619 6987
rect 9768 6953 9802 6987
rect 11621 6953 11655 6987
rect 13001 6953 13035 6987
rect 13369 6953 13403 6987
rect 14105 6953 14139 6987
rect 17785 6953 17819 6987
rect 17969 6953 18003 6987
rect 27077 6953 27111 6987
rect 27537 6953 27571 6987
rect 32597 6953 32631 6987
rect 18245 6885 18279 6919
rect 18797 6885 18831 6919
rect 19533 6885 19567 6919
rect 32781 6885 32815 6919
rect 4077 6817 4111 6851
rect 4261 6817 4295 6851
rect 4629 6817 4663 6851
rect 4905 6817 4939 6851
rect 4997 6817 5031 6851
rect 5641 6817 5675 6851
rect 5825 6817 5859 6851
rect 6837 6817 6871 6851
rect 6930 6817 6964 6851
rect 7021 6817 7055 6851
rect 9505 6817 9539 6851
rect 11529 6817 11563 6851
rect 14473 6817 14507 6851
rect 18613 6817 18647 6851
rect 18705 6817 18739 6851
rect 19625 6817 19659 6851
rect 29929 6817 29963 6851
rect 32689 6817 32723 6851
rect 4169 6749 4203 6783
rect 4353 6749 4387 6783
rect 4813 6749 4847 6783
rect 5089 6749 5123 6783
rect 5273 6749 5307 6783
rect 5365 6749 5399 6783
rect 5549 6749 5583 6783
rect 5733 6749 5767 6783
rect 6101 6749 6135 6783
rect 6377 6749 6411 6783
rect 7106 6749 7140 6783
rect 7665 6749 7699 6783
rect 7941 6749 7975 6783
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 8953 6749 8987 6783
rect 9229 6749 9263 6783
rect 11805 6749 11839 6783
rect 11989 6749 12023 6783
rect 12081 6749 12115 6783
rect 12909 6749 12943 6783
rect 13185 6749 13219 6783
rect 13369 6749 13403 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 18521 6749 18555 6783
rect 18981 6749 19015 6783
rect 19441 6749 19475 6783
rect 19717 6749 19751 6783
rect 19901 6749 19935 6783
rect 20269 6749 20303 6783
rect 29837 6749 29871 6783
rect 30021 6749 30055 6783
rect 33149 6749 33183 6783
rect 33241 6749 33275 6783
rect 5917 6681 5951 6715
rect 13553 6681 13587 6715
rect 18153 6681 18187 6715
rect 26893 6681 26927 6715
rect 27521 6681 27555 6715
rect 27721 6681 27755 6715
rect 6285 6613 6319 6647
rect 6653 6613 6687 6647
rect 7297 6613 7331 6647
rect 9045 6613 9079 6647
rect 9321 6613 9355 6647
rect 12265 6613 12299 6647
rect 17969 6613 18003 6647
rect 19257 6613 19291 6647
rect 27098 6613 27132 6647
rect 27261 6613 27295 6647
rect 27353 6613 27387 6647
rect 4353 6409 4387 6443
rect 5089 6409 5123 6443
rect 5365 6409 5399 6443
rect 6009 6409 6043 6443
rect 6469 6409 6503 6443
rect 8769 6409 8803 6443
rect 11345 6409 11379 6443
rect 12265 6409 12299 6443
rect 13553 6409 13587 6443
rect 13737 6409 13771 6443
rect 14105 6409 14139 6443
rect 18153 6409 18187 6443
rect 21373 6409 21407 6443
rect 23581 6409 23615 6443
rect 23949 6409 23983 6443
rect 24777 6409 24811 6443
rect 25881 6409 25915 6443
rect 26265 6409 26299 6443
rect 26433 6409 26467 6443
rect 29469 6409 29503 6443
rect 29929 6409 29963 6443
rect 33333 6409 33367 6443
rect 33609 6409 33643 6443
rect 5181 6341 5215 6375
rect 7297 6341 7331 6375
rect 9045 6341 9079 6375
rect 12909 6341 12943 6375
rect 15209 6341 15243 6375
rect 15425 6341 15459 6375
rect 17785 6341 17819 6375
rect 17985 6341 18019 6375
rect 21005 6341 21039 6375
rect 21221 6341 21255 6375
rect 24041 6341 24075 6375
rect 26065 6341 26099 6375
rect 29837 6341 29871 6375
rect 32229 6341 32263 6375
rect 32321 6341 32355 6375
rect 34069 6341 34103 6375
rect 4169 6273 4203 6307
rect 4261 6273 4295 6307
rect 4445 6273 4479 6307
rect 4721 6273 4755 6307
rect 5365 6273 5399 6307
rect 5457 6273 5491 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7021 6273 7055 6307
rect 9321 6273 9355 6307
rect 9597 6273 9631 6307
rect 11713 6273 11747 6307
rect 12173 6273 12207 6307
rect 12357 6273 12391 6307
rect 12817 6273 12851 6307
rect 13277 6273 13311 6307
rect 13829 6273 13863 6307
rect 14289 6273 14323 6307
rect 14381 6273 14415 6307
rect 14657 6273 14691 6307
rect 18613 6273 18647 6307
rect 18705 6273 18739 6307
rect 18797 6273 18831 6307
rect 18981 6273 19015 6307
rect 23857 6273 23891 6307
rect 24317 6273 24351 6307
rect 24691 6273 24725 6307
rect 24869 6273 24903 6307
rect 25329 6273 25363 6307
rect 25513 6273 25547 6307
rect 25789 6273 25823 6307
rect 27353 6273 27387 6307
rect 27721 6273 27755 6307
rect 28089 6273 28123 6307
rect 28457 6273 28491 6307
rect 29193 6273 29227 6307
rect 30021 6273 30055 6307
rect 30573 6273 30607 6307
rect 30849 6273 30883 6307
rect 31217 6273 31251 6307
rect 32689 6273 32723 6307
rect 32781 6273 32815 6307
rect 33241 6273 33275 6307
rect 33517 6273 33551 6307
rect 4813 6205 4847 6239
rect 5641 6205 5675 6239
rect 9137 6205 9171 6239
rect 9873 6205 9907 6239
rect 13093 6205 13127 6239
rect 13553 6205 13587 6239
rect 18337 6205 18371 6239
rect 27261 6205 27295 6239
rect 29285 6205 29319 6239
rect 30481 6205 30515 6239
rect 13369 6137 13403 6171
rect 24961 6137 24995 6171
rect 30205 6137 30239 6171
rect 34069 6137 34103 6171
rect 9045 6069 9079 6103
rect 9505 6069 9539 6103
rect 12449 6069 12483 6103
rect 14565 6069 14599 6103
rect 15393 6069 15427 6103
rect 15577 6069 15611 6103
rect 17969 6069 18003 6103
rect 21189 6069 21223 6103
rect 24225 6069 24259 6103
rect 26249 6069 26283 6103
rect 5273 5865 5307 5899
rect 7573 5865 7607 5899
rect 10885 5865 10919 5899
rect 12068 5865 12102 5899
rect 16221 5865 16255 5899
rect 17325 5865 17359 5899
rect 17509 5865 17543 5899
rect 20821 5865 20855 5899
rect 21005 5865 21039 5899
rect 22845 5865 22879 5899
rect 27905 5865 27939 5899
rect 31125 5865 31159 5899
rect 31953 5865 31987 5899
rect 10149 5797 10183 5831
rect 13829 5797 13863 5831
rect 21465 5797 21499 5831
rect 30665 5797 30699 5831
rect 31033 5797 31067 5831
rect 31493 5797 31527 5831
rect 9597 5729 9631 5763
rect 11529 5729 11563 5763
rect 11805 5729 11839 5763
rect 24501 5729 24535 5763
rect 24685 5729 24719 5763
rect 24869 5729 24903 5763
rect 26433 5729 26467 5763
rect 28457 5729 28491 5763
rect 29837 5729 29871 5763
rect 30941 5729 30975 5763
rect 32413 5729 32447 5763
rect 5181 5661 5215 5695
rect 5365 5661 5399 5695
rect 7573 5661 7607 5695
rect 7757 5661 7791 5695
rect 8585 5661 8619 5695
rect 9413 5661 9447 5695
rect 9505 5661 9539 5695
rect 10977 5661 11011 5695
rect 13737 5661 13771 5695
rect 14105 5661 14139 5695
rect 15025 5661 15059 5695
rect 15209 5661 15243 5695
rect 15301 5661 15335 5695
rect 15485 5661 15519 5695
rect 15577 5661 15611 5695
rect 16221 5661 16255 5695
rect 16497 5661 16531 5695
rect 19625 5661 19659 5695
rect 19717 5661 19751 5695
rect 19947 5661 19981 5695
rect 20085 5661 20119 5695
rect 21097 5661 21131 5695
rect 21373 5661 21407 5695
rect 21557 5661 21591 5695
rect 21649 5661 21683 5695
rect 21833 5661 21867 5695
rect 22845 5661 22879 5695
rect 23397 5661 23431 5695
rect 23765 5661 23799 5695
rect 24225 5661 24259 5695
rect 24777 5661 24811 5695
rect 24961 5661 24995 5695
rect 26893 5661 26927 5695
rect 26985 5661 27019 5695
rect 27077 5661 27111 5695
rect 27445 5661 27479 5695
rect 27813 5661 27847 5695
rect 27997 5661 28031 5695
rect 28825 5661 28859 5695
rect 29653 5661 29687 5695
rect 30205 5661 30239 5695
rect 30297 5661 30331 5695
rect 31585 5661 31619 5695
rect 31769 5661 31803 5695
rect 32229 5661 32263 5695
rect 32873 5661 32907 5695
rect 32965 5661 32999 5695
rect 10149 5593 10183 5627
rect 10609 5593 10643 5627
rect 17477 5593 17511 5627
rect 17693 5593 17727 5627
rect 19809 5593 19843 5627
rect 20637 5593 20671 5627
rect 20853 5593 20887 5627
rect 26525 5593 26559 5627
rect 28340 5593 28374 5627
rect 28549 5593 28583 5627
rect 30389 5593 30423 5627
rect 32781 5593 32815 5627
rect 8677 5525 8711 5559
rect 9045 5525 9079 5559
rect 10701 5525 10735 5559
rect 13553 5525 13587 5559
rect 14749 5525 14783 5559
rect 16405 5525 16439 5559
rect 19441 5525 19475 5559
rect 27629 5525 27663 5559
rect 28181 5525 28215 5559
rect 8125 5321 8159 5355
rect 19533 5321 19567 5355
rect 9597 5253 9631 5287
rect 10241 5253 10275 5287
rect 11069 5253 11103 5287
rect 14286 5253 14320 5287
rect 19685 5253 19719 5287
rect 19901 5253 19935 5287
rect 22109 5253 22143 5287
rect 9873 5185 9907 5219
rect 10977 5185 11011 5219
rect 11345 5185 11379 5219
rect 11529 5185 11563 5219
rect 15209 5185 15243 5219
rect 19073 5185 19107 5219
rect 19165 5185 19199 5219
rect 21925 5185 21959 5219
rect 22201 5185 22235 5219
rect 22293 5185 22327 5219
rect 22937 5185 22971 5219
rect 27169 5185 27203 5219
rect 27353 5185 27387 5219
rect 30205 5185 30239 5219
rect 30389 5185 30423 5219
rect 11069 5117 11103 5151
rect 11805 5117 11839 5151
rect 13461 5117 13495 5151
rect 15025 5117 15059 5151
rect 19441 5049 19475 5083
rect 22661 5049 22695 5083
rect 30389 5049 30423 5083
rect 11253 4981 11287 5015
rect 13277 4981 13311 5015
rect 14381 4981 14415 5015
rect 19257 4981 19291 5015
rect 19717 4981 19751 5015
rect 22477 4981 22511 5015
rect 26985 4981 27019 5015
rect 27353 4981 27387 5015
rect 11529 4777 11563 4811
rect 11713 4777 11747 4811
rect 16313 4777 16347 4811
rect 18521 4777 18555 4811
rect 21465 4777 21499 4811
rect 23949 4777 23983 4811
rect 14657 4709 14691 4743
rect 17509 4709 17543 4743
rect 17877 4709 17911 4743
rect 23213 4709 23247 4743
rect 8769 4641 8803 4675
rect 10977 4641 11011 4675
rect 11069 4641 11103 4675
rect 12449 4641 12483 4675
rect 13277 4641 13311 4675
rect 13369 4641 13403 4675
rect 15485 4641 15519 4675
rect 22661 4641 22695 4675
rect 8125 4573 8159 4607
rect 10701 4573 10735 4607
rect 11805 4573 11839 4607
rect 12265 4573 12299 4607
rect 13185 4573 13219 4607
rect 13645 4573 13679 4607
rect 14289 4573 14323 4607
rect 14381 4573 14415 4607
rect 14749 4573 14783 4607
rect 16037 4573 16071 4607
rect 16589 4573 16623 4607
rect 17601 4573 17635 4607
rect 17969 4573 18003 4607
rect 18153 4573 18187 4607
rect 18337 4573 18371 4607
rect 21649 4573 21683 4607
rect 21833 4573 21867 4607
rect 22293 4573 22327 4607
rect 23029 4573 23063 4607
rect 10425 4505 10459 4539
rect 14657 4505 14691 4539
rect 15393 4505 15427 4539
rect 17141 4505 17175 4539
rect 17325 4505 17359 4539
rect 17877 4505 17911 4539
rect 18245 4505 18279 4539
rect 23857 4505 23891 4539
rect 8953 4437 8987 4471
rect 11161 4437 11195 4471
rect 11897 4437 11931 4471
rect 12357 4437 12391 4471
rect 12817 4437 12851 4471
rect 13829 4437 13863 4471
rect 14197 4437 14231 4471
rect 14473 4437 14507 4471
rect 17693 4437 17727 4471
rect 21833 4437 21867 4471
rect 10701 4233 10735 4267
rect 15577 4233 15611 4267
rect 18429 4233 18463 4267
rect 21649 4233 21683 4267
rect 9873 4165 9907 4199
rect 24317 4165 24351 4199
rect 24409 4165 24443 4199
rect 9965 4097 9999 4131
rect 11529 4097 11563 4131
rect 11805 4097 11839 4131
rect 13829 4097 13863 4131
rect 15853 4097 15887 4131
rect 16129 4097 16163 4131
rect 16313 4097 16347 4131
rect 18061 4097 18095 4131
rect 18153 4097 18187 4131
rect 18337 4097 18371 4131
rect 18613 4097 18647 4131
rect 19257 4097 19291 4131
rect 21097 4097 21131 4131
rect 21281 4097 21315 4131
rect 21373 4097 21407 4131
rect 21465 4097 21499 4131
rect 24133 4097 24167 4131
rect 24501 4097 24535 4131
rect 25329 4097 25363 4131
rect 25697 4097 25731 4131
rect 28641 4097 28675 4131
rect 29009 4097 29043 4131
rect 8677 4029 8711 4063
rect 8861 4029 8895 4063
rect 10149 4029 10183 4063
rect 10793 4029 10827 4063
rect 10977 4029 11011 4063
rect 12081 4029 12115 4063
rect 14105 4029 14139 4063
rect 15945 4029 15979 4063
rect 16037 4029 16071 4063
rect 16681 4029 16715 4063
rect 17417 4029 17451 4063
rect 22201 4029 22235 4063
rect 22477 4029 22511 4063
rect 9413 3961 9447 3995
rect 19073 3961 19107 3995
rect 8033 3893 8067 3927
rect 9505 3893 9539 3927
rect 10333 3893 10367 3927
rect 11621 3893 11655 3927
rect 13553 3893 13587 3927
rect 15669 3893 15703 3927
rect 17325 3893 17359 3927
rect 18797 3893 18831 3927
rect 23949 3893 23983 3927
rect 24685 3893 24719 3927
rect 25697 3893 25731 3927
rect 25881 3893 25915 3927
rect 28457 3893 28491 3927
rect 28641 3893 28675 3927
rect 9413 3689 9447 3723
rect 13921 3689 13955 3723
rect 15301 3689 15335 3723
rect 19625 3689 19659 3723
rect 21557 3689 21591 3723
rect 24041 3689 24075 3723
rect 26617 3689 26651 3723
rect 27445 3689 27479 3723
rect 35909 3689 35943 3723
rect 7757 3621 7791 3655
rect 13185 3621 13219 3655
rect 14105 3621 14139 3655
rect 14933 3621 14967 3655
rect 20177 3621 20211 3655
rect 27169 3621 27203 3655
rect 8217 3553 8251 3587
rect 8309 3553 8343 3587
rect 10885 3553 10919 3587
rect 11161 3553 11195 3587
rect 11437 3553 11471 3587
rect 14565 3553 14599 3587
rect 14749 3553 14783 3587
rect 15577 3553 15611 3587
rect 17325 3553 17359 3587
rect 18245 3553 18279 3587
rect 21373 3553 21407 3587
rect 22293 3553 22327 3587
rect 22569 3553 22603 3587
rect 24409 3553 24443 3587
rect 25881 3553 25915 3587
rect 7941 3485 7975 3519
rect 8401 3485 8435 3519
rect 9321 3485 9355 3519
rect 13277 3485 13311 3519
rect 14473 3485 14507 3519
rect 15209 3485 15243 3519
rect 15485 3485 15519 3519
rect 17601 3485 17635 3519
rect 18981 3485 19015 3519
rect 19809 3485 19843 3519
rect 19901 3485 19935 3519
rect 20821 3485 20855 3519
rect 21097 3485 21131 3519
rect 21281 3485 21315 3519
rect 21833 3485 21867 3519
rect 21925 3485 21959 3519
rect 22017 3485 22051 3519
rect 22201 3485 22235 3519
rect 26157 3485 26191 3519
rect 26985 3485 27019 3519
rect 27537 3485 27571 3519
rect 27813 3485 27847 3519
rect 36093 3485 36127 3519
rect 11713 3417 11747 3451
rect 26801 3417 26835 3451
rect 8769 3349 8803 3383
rect 9137 3349 9171 3383
rect 17693 3349 17727 3383
rect 18429 3349 18463 3383
rect 26893 3349 26927 3383
rect 27261 3349 27295 3383
rect 12265 3145 12299 3179
rect 16129 3145 16163 3179
rect 16405 3145 16439 3179
rect 16957 3145 16991 3179
rect 9045 3077 9079 3111
rect 10977 3077 11011 3111
rect 12173 3077 12207 3111
rect 15577 3077 15611 3111
rect 19901 3077 19935 3111
rect 20453 3077 20487 3111
rect 20637 3077 20671 3111
rect 7849 3009 7883 3043
rect 8953 3009 8987 3043
rect 11253 3009 11287 3043
rect 14013 3009 14047 3043
rect 15853 3009 15887 3043
rect 15945 3009 15979 3043
rect 16221 3009 16255 3043
rect 16313 3009 16347 3043
rect 16497 3009 16531 3043
rect 16865 3009 16899 3043
rect 17141 3009 17175 3043
rect 17233 3009 17267 3043
rect 20361 3009 20395 3043
rect 21465 3009 21499 3043
rect 21649 3009 21683 3043
rect 21833 3009 21867 3043
rect 25421 3009 25455 3043
rect 8033 2941 8067 2975
rect 8861 2941 8895 2975
rect 11529 2941 11563 2975
rect 13737 2941 13771 2975
rect 14105 2941 14139 2975
rect 17509 2941 17543 2975
rect 19625 2941 19659 2975
rect 20177 2941 20211 2975
rect 22109 2941 22143 2975
rect 25145 2941 25179 2975
rect 9505 2873 9539 2907
rect 15945 2873 15979 2907
rect 17141 2873 17175 2907
rect 7665 2805 7699 2839
rect 8585 2805 8619 2839
rect 9413 2805 9447 2839
rect 18981 2805 19015 2839
rect 19073 2805 19107 2839
rect 20545 2805 20579 2839
rect 21281 2805 21315 2839
rect 23581 2805 23615 2839
rect 23673 2805 23707 2839
rect 7849 2601 7883 2635
rect 10701 2601 10735 2635
rect 13277 2601 13311 2635
rect 13461 2601 13495 2635
rect 18429 2601 18463 2635
rect 24869 2601 24903 2635
rect 16221 2533 16255 2567
rect 23949 2533 23983 2567
rect 24685 2533 24719 2567
rect 8953 2465 8987 2499
rect 11529 2465 11563 2499
rect 11805 2465 11839 2499
rect 14473 2465 14507 2499
rect 14749 2465 14783 2499
rect 16405 2465 16439 2499
rect 16681 2465 16715 2499
rect 16957 2465 16991 2499
rect 22753 2465 22787 2499
rect 23397 2465 23431 2499
rect 24409 2465 24443 2499
rect 8033 2397 8067 2431
rect 8401 2397 8435 2431
rect 8493 2397 8527 2431
rect 10793 2397 10827 2431
rect 11161 2397 11195 2431
rect 13553 2397 13587 2431
rect 13645 2397 13679 2431
rect 14105 2397 14139 2431
rect 16313 2397 16347 2431
rect 20729 2397 20763 2431
rect 21833 2397 21867 2431
rect 22201 2397 22235 2431
rect 22569 2397 22603 2431
rect 23029 2397 23063 2431
rect 23213 2397 23247 2431
rect 9229 2329 9263 2363
rect 8217 2261 8251 2295
rect 8677 2261 8711 2295
rect 13829 2261 13863 2295
rect 14289 2261 14323 2295
rect 20913 2261 20947 2295
<< metal1 >>
rect 1104 37562 36432 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 36432 37562
rect 1104 37488 36432 37510
rect 20809 37315 20867 37321
rect 16960 37284 17724 37312
rect 16960 37256 16988 37284
rect 16942 37204 16948 37256
rect 17000 37204 17006 37256
rect 17034 37204 17040 37256
rect 17092 37244 17098 37256
rect 17589 37247 17647 37253
rect 17589 37244 17601 37247
rect 17092 37216 17601 37244
rect 17092 37204 17098 37216
rect 17589 37213 17601 37216
rect 17635 37213 17647 37247
rect 17696 37244 17724 37284
rect 20809 37281 20821 37315
rect 20855 37312 20867 37315
rect 21082 37312 21088 37324
rect 20855 37284 21088 37312
rect 20855 37281 20867 37284
rect 20809 37275 20867 37281
rect 21082 37272 21088 37284
rect 21140 37272 21146 37324
rect 23569 37315 23627 37321
rect 23569 37281 23581 37315
rect 23615 37312 23627 37315
rect 25222 37312 25228 37324
rect 23615 37284 25228 37312
rect 23615 37281 23627 37284
rect 23569 37275 23627 37281
rect 25222 37272 25228 37284
rect 25280 37272 25286 37324
rect 22278 37244 22284 37256
rect 17696 37216 22284 37244
rect 17589 37207 17647 37213
rect 22278 37204 22284 37216
rect 22336 37204 22342 37256
rect 22462 37204 22468 37256
rect 22520 37204 22526 37256
rect 23842 37204 23848 37256
rect 23900 37204 23906 37256
rect 28994 37204 29000 37256
rect 29052 37244 29058 37256
rect 29089 37247 29147 37253
rect 29089 37244 29101 37247
rect 29052 37216 29101 37244
rect 29052 37204 29058 37216
rect 29089 37213 29101 37216
rect 29135 37213 29147 37247
rect 29089 37207 29147 37213
rect 29638 37204 29644 37256
rect 29696 37244 29702 37256
rect 29825 37247 29883 37253
rect 29825 37244 29837 37247
rect 29696 37216 29837 37244
rect 29696 37204 29702 37216
rect 29825 37213 29837 37216
rect 29871 37213 29883 37247
rect 29825 37207 29883 37213
rect 16574 37136 16580 37188
rect 16632 37176 16638 37188
rect 17310 37176 17316 37188
rect 16632 37148 17316 37176
rect 16632 37136 16638 37148
rect 17310 37136 17316 37148
rect 17368 37176 17374 37188
rect 17405 37179 17463 37185
rect 17405 37176 17417 37179
rect 17368 37148 17417 37176
rect 17368 37136 17374 37148
rect 17405 37145 17417 37148
rect 17451 37145 17463 37179
rect 17405 37139 17463 37145
rect 18874 37136 18880 37188
rect 18932 37176 18938 37188
rect 20533 37179 20591 37185
rect 20533 37176 20545 37179
rect 18932 37148 20545 37176
rect 18932 37136 18938 37148
rect 20533 37145 20545 37148
rect 20579 37145 20591 37179
rect 20533 37139 20591 37145
rect 21821 37179 21879 37185
rect 21821 37145 21833 37179
rect 21867 37176 21879 37179
rect 22186 37176 22192 37188
rect 21867 37148 22192 37176
rect 21867 37145 21879 37148
rect 21821 37139 21879 37145
rect 22186 37136 22192 37148
rect 22244 37136 22250 37188
rect 17494 37068 17500 37120
rect 17552 37108 17558 37120
rect 17773 37111 17831 37117
rect 17773 37108 17785 37111
rect 17552 37080 17785 37108
rect 17552 37068 17558 37080
rect 17773 37077 17785 37080
rect 17819 37108 17831 37111
rect 18782 37108 18788 37120
rect 17819 37080 18788 37108
rect 17819 37077 17831 37080
rect 17773 37071 17831 37077
rect 18782 37068 18788 37080
rect 18840 37068 18846 37120
rect 20162 37068 20168 37120
rect 20220 37068 20226 37120
rect 20625 37111 20683 37117
rect 20625 37077 20637 37111
rect 20671 37108 20683 37111
rect 21910 37108 21916 37120
rect 20671 37080 21916 37108
rect 20671 37077 20683 37080
rect 20625 37071 20683 37077
rect 21910 37068 21916 37080
rect 21968 37108 21974 37120
rect 23750 37108 23756 37120
rect 21968 37080 23756 37108
rect 21968 37068 21974 37080
rect 23750 37068 23756 37080
rect 23808 37068 23814 37120
rect 29270 37068 29276 37120
rect 29328 37068 29334 37120
rect 29730 37068 29736 37120
rect 29788 37108 29794 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29788 37080 29929 37108
rect 29788 37068 29794 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 1104 37018 36432 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 36432 37018
rect 1104 36944 36432 36966
rect 15473 36907 15531 36913
rect 9784 36876 14044 36904
rect 9674 36796 9680 36848
rect 9732 36836 9738 36848
rect 9784 36836 9812 36876
rect 9732 36808 9890 36836
rect 9732 36796 9738 36808
rect 14016 36768 14044 36876
rect 15473 36873 15485 36907
rect 15519 36904 15531 36907
rect 16114 36904 16120 36916
rect 15519 36876 16120 36904
rect 15519 36873 15531 36876
rect 15473 36867 15531 36873
rect 16114 36864 16120 36876
rect 16172 36904 16178 36916
rect 22554 36904 22560 36916
rect 16172 36876 16712 36904
rect 16172 36864 16178 36876
rect 15105 36839 15163 36845
rect 15105 36805 15117 36839
rect 15151 36836 15163 36839
rect 16574 36836 16580 36848
rect 15151 36808 16068 36836
rect 15151 36805 15163 36808
rect 15105 36799 15163 36805
rect 14826 36768 14832 36780
rect 14016 36754 14832 36768
rect 14030 36740 14832 36754
rect 14826 36728 14832 36740
rect 14884 36728 14890 36780
rect 14918 36728 14924 36780
rect 14976 36728 14982 36780
rect 15197 36771 15255 36777
rect 15197 36737 15209 36771
rect 15243 36768 15255 36771
rect 15286 36768 15292 36780
rect 15243 36740 15292 36768
rect 15243 36737 15255 36740
rect 15197 36731 15255 36737
rect 15286 36728 15292 36740
rect 15344 36728 15350 36780
rect 15565 36771 15623 36777
rect 15565 36768 15577 36771
rect 15396 36740 15577 36768
rect 9309 36703 9367 36709
rect 9309 36669 9321 36703
rect 9355 36700 9367 36703
rect 10686 36700 10692 36712
rect 9355 36672 10692 36700
rect 9355 36669 9367 36672
rect 9309 36663 9367 36669
rect 10686 36660 10692 36672
rect 10744 36660 10750 36712
rect 11054 36660 11060 36712
rect 11112 36660 11118 36712
rect 11333 36703 11391 36709
rect 11333 36669 11345 36703
rect 11379 36700 11391 36703
rect 12618 36700 12624 36712
rect 11379 36672 12624 36700
rect 11379 36669 11391 36672
rect 11333 36663 11391 36669
rect 12618 36660 12624 36672
rect 12676 36660 12682 36712
rect 12897 36703 12955 36709
rect 12897 36669 12909 36703
rect 12943 36700 12955 36703
rect 13262 36700 13268 36712
rect 12943 36672 13268 36700
rect 12943 36669 12955 36672
rect 12897 36663 12955 36669
rect 13262 36660 13268 36672
rect 13320 36660 13326 36712
rect 14090 36660 14096 36712
rect 14148 36700 14154 36712
rect 14645 36703 14703 36709
rect 14645 36700 14657 36703
rect 14148 36672 14657 36700
rect 14148 36660 14154 36672
rect 14645 36669 14657 36672
rect 14691 36669 14703 36703
rect 14645 36663 14703 36669
rect 14734 36660 14740 36712
rect 14792 36700 14798 36712
rect 15396 36700 15424 36740
rect 15565 36737 15577 36740
rect 15611 36737 15623 36771
rect 15565 36731 15623 36737
rect 15749 36771 15807 36777
rect 15749 36737 15761 36771
rect 15795 36737 15807 36771
rect 15749 36731 15807 36737
rect 14792 36672 15424 36700
rect 15473 36703 15531 36709
rect 14792 36660 14798 36672
rect 15473 36669 15485 36703
rect 15519 36700 15531 36703
rect 15657 36703 15715 36709
rect 15657 36700 15669 36703
rect 15519 36672 15669 36700
rect 15519 36669 15531 36672
rect 15473 36663 15531 36669
rect 15657 36669 15669 36672
rect 15703 36669 15715 36703
rect 15764 36700 15792 36731
rect 15838 36728 15844 36780
rect 15896 36728 15902 36780
rect 16040 36777 16068 36808
rect 16316 36808 16580 36836
rect 16316 36777 16344 36808
rect 16574 36796 16580 36808
rect 16632 36796 16638 36848
rect 16025 36771 16083 36777
rect 16025 36737 16037 36771
rect 16071 36737 16083 36771
rect 16025 36731 16083 36737
rect 16301 36771 16359 36777
rect 16301 36737 16313 36771
rect 16347 36737 16359 36771
rect 16301 36731 16359 36737
rect 16316 36700 16344 36731
rect 16482 36728 16488 36780
rect 16540 36728 16546 36780
rect 16684 36777 16712 36876
rect 17328 36876 19104 36904
rect 17328 36777 17356 36876
rect 17405 36839 17463 36845
rect 17405 36805 17417 36839
rect 17451 36836 17463 36839
rect 17770 36836 17776 36848
rect 17451 36808 17776 36836
rect 17451 36805 17463 36808
rect 17405 36799 17463 36805
rect 17770 36796 17776 36808
rect 17828 36796 17834 36848
rect 18037 36781 18095 36787
rect 16669 36771 16727 36777
rect 16669 36737 16681 36771
rect 16715 36737 16727 36771
rect 16669 36731 16727 36737
rect 16823 36771 16881 36777
rect 16823 36737 16835 36771
rect 16869 36768 16881 36771
rect 17037 36771 17095 36777
rect 16869 36737 16896 36768
rect 16823 36731 16896 36737
rect 17037 36737 17049 36771
rect 17083 36768 17095 36771
rect 17313 36771 17371 36777
rect 17313 36768 17325 36771
rect 17083 36740 17325 36768
rect 17083 36737 17095 36740
rect 17037 36731 17095 36737
rect 17313 36737 17325 36740
rect 17359 36737 17371 36771
rect 17313 36731 17371 36737
rect 15764 36672 16344 36700
rect 16393 36703 16451 36709
rect 15657 36663 15715 36669
rect 16393 36669 16405 36703
rect 16439 36700 16451 36703
rect 16868 36700 16896 36731
rect 17494 36728 17500 36780
rect 17552 36728 17558 36780
rect 17586 36728 17592 36780
rect 17644 36777 17650 36780
rect 18037 36778 18049 36781
rect 17644 36771 17673 36777
rect 17661 36737 17673 36771
rect 17644 36731 17673 36737
rect 17972 36750 18049 36778
rect 17644 36728 17650 36731
rect 17218 36700 17224 36712
rect 16439 36672 17224 36700
rect 16439 36669 16451 36672
rect 16393 36663 16451 36669
rect 17218 36660 17224 36672
rect 17276 36660 17282 36712
rect 17773 36703 17831 36709
rect 17773 36669 17785 36703
rect 17819 36700 17831 36703
rect 17862 36700 17868 36712
rect 17819 36672 17868 36700
rect 17819 36669 17831 36672
rect 17773 36663 17831 36669
rect 17862 36660 17868 36672
rect 17920 36660 17926 36712
rect 14274 36592 14280 36644
rect 14332 36632 14338 36644
rect 15841 36635 15899 36641
rect 15841 36632 15853 36635
rect 14332 36604 15853 36632
rect 14332 36592 14338 36604
rect 15841 36601 15853 36604
rect 15887 36601 15899 36635
rect 15841 36595 15899 36601
rect 17972 36576 18000 36750
rect 18037 36747 18049 36750
rect 18083 36747 18095 36781
rect 18037 36741 18095 36747
rect 18230 36728 18236 36780
rect 18288 36728 18294 36780
rect 18601 36771 18659 36777
rect 18601 36768 18613 36771
rect 18524 36740 18613 36768
rect 18138 36660 18144 36712
rect 18196 36660 18202 36712
rect 18322 36660 18328 36712
rect 18380 36660 18386 36712
rect 18414 36660 18420 36712
rect 18472 36660 18478 36712
rect 18156 36632 18184 36660
rect 18524 36632 18552 36740
rect 18601 36737 18613 36740
rect 18647 36737 18659 36771
rect 18601 36731 18659 36737
rect 18782 36728 18788 36780
rect 18840 36768 18846 36780
rect 19076 36777 19104 36876
rect 21836 36876 22560 36904
rect 21836 36845 21864 36876
rect 22554 36864 22560 36876
rect 22612 36864 22618 36916
rect 21821 36839 21879 36845
rect 21821 36805 21833 36839
rect 21867 36805 21879 36839
rect 21821 36799 21879 36805
rect 23290 36796 23296 36848
rect 23348 36836 23354 36848
rect 25774 36836 25780 36848
rect 23348 36808 25780 36836
rect 23348 36796 23354 36808
rect 25774 36796 25780 36808
rect 25832 36796 25838 36848
rect 18877 36771 18935 36777
rect 18877 36768 18889 36771
rect 18840 36740 18889 36768
rect 18840 36728 18846 36740
rect 18877 36737 18889 36740
rect 18923 36737 18935 36771
rect 18877 36731 18935 36737
rect 19061 36771 19119 36777
rect 19061 36737 19073 36771
rect 19107 36737 19119 36771
rect 22094 36768 22100 36780
rect 20746 36740 22100 36768
rect 19061 36731 19119 36737
rect 22094 36728 22100 36740
rect 22152 36768 22158 36780
rect 22462 36768 22468 36780
rect 22152 36740 22468 36768
rect 22152 36728 22158 36740
rect 22462 36728 22468 36740
rect 22520 36728 22526 36780
rect 23842 36728 23848 36780
rect 23900 36728 23906 36780
rect 18690 36660 18696 36712
rect 18748 36700 18754 36712
rect 19337 36703 19395 36709
rect 19337 36700 19349 36703
rect 18748 36672 19349 36700
rect 18748 36660 18754 36672
rect 19337 36669 19349 36672
rect 19383 36669 19395 36703
rect 19337 36663 19395 36669
rect 19610 36660 19616 36712
rect 19668 36660 19674 36712
rect 21361 36703 21419 36709
rect 21361 36669 21373 36703
rect 21407 36669 21419 36703
rect 23474 36700 23480 36712
rect 21361 36663 21419 36669
rect 22066 36672 23480 36700
rect 18156 36604 18552 36632
rect 18598 36592 18604 36644
rect 18656 36632 18662 36644
rect 18969 36635 19027 36641
rect 18969 36632 18981 36635
rect 18656 36604 18981 36632
rect 18656 36592 18662 36604
rect 18969 36601 18981 36604
rect 19015 36601 19027 36635
rect 21376 36632 21404 36663
rect 22066 36632 22094 36672
rect 23474 36660 23480 36672
rect 23532 36660 23538 36712
rect 23569 36703 23627 36709
rect 23569 36669 23581 36703
rect 23615 36700 23627 36703
rect 24394 36700 24400 36712
rect 23615 36672 24400 36700
rect 23615 36669 23627 36672
rect 23569 36663 23627 36669
rect 24394 36660 24400 36672
rect 24452 36660 24458 36712
rect 21376 36604 22094 36632
rect 18969 36595 19027 36601
rect 12710 36524 12716 36576
rect 12768 36564 12774 36576
rect 13630 36564 13636 36576
rect 12768 36536 13636 36564
rect 12768 36524 12774 36536
rect 13630 36524 13636 36536
rect 13688 36524 13694 36576
rect 14182 36524 14188 36576
rect 14240 36564 14246 36576
rect 15289 36567 15347 36573
rect 15289 36564 15301 36567
rect 14240 36536 15301 36564
rect 14240 36524 14246 36536
rect 15289 36533 15301 36536
rect 15335 36533 15347 36567
rect 15289 36527 15347 36533
rect 17126 36524 17132 36576
rect 17184 36524 17190 36576
rect 17954 36524 17960 36576
rect 18012 36524 18018 36576
rect 18138 36524 18144 36576
rect 18196 36564 18202 36576
rect 18322 36564 18328 36576
rect 18196 36536 18328 36564
rect 18196 36524 18202 36536
rect 18322 36524 18328 36536
rect 18380 36524 18386 36576
rect 18782 36524 18788 36576
rect 18840 36524 18846 36576
rect 22186 36524 22192 36576
rect 22244 36564 22250 36576
rect 23198 36564 23204 36576
rect 22244 36536 23204 36564
rect 22244 36524 22250 36536
rect 23198 36524 23204 36536
rect 23256 36564 23262 36576
rect 23382 36564 23388 36576
rect 23256 36536 23388 36564
rect 23256 36524 23262 36536
rect 23382 36524 23388 36536
rect 23440 36524 23446 36576
rect 1104 36474 36432 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 36432 36474
rect 1104 36400 36432 36422
rect 13262 36320 13268 36372
rect 13320 36320 13326 36372
rect 13630 36320 13636 36372
rect 13688 36360 13694 36372
rect 16666 36360 16672 36372
rect 13688 36332 16672 36360
rect 13688 36320 13694 36332
rect 16666 36320 16672 36332
rect 16724 36360 16730 36372
rect 16945 36363 17003 36369
rect 16945 36360 16957 36363
rect 16724 36332 16957 36360
rect 16724 36320 16730 36332
rect 16945 36329 16957 36332
rect 16991 36360 17003 36363
rect 17034 36360 17040 36372
rect 16991 36332 17040 36360
rect 16991 36329 17003 36332
rect 16945 36323 17003 36329
rect 17034 36320 17040 36332
rect 17092 36320 17098 36372
rect 17954 36320 17960 36372
rect 18012 36360 18018 36372
rect 19245 36363 19303 36369
rect 19245 36360 19257 36363
rect 18012 36332 19257 36360
rect 18012 36320 18018 36332
rect 19245 36329 19257 36332
rect 19291 36329 19303 36363
rect 19245 36323 19303 36329
rect 19610 36320 19616 36372
rect 19668 36360 19674 36372
rect 22833 36363 22891 36369
rect 22833 36360 22845 36363
rect 19668 36332 22845 36360
rect 19668 36320 19674 36332
rect 22833 36329 22845 36332
rect 22879 36329 22891 36363
rect 22833 36323 22891 36329
rect 24394 36320 24400 36372
rect 24452 36320 24458 36372
rect 25222 36320 25228 36372
rect 25280 36320 25286 36372
rect 8938 36252 8944 36304
rect 8996 36292 9002 36304
rect 9401 36295 9459 36301
rect 9401 36292 9413 36295
rect 8996 36264 9413 36292
rect 8996 36252 9002 36264
rect 9401 36261 9413 36264
rect 9447 36261 9459 36295
rect 9401 36255 9459 36261
rect 12618 36252 12624 36304
rect 12676 36292 12682 36304
rect 12676 36264 15516 36292
rect 12676 36252 12682 36264
rect 8294 36184 8300 36236
rect 8352 36224 8358 36236
rect 10137 36227 10195 36233
rect 10137 36224 10149 36227
rect 8352 36196 10149 36224
rect 8352 36184 8358 36196
rect 10137 36193 10149 36196
rect 10183 36193 10195 36227
rect 10137 36187 10195 36193
rect 13354 36184 13360 36236
rect 13412 36184 13418 36236
rect 13538 36184 13544 36236
rect 13596 36224 13602 36236
rect 13633 36227 13691 36233
rect 13633 36224 13645 36227
rect 13596 36196 13645 36224
rect 13596 36184 13602 36196
rect 13633 36193 13645 36196
rect 13679 36193 13691 36227
rect 13633 36187 13691 36193
rect 14182 36184 14188 36236
rect 14240 36184 14246 36236
rect 15488 36224 15516 36264
rect 18708 36264 19932 36292
rect 18708 36236 18736 36264
rect 16761 36227 16819 36233
rect 16761 36224 16773 36227
rect 15488 36196 16773 36224
rect 16761 36193 16773 36196
rect 16807 36224 16819 36227
rect 18414 36224 18420 36236
rect 16807 36196 18420 36224
rect 16807 36193 16819 36196
rect 16761 36187 16819 36193
rect 18414 36184 18420 36196
rect 18472 36224 18478 36236
rect 18690 36224 18696 36236
rect 18472 36196 18696 36224
rect 18472 36184 18478 36196
rect 18690 36184 18696 36196
rect 18748 36184 18754 36236
rect 18785 36227 18843 36233
rect 18785 36193 18797 36227
rect 18831 36193 18843 36227
rect 18785 36187 18843 36193
rect 18969 36227 19027 36233
rect 18969 36193 18981 36227
rect 19015 36224 19027 36227
rect 19015 36196 19196 36224
rect 19015 36193 19027 36196
rect 18969 36187 19027 36193
rect 5994 36116 6000 36168
rect 6052 36156 6058 36168
rect 7193 36159 7251 36165
rect 7193 36156 7205 36159
rect 6052 36128 7205 36156
rect 6052 36116 6058 36128
rect 7193 36125 7205 36128
rect 7239 36125 7251 36159
rect 7193 36119 7251 36125
rect 7377 36159 7435 36165
rect 7377 36125 7389 36159
rect 7423 36156 7435 36159
rect 7834 36156 7840 36168
rect 7423 36128 7840 36156
rect 7423 36125 7435 36128
rect 7377 36119 7435 36125
rect 7834 36116 7840 36128
rect 7892 36116 7898 36168
rect 9306 36116 9312 36168
rect 9364 36116 9370 36168
rect 9677 36159 9735 36165
rect 9677 36125 9689 36159
rect 9723 36125 9735 36159
rect 9677 36119 9735 36125
rect 9582 36048 9588 36100
rect 9640 36048 9646 36100
rect 7098 35980 7104 36032
rect 7156 36020 7162 36032
rect 7285 36023 7343 36029
rect 7285 36020 7297 36023
rect 7156 35992 7297 36020
rect 7156 35980 7162 35992
rect 7285 35989 7297 35992
rect 7331 35989 7343 36023
rect 7285 35983 7343 35989
rect 9309 36023 9367 36029
rect 9309 35989 9321 36023
rect 9355 36020 9367 36023
rect 9692 36020 9720 36119
rect 9766 36116 9772 36168
rect 9824 36116 9830 36168
rect 9858 36116 9864 36168
rect 9916 36116 9922 36168
rect 12618 36116 12624 36168
rect 12676 36116 12682 36168
rect 12802 36116 12808 36168
rect 12860 36116 12866 36168
rect 12894 36116 12900 36168
rect 12952 36116 12958 36168
rect 12986 36116 12992 36168
rect 13044 36116 13050 36168
rect 13170 36116 13176 36168
rect 13228 36156 13234 36168
rect 13725 36159 13783 36165
rect 13725 36156 13737 36159
rect 13228 36128 13737 36156
rect 13228 36116 13234 36128
rect 13725 36125 13737 36128
rect 13771 36156 13783 36159
rect 14090 36156 14096 36168
rect 13771 36128 14096 36156
rect 13771 36125 13783 36128
rect 13725 36119 13783 36125
rect 14090 36116 14096 36128
rect 14148 36116 14154 36168
rect 14274 36116 14280 36168
rect 14332 36116 14338 36168
rect 14826 36116 14832 36168
rect 14884 36156 14890 36168
rect 14884 36142 15410 36156
rect 14884 36128 15424 36142
rect 14884 36116 14890 36128
rect 9784 36088 9812 36116
rect 9784 36060 10364 36088
rect 9355 35992 9720 36020
rect 9769 36023 9827 36029
rect 9355 35989 9367 35992
rect 9309 35983 9367 35989
rect 9769 35989 9781 36023
rect 9815 36020 9827 36023
rect 10134 36020 10140 36032
rect 9815 35992 10140 36020
rect 9815 35989 9827 35992
rect 9769 35983 9827 35989
rect 10134 35980 10140 35992
rect 10192 35980 10198 36032
rect 10336 36020 10364 36060
rect 10410 36048 10416 36100
rect 10468 36048 10474 36100
rect 10520 36060 10902 36088
rect 10520 36020 10548 36060
rect 12158 36048 12164 36100
rect 12216 36048 12222 36100
rect 14734 36048 14740 36100
rect 14792 36048 14798 36100
rect 10336 35992 10548 36020
rect 14645 36023 14703 36029
rect 14645 35989 14657 36023
rect 14691 36020 14703 36023
rect 15194 36020 15200 36032
rect 14691 35992 15200 36020
rect 14691 35989 14703 35992
rect 14645 35983 14703 35989
rect 15194 35980 15200 35992
rect 15252 35980 15258 36032
rect 15396 36020 15424 36128
rect 16482 36048 16488 36100
rect 16540 36048 16546 36100
rect 16592 36060 17250 36088
rect 16592 36020 16620 36060
rect 18322 36048 18328 36100
rect 18380 36088 18386 36100
rect 18417 36091 18475 36097
rect 18417 36088 18429 36091
rect 18380 36060 18429 36088
rect 18380 36048 18386 36060
rect 18417 36057 18429 36060
rect 18463 36057 18475 36091
rect 18417 36051 18475 36057
rect 18506 36048 18512 36100
rect 18564 36088 18570 36100
rect 18800 36088 18828 36187
rect 19058 36116 19064 36168
rect 19116 36116 19122 36168
rect 19168 36156 19196 36196
rect 19242 36184 19248 36236
rect 19300 36224 19306 36236
rect 19794 36224 19800 36236
rect 19300 36196 19800 36224
rect 19300 36184 19306 36196
rect 19794 36184 19800 36196
rect 19852 36184 19858 36236
rect 19904 36233 19932 36264
rect 21192 36264 22692 36292
rect 19889 36227 19947 36233
rect 19889 36193 19901 36227
rect 19935 36193 19947 36227
rect 19889 36187 19947 36193
rect 20162 36184 20168 36236
rect 20220 36184 20226 36236
rect 20254 36184 20260 36236
rect 20312 36224 20318 36236
rect 21192 36224 21220 36264
rect 20312 36196 21220 36224
rect 20312 36184 20318 36196
rect 21910 36184 21916 36236
rect 21968 36184 21974 36236
rect 22186 36184 22192 36236
rect 22244 36224 22250 36236
rect 22557 36227 22615 36233
rect 22557 36224 22569 36227
rect 22244 36196 22569 36224
rect 22244 36184 22250 36196
rect 22557 36193 22569 36196
rect 22603 36193 22615 36227
rect 22557 36187 22615 36193
rect 19334 36156 19340 36168
rect 19168 36128 19340 36156
rect 19334 36116 19340 36128
rect 19392 36116 19398 36168
rect 19429 36159 19487 36165
rect 19429 36125 19441 36159
rect 19475 36125 19487 36159
rect 19429 36119 19487 36125
rect 18564 36060 18828 36088
rect 18564 36048 18570 36060
rect 19150 36048 19156 36100
rect 19208 36088 19214 36100
rect 19444 36088 19472 36119
rect 19518 36116 19524 36168
rect 19576 36156 19582 36168
rect 19705 36159 19763 36165
rect 19705 36156 19717 36159
rect 19576 36128 19717 36156
rect 19576 36116 19582 36128
rect 19705 36125 19717 36128
rect 19751 36125 19763 36159
rect 21298 36128 22048 36156
rect 19705 36119 19763 36125
rect 19208 36060 19472 36088
rect 19720 36088 19748 36119
rect 20254 36088 20260 36100
rect 19720 36060 20260 36088
rect 19208 36048 19214 36060
rect 20254 36048 20260 36060
rect 20312 36048 20318 36100
rect 22020 36088 22048 36128
rect 22278 36116 22284 36168
rect 22336 36156 22342 36168
rect 22373 36159 22431 36165
rect 22373 36156 22385 36159
rect 22336 36128 22385 36156
rect 22336 36116 22342 36128
rect 22373 36125 22385 36128
rect 22419 36125 22431 36159
rect 22664 36156 22692 36264
rect 22738 36184 22744 36236
rect 22796 36224 22802 36236
rect 22796 36196 23336 36224
rect 22796 36184 22802 36196
rect 23201 36159 23259 36165
rect 23201 36156 23213 36159
rect 22664 36128 23213 36156
rect 22373 36119 22431 36125
rect 23201 36125 23213 36128
rect 23247 36125 23259 36159
rect 23308 36156 23336 36196
rect 23474 36184 23480 36236
rect 23532 36224 23538 36236
rect 25038 36224 25044 36236
rect 23532 36196 25044 36224
rect 23532 36184 23538 36196
rect 25038 36184 25044 36196
rect 25096 36224 25102 36236
rect 25777 36227 25835 36233
rect 25777 36224 25789 36227
rect 25096 36196 25789 36224
rect 25096 36184 25102 36196
rect 25777 36193 25789 36196
rect 25823 36193 25835 36227
rect 25777 36187 25835 36193
rect 24857 36159 24915 36165
rect 24857 36156 24869 36159
rect 23308 36128 24869 36156
rect 23201 36119 23259 36125
rect 24857 36125 24869 36128
rect 24903 36125 24915 36159
rect 24857 36119 24915 36125
rect 22094 36088 22100 36100
rect 22020 36060 22100 36088
rect 22094 36048 22100 36060
rect 22152 36048 22158 36100
rect 22738 36048 22744 36100
rect 22796 36088 22802 36100
rect 24765 36091 24823 36097
rect 24765 36088 24777 36091
rect 22796 36060 24777 36088
rect 22796 36048 22802 36060
rect 24765 36057 24777 36060
rect 24811 36057 24823 36091
rect 24765 36051 24823 36057
rect 25590 36048 25596 36100
rect 25648 36048 25654 36100
rect 15396 35992 16620 36020
rect 17678 35980 17684 36032
rect 17736 36020 17742 36032
rect 18598 36020 18604 36032
rect 17736 35992 18604 36020
rect 17736 35980 17742 35992
rect 18598 35980 18604 35992
rect 18656 35980 18662 36032
rect 18785 36023 18843 36029
rect 18785 35989 18797 36023
rect 18831 36020 18843 36023
rect 18966 36020 18972 36032
rect 18831 35992 18972 36020
rect 18831 35989 18843 35992
rect 18785 35983 18843 35989
rect 18966 35980 18972 35992
rect 19024 35980 19030 36032
rect 19242 35980 19248 36032
rect 19300 36020 19306 36032
rect 19613 36023 19671 36029
rect 19613 36020 19625 36023
rect 19300 35992 19625 36020
rect 19300 35980 19306 35992
rect 19613 35989 19625 35992
rect 19659 35989 19671 36023
rect 19613 35983 19671 35989
rect 21542 35980 21548 36032
rect 21600 36020 21606 36032
rect 22005 36023 22063 36029
rect 22005 36020 22017 36023
rect 21600 35992 22017 36020
rect 21600 35980 21606 35992
rect 22005 35989 22017 35992
rect 22051 35989 22063 36023
rect 22005 35983 22063 35989
rect 22465 36023 22523 36029
rect 22465 35989 22477 36023
rect 22511 36020 22523 36023
rect 22646 36020 22652 36032
rect 22511 35992 22652 36020
rect 22511 35989 22523 35992
rect 22465 35983 22523 35989
rect 22646 35980 22652 35992
rect 22704 35980 22710 36032
rect 23290 35980 23296 36032
rect 23348 35980 23354 36032
rect 23382 35980 23388 36032
rect 23440 36020 23446 36032
rect 25685 36023 25743 36029
rect 25685 36020 25697 36023
rect 23440 35992 25697 36020
rect 23440 35980 23446 35992
rect 25685 35989 25697 35992
rect 25731 35989 25743 36023
rect 25685 35983 25743 35989
rect 1104 35930 36432 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 36432 35930
rect 1104 35856 36432 35878
rect 8294 35816 8300 35828
rect 6472 35788 8300 35816
rect 6472 35748 6500 35788
rect 8294 35776 8300 35788
rect 8352 35776 8358 35828
rect 8404 35788 10364 35816
rect 6380 35720 6500 35748
rect 6380 35689 6408 35720
rect 7926 35708 7932 35760
rect 7984 35748 7990 35760
rect 8404 35748 8432 35788
rect 9674 35748 9680 35760
rect 7984 35720 8432 35748
rect 9048 35720 9680 35748
rect 7984 35708 7990 35720
rect 6365 35683 6423 35689
rect 6365 35649 6377 35683
rect 6411 35649 6423 35683
rect 6365 35643 6423 35649
rect 6641 35615 6699 35621
rect 6641 35581 6653 35615
rect 6687 35612 6699 35615
rect 6730 35612 6736 35624
rect 6687 35584 6736 35612
rect 6687 35581 6699 35584
rect 6641 35575 6699 35581
rect 6730 35572 6736 35584
rect 6788 35572 6794 35624
rect 7760 35612 7788 35666
rect 8754 35640 8760 35692
rect 8812 35640 8818 35692
rect 8938 35640 8944 35692
rect 8996 35640 9002 35692
rect 9048 35612 9076 35720
rect 9674 35708 9680 35720
rect 9732 35708 9738 35760
rect 10336 35748 10364 35788
rect 10410 35776 10416 35828
rect 10468 35816 10474 35828
rect 10505 35819 10563 35825
rect 10505 35816 10517 35819
rect 10468 35788 10517 35816
rect 10468 35776 10474 35788
rect 10505 35785 10517 35788
rect 10551 35785 10563 35819
rect 10505 35779 10563 35785
rect 11054 35776 11060 35828
rect 11112 35816 11118 35828
rect 11517 35819 11575 35825
rect 11517 35816 11529 35819
rect 11112 35788 11529 35816
rect 11112 35776 11118 35788
rect 11517 35785 11529 35788
rect 11563 35785 11575 35819
rect 11517 35779 11575 35785
rect 11885 35819 11943 35825
rect 11885 35785 11897 35819
rect 11931 35816 11943 35819
rect 12434 35816 12440 35828
rect 11931 35788 12440 35816
rect 11931 35785 11943 35788
rect 11885 35779 11943 35785
rect 12434 35776 12440 35788
rect 12492 35776 12498 35828
rect 12713 35819 12771 35825
rect 12713 35785 12725 35819
rect 12759 35816 12771 35819
rect 12802 35816 12808 35828
rect 12759 35788 12808 35816
rect 12759 35785 12771 35788
rect 12713 35779 12771 35785
rect 12802 35776 12808 35788
rect 12860 35776 12866 35828
rect 12894 35776 12900 35828
rect 12952 35816 12958 35828
rect 14461 35819 14519 35825
rect 14461 35816 14473 35819
rect 12952 35788 14473 35816
rect 12952 35776 12958 35788
rect 14461 35785 14473 35788
rect 14507 35785 14519 35819
rect 14461 35779 14519 35785
rect 14921 35819 14979 35825
rect 14921 35785 14933 35819
rect 14967 35816 14979 35819
rect 15286 35816 15292 35828
rect 14967 35788 15292 35816
rect 14967 35785 14979 35788
rect 14921 35779 14979 35785
rect 15286 35776 15292 35788
rect 15344 35776 15350 35828
rect 15470 35776 15476 35828
rect 15528 35816 15534 35828
rect 15841 35819 15899 35825
rect 15528 35788 15792 35816
rect 15528 35776 15534 35788
rect 13354 35748 13360 35760
rect 9968 35720 10272 35748
rect 9217 35683 9275 35689
rect 9217 35649 9229 35683
rect 9263 35680 9275 35683
rect 9263 35652 9720 35680
rect 9263 35649 9275 35652
rect 9217 35643 9275 35649
rect 7760 35584 9076 35612
rect 9125 35615 9183 35621
rect 9125 35581 9137 35615
rect 9171 35581 9183 35615
rect 9125 35575 9183 35581
rect 7650 35504 7656 35556
rect 7708 35544 7714 35556
rect 7708 35516 8892 35544
rect 7708 35504 7714 35516
rect 6822 35436 6828 35488
rect 6880 35476 6886 35488
rect 8113 35479 8171 35485
rect 8113 35476 8125 35479
rect 6880 35448 8125 35476
rect 6880 35436 6886 35448
rect 8113 35445 8125 35448
rect 8159 35445 8171 35479
rect 8113 35439 8171 35445
rect 8570 35436 8576 35488
rect 8628 35476 8634 35488
rect 8757 35479 8815 35485
rect 8757 35476 8769 35479
rect 8628 35448 8769 35476
rect 8628 35436 8634 35448
rect 8757 35445 8769 35448
rect 8803 35445 8815 35479
rect 8864 35476 8892 35516
rect 8938 35504 8944 35556
rect 8996 35544 9002 35556
rect 9140 35544 9168 35575
rect 9582 35572 9588 35624
rect 9640 35572 9646 35624
rect 9692 35612 9720 35652
rect 9766 35640 9772 35692
rect 9824 35640 9830 35692
rect 9968 35689 9996 35720
rect 9953 35683 10011 35689
rect 9953 35649 9965 35683
rect 9999 35649 10011 35683
rect 9953 35643 10011 35649
rect 10134 35640 10140 35692
rect 10192 35640 10198 35692
rect 10045 35615 10103 35621
rect 10045 35612 10057 35615
rect 9692 35584 10057 35612
rect 10045 35581 10057 35584
rect 10091 35581 10103 35615
rect 10244 35612 10272 35720
rect 10336 35720 12480 35748
rect 10336 35689 10364 35720
rect 10321 35683 10379 35689
rect 10321 35649 10333 35683
rect 10367 35649 10379 35683
rect 10321 35643 10379 35649
rect 10870 35640 10876 35692
rect 10928 35640 10934 35692
rect 12345 35683 12403 35689
rect 12345 35649 12357 35683
rect 12391 35649 12403 35683
rect 12345 35643 12403 35649
rect 10778 35612 10784 35624
rect 10244 35584 10784 35612
rect 10045 35575 10103 35581
rect 8996 35516 9168 35544
rect 10060 35544 10088 35575
rect 10778 35572 10784 35584
rect 10836 35572 10842 35624
rect 10962 35572 10968 35624
rect 11020 35572 11026 35624
rect 11974 35572 11980 35624
rect 12032 35572 12038 35624
rect 12069 35615 12127 35621
rect 12069 35581 12081 35615
rect 12115 35612 12127 35615
rect 12360 35612 12388 35643
rect 12115 35584 12388 35612
rect 12115 35581 12127 35584
rect 12069 35575 12127 35581
rect 11054 35544 11060 35556
rect 10060 35516 11060 35544
rect 8996 35504 9002 35516
rect 11054 35504 11060 35516
rect 11112 35504 11118 35556
rect 11422 35504 11428 35556
rect 11480 35544 11486 35556
rect 12084 35544 12112 35575
rect 11480 35516 12112 35544
rect 12452 35544 12480 35720
rect 12912 35720 13360 35748
rect 12912 35692 12940 35720
rect 13354 35708 13360 35720
rect 13412 35748 13418 35760
rect 15764 35748 15792 35788
rect 15841 35785 15853 35819
rect 15887 35816 15899 35819
rect 16482 35816 16488 35828
rect 15887 35788 16488 35816
rect 15887 35785 15899 35788
rect 15841 35779 15899 35785
rect 16482 35776 16488 35788
rect 16540 35776 16546 35828
rect 18141 35819 18199 35825
rect 18141 35785 18153 35819
rect 18187 35816 18199 35819
rect 18230 35816 18236 35828
rect 18187 35788 18236 35816
rect 18187 35785 18199 35788
rect 18141 35779 18199 35785
rect 18230 35776 18236 35788
rect 18288 35776 18294 35828
rect 21453 35819 21511 35825
rect 21453 35785 21465 35819
rect 21499 35816 21511 35819
rect 22554 35816 22560 35828
rect 21499 35788 22560 35816
rect 21499 35785 21511 35788
rect 21453 35779 21511 35785
rect 22554 35776 22560 35788
rect 22612 35776 22618 35828
rect 24489 35819 24547 35825
rect 24489 35816 24501 35819
rect 22664 35788 24501 35816
rect 13412 35720 14136 35748
rect 13412 35708 13418 35720
rect 12529 35683 12587 35689
rect 12529 35649 12541 35683
rect 12575 35680 12587 35683
rect 12802 35680 12808 35692
rect 12575 35652 12808 35680
rect 12575 35649 12587 35652
rect 12529 35643 12587 35649
rect 12802 35640 12808 35652
rect 12860 35640 12866 35692
rect 12894 35640 12900 35692
rect 12952 35640 12958 35692
rect 12986 35640 12992 35692
rect 13044 35640 13050 35692
rect 13538 35640 13544 35692
rect 13596 35640 13602 35692
rect 13998 35680 14004 35692
rect 13648 35652 14004 35680
rect 12820 35612 12848 35640
rect 13170 35612 13176 35624
rect 12820 35584 13176 35612
rect 13170 35572 13176 35584
rect 13228 35572 13234 35624
rect 13262 35572 13268 35624
rect 13320 35572 13326 35624
rect 13357 35615 13415 35621
rect 13357 35581 13369 35615
rect 13403 35612 13415 35615
rect 13648 35612 13676 35652
rect 13998 35640 14004 35652
rect 14056 35640 14062 35692
rect 14108 35689 14136 35720
rect 14844 35720 15700 35748
rect 15764 35720 16988 35748
rect 14844 35692 14872 35720
rect 14093 35683 14151 35689
rect 14093 35649 14105 35683
rect 14139 35649 14151 35683
rect 14093 35643 14151 35649
rect 14366 35640 14372 35692
rect 14424 35640 14430 35692
rect 14553 35683 14611 35689
rect 14553 35649 14565 35683
rect 14599 35649 14611 35683
rect 14553 35643 14611 35649
rect 13817 35615 13875 35621
rect 13817 35612 13829 35615
rect 13403 35584 13676 35612
rect 13740 35584 13829 35612
rect 13403 35581 13415 35584
rect 13357 35575 13415 35581
rect 13078 35544 13084 35556
rect 12452 35516 13084 35544
rect 11480 35504 11486 35516
rect 13078 35504 13084 35516
rect 13136 35504 13142 35556
rect 10226 35476 10232 35488
rect 8864 35448 10232 35476
rect 8757 35439 8815 35445
rect 10226 35436 10232 35448
rect 10284 35436 10290 35488
rect 11149 35479 11207 35485
rect 11149 35445 11161 35479
rect 11195 35476 11207 35479
rect 11606 35476 11612 35488
rect 11195 35448 11612 35476
rect 11195 35445 11207 35448
rect 11149 35439 11207 35445
rect 11606 35436 11612 35448
rect 11664 35436 11670 35488
rect 13170 35436 13176 35488
rect 13228 35436 13234 35488
rect 13630 35436 13636 35488
rect 13688 35476 13694 35488
rect 13740 35485 13768 35584
rect 13817 35581 13829 35584
rect 13863 35581 13875 35615
rect 14568 35612 14596 35643
rect 14826 35640 14832 35692
rect 14884 35640 14890 35692
rect 14918 35640 14924 35692
rect 14976 35680 14982 35692
rect 15013 35683 15071 35689
rect 15013 35680 15025 35683
rect 14976 35652 15025 35680
rect 14976 35640 14982 35652
rect 15013 35649 15025 35652
rect 15059 35649 15071 35683
rect 15013 35643 15071 35649
rect 15102 35640 15108 35692
rect 15160 35640 15166 35692
rect 15194 35640 15200 35692
rect 15252 35680 15258 35692
rect 15672 35689 15700 35720
rect 15289 35683 15347 35689
rect 15289 35680 15301 35683
rect 15252 35652 15301 35680
rect 15252 35640 15258 35652
rect 15289 35649 15301 35652
rect 15335 35649 15347 35683
rect 15289 35643 15347 35649
rect 15657 35683 15715 35689
rect 15657 35649 15669 35683
rect 15703 35649 15715 35683
rect 15657 35643 15715 35649
rect 16114 35640 16120 35692
rect 16172 35640 16178 35692
rect 16666 35640 16672 35692
rect 16724 35640 16730 35692
rect 16960 35689 16988 35720
rect 17034 35708 17040 35760
rect 17092 35748 17098 35760
rect 17405 35751 17463 35757
rect 17092 35720 17264 35748
rect 17092 35708 17098 35720
rect 17236 35689 17264 35720
rect 17405 35717 17417 35751
rect 17451 35748 17463 35751
rect 18322 35748 18328 35760
rect 17451 35720 18328 35748
rect 17451 35717 17463 35720
rect 17405 35711 17463 35717
rect 18322 35708 18328 35720
rect 18380 35708 18386 35760
rect 18693 35751 18751 35757
rect 18693 35717 18705 35751
rect 18739 35748 18751 35751
rect 18782 35748 18788 35760
rect 18739 35720 18788 35748
rect 18739 35717 18751 35720
rect 18693 35711 18751 35717
rect 18782 35708 18788 35720
rect 18840 35708 18846 35760
rect 22664 35757 22692 35788
rect 24489 35785 24501 35788
rect 24535 35785 24547 35819
rect 24489 35779 24547 35785
rect 22649 35751 22707 35757
rect 22649 35717 22661 35751
rect 22695 35717 22707 35751
rect 24949 35751 25007 35757
rect 24949 35748 24961 35751
rect 22649 35711 22707 35717
rect 24504 35720 24961 35748
rect 24504 35692 24532 35720
rect 24949 35717 24961 35720
rect 24995 35717 25007 35751
rect 24949 35711 25007 35717
rect 16853 35683 16911 35689
rect 16853 35649 16865 35683
rect 16899 35649 16911 35683
rect 16853 35643 16911 35649
rect 16945 35683 17003 35689
rect 16945 35649 16957 35683
rect 16991 35649 17003 35683
rect 16945 35643 17003 35649
rect 17221 35683 17279 35689
rect 17221 35649 17233 35683
rect 17267 35649 17279 35683
rect 17221 35643 17279 35649
rect 13817 35575 13875 35581
rect 14292 35584 14596 35612
rect 14292 35488 14320 35584
rect 15378 35572 15384 35624
rect 15436 35572 15442 35624
rect 15473 35615 15531 35621
rect 15473 35581 15485 35615
rect 15519 35581 15531 35615
rect 15473 35575 15531 35581
rect 16209 35615 16267 35621
rect 16209 35581 16221 35615
rect 16255 35612 16267 35615
rect 16298 35612 16304 35624
rect 16255 35584 16304 35612
rect 16255 35581 16267 35584
rect 16209 35575 16267 35581
rect 14642 35504 14648 35556
rect 14700 35544 14706 35556
rect 15488 35544 15516 35575
rect 16298 35572 16304 35584
rect 16356 35572 16362 35624
rect 16574 35572 16580 35624
rect 16632 35612 16638 35624
rect 16868 35612 16896 35643
rect 17770 35640 17776 35692
rect 17828 35640 17834 35692
rect 18414 35640 18420 35692
rect 18472 35640 18478 35692
rect 20346 35680 20352 35692
rect 19826 35652 20352 35680
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 20901 35683 20959 35689
rect 20901 35649 20913 35683
rect 20947 35649 20959 35683
rect 20901 35643 20959 35649
rect 16632 35584 16896 35612
rect 17037 35615 17095 35621
rect 16632 35572 16638 35584
rect 17037 35581 17049 35615
rect 17083 35612 17095 35615
rect 17402 35612 17408 35624
rect 17083 35584 17408 35612
rect 17083 35581 17095 35584
rect 17037 35575 17095 35581
rect 17052 35544 17080 35575
rect 17402 35572 17408 35584
rect 17460 35572 17466 35624
rect 17678 35572 17684 35624
rect 17736 35572 17742 35624
rect 17862 35572 17868 35624
rect 17920 35612 17926 35624
rect 20441 35615 20499 35621
rect 20441 35612 20453 35615
rect 17920 35584 20453 35612
rect 17920 35572 17926 35584
rect 20441 35581 20453 35584
rect 20487 35581 20499 35615
rect 20441 35575 20499 35581
rect 20916 35544 20944 35643
rect 21358 35640 21364 35692
rect 21416 35640 21422 35692
rect 23934 35680 23940 35692
rect 23782 35652 23940 35680
rect 23934 35640 23940 35652
rect 23992 35640 23998 35692
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35680 24455 35683
rect 24486 35680 24492 35692
rect 24443 35652 24492 35680
rect 24443 35649 24455 35652
rect 24397 35643 24455 35649
rect 24486 35640 24492 35652
rect 24544 35640 24550 35692
rect 24854 35640 24860 35692
rect 24912 35640 24918 35692
rect 26418 35680 26424 35692
rect 24964 35652 26424 35680
rect 20993 35615 21051 35621
rect 20993 35581 21005 35615
rect 21039 35581 21051 35615
rect 20993 35575 21051 35581
rect 14700 35516 17080 35544
rect 19720 35516 20944 35544
rect 21008 35544 21036 35575
rect 21082 35572 21088 35624
rect 21140 35612 21146 35624
rect 22186 35612 22192 35624
rect 21140 35584 22192 35612
rect 21140 35572 21146 35584
rect 22186 35572 22192 35584
rect 22244 35572 22250 35624
rect 22278 35572 22284 35624
rect 22336 35612 22342 35624
rect 22373 35615 22431 35621
rect 22373 35612 22385 35615
rect 22336 35584 22385 35612
rect 22336 35572 22342 35584
rect 22373 35581 22385 35584
rect 22419 35581 22431 35615
rect 22373 35575 22431 35581
rect 22646 35572 22652 35624
rect 22704 35612 22710 35624
rect 23014 35612 23020 35624
rect 22704 35584 23020 35612
rect 22704 35572 22710 35584
rect 23014 35572 23020 35584
rect 23072 35612 23078 35624
rect 24964 35612 24992 35652
rect 26418 35640 26424 35652
rect 26476 35640 26482 35692
rect 23072 35584 24992 35612
rect 23072 35572 23078 35584
rect 25038 35572 25044 35624
rect 25096 35572 25102 35624
rect 21634 35544 21640 35556
rect 21008 35516 21640 35544
rect 14700 35504 14706 35516
rect 13725 35479 13783 35485
rect 13725 35476 13737 35479
rect 13688 35448 13737 35476
rect 13688 35436 13694 35448
rect 13725 35445 13737 35448
rect 13771 35445 13783 35479
rect 13725 35439 13783 35445
rect 13906 35436 13912 35488
rect 13964 35436 13970 35488
rect 14274 35436 14280 35488
rect 14332 35436 14338 35488
rect 16393 35479 16451 35485
rect 16393 35445 16405 35479
rect 16439 35476 16451 35479
rect 16482 35476 16488 35488
rect 16439 35448 16488 35476
rect 16439 35445 16451 35448
rect 16393 35439 16451 35445
rect 16482 35436 16488 35448
rect 16540 35436 16546 35488
rect 16574 35436 16580 35488
rect 16632 35476 16638 35488
rect 19720 35476 19748 35516
rect 21634 35504 21640 35516
rect 21692 35504 21698 35556
rect 16632 35448 19748 35476
rect 16632 35436 16638 35448
rect 19886 35436 19892 35488
rect 19944 35476 19950 35488
rect 20533 35479 20591 35485
rect 20533 35476 20545 35479
rect 19944 35448 20545 35476
rect 19944 35436 19950 35448
rect 20533 35445 20545 35448
rect 20579 35445 20591 35479
rect 20533 35439 20591 35445
rect 1104 35386 36432 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 36432 35386
rect 1104 35312 36432 35334
rect 5994 35232 6000 35284
rect 6052 35232 6058 35284
rect 6730 35232 6736 35284
rect 6788 35232 6794 35284
rect 7834 35232 7840 35284
rect 7892 35272 7898 35284
rect 8202 35272 8208 35284
rect 7892 35244 8208 35272
rect 7892 35232 7898 35244
rect 8202 35232 8208 35244
rect 8260 35272 8266 35284
rect 8260 35244 8524 35272
rect 8260 35232 8266 35244
rect 7285 35207 7343 35213
rect 7285 35173 7297 35207
rect 7331 35204 7343 35207
rect 7374 35204 7380 35216
rect 7331 35176 7380 35204
rect 7331 35173 7343 35176
rect 7285 35167 7343 35173
rect 7374 35164 7380 35176
rect 7432 35164 7438 35216
rect 8496 35213 8524 35244
rect 8754 35232 8760 35284
rect 8812 35272 8818 35284
rect 8941 35275 8999 35281
rect 8941 35272 8953 35275
rect 8812 35244 8953 35272
rect 8812 35232 8818 35244
rect 8941 35241 8953 35244
rect 8987 35241 8999 35275
rect 8941 35235 8999 35241
rect 9306 35232 9312 35284
rect 9364 35232 9370 35284
rect 10505 35275 10563 35281
rect 10505 35241 10517 35275
rect 10551 35272 10563 35275
rect 10870 35272 10876 35284
rect 10551 35244 10876 35272
rect 10551 35241 10563 35244
rect 10505 35235 10563 35241
rect 10870 35232 10876 35244
rect 10928 35232 10934 35284
rect 11974 35232 11980 35284
rect 12032 35232 12038 35284
rect 13357 35275 13415 35281
rect 13357 35241 13369 35275
rect 13403 35272 13415 35275
rect 14366 35272 14372 35284
rect 13403 35244 14372 35272
rect 13403 35241 13415 35244
rect 13357 35235 13415 35241
rect 14366 35232 14372 35244
rect 14424 35232 14430 35284
rect 15102 35232 15108 35284
rect 15160 35272 15166 35284
rect 15565 35275 15623 35281
rect 15565 35272 15577 35275
rect 15160 35244 15577 35272
rect 15160 35232 15166 35244
rect 15565 35241 15577 35244
rect 15611 35241 15623 35275
rect 15565 35235 15623 35241
rect 16298 35232 16304 35284
rect 16356 35272 16362 35284
rect 17402 35272 17408 35284
rect 16356 35244 17408 35272
rect 16356 35232 16362 35244
rect 17402 35232 17408 35244
rect 17460 35232 17466 35284
rect 17770 35232 17776 35284
rect 17828 35272 17834 35284
rect 17865 35275 17923 35281
rect 17865 35272 17877 35275
rect 17828 35244 17877 35272
rect 17828 35232 17834 35244
rect 17865 35241 17877 35244
rect 17911 35241 17923 35275
rect 17865 35235 17923 35241
rect 21634 35232 21640 35284
rect 21692 35272 21698 35284
rect 27062 35272 27068 35284
rect 21692 35244 27068 35272
rect 21692 35232 21698 35244
rect 27062 35232 27068 35244
rect 27120 35232 27126 35284
rect 8481 35207 8539 35213
rect 8481 35173 8493 35207
rect 8527 35173 8539 35207
rect 9324 35204 9352 35232
rect 8481 35167 8539 35173
rect 8588 35176 9352 35204
rect 6822 35136 6828 35148
rect 5828 35108 6828 35136
rect 5828 35077 5856 35108
rect 6472 35080 6500 35108
rect 6822 35096 6828 35108
rect 6880 35136 6886 35148
rect 7469 35139 7527 35145
rect 7469 35136 7481 35139
rect 6880 35108 7481 35136
rect 6880 35096 6886 35108
rect 7469 35105 7481 35108
rect 7515 35105 7527 35139
rect 8588 35136 8616 35176
rect 10962 35164 10968 35216
rect 11020 35204 11026 35216
rect 11149 35207 11207 35213
rect 11149 35204 11161 35207
rect 11020 35176 11161 35204
rect 11020 35164 11026 35176
rect 11149 35173 11161 35176
rect 11195 35204 11207 35207
rect 13265 35207 13323 35213
rect 11195 35176 12296 35204
rect 11195 35173 11207 35176
rect 11149 35167 11207 35173
rect 7469 35099 7527 35105
rect 8128 35108 8616 35136
rect 5813 35071 5871 35077
rect 5813 35037 5825 35071
rect 5859 35037 5871 35071
rect 5813 35031 5871 35037
rect 5997 35071 6055 35077
rect 5997 35037 6009 35071
rect 6043 35037 6055 35071
rect 5997 35031 6055 35037
rect 6012 34932 6040 35031
rect 6086 35028 6092 35080
rect 6144 35028 6150 35080
rect 6270 35028 6276 35080
rect 6328 35028 6334 35080
rect 6362 35028 6368 35080
rect 6420 35028 6426 35080
rect 6454 35028 6460 35080
rect 6512 35028 6518 35080
rect 7098 35028 7104 35080
rect 7156 35028 7162 35080
rect 7282 35028 7288 35080
rect 7340 35068 7346 35080
rect 7377 35071 7435 35077
rect 7377 35068 7389 35071
rect 7340 35040 7389 35068
rect 7340 35028 7346 35040
rect 7377 35037 7389 35040
rect 7423 35037 7435 35071
rect 7377 35031 7435 35037
rect 7650 35028 7656 35080
rect 7708 35028 7714 35080
rect 7926 35028 7932 35080
rect 7984 35077 7990 35080
rect 8128 35077 8156 35108
rect 9030 35096 9036 35148
rect 9088 35136 9094 35148
rect 9217 35139 9275 35145
rect 9217 35136 9229 35139
rect 9088 35108 9229 35136
rect 9088 35096 9094 35108
rect 9217 35105 9229 35108
rect 9263 35105 9275 35139
rect 10873 35139 10931 35145
rect 10873 35136 10885 35139
rect 9217 35099 9275 35105
rect 10244 35108 10885 35136
rect 10244 35080 10272 35108
rect 10873 35105 10885 35108
rect 10919 35105 10931 35139
rect 10873 35099 10931 35105
rect 11330 35096 11336 35148
rect 11388 35096 11394 35148
rect 7984 35068 7993 35077
rect 8113 35071 8171 35077
rect 7984 35040 8029 35068
rect 7984 35031 7993 35040
rect 8113 35037 8125 35071
rect 8159 35037 8171 35071
rect 8113 35031 8171 35037
rect 8297 35071 8355 35077
rect 8297 35037 8309 35071
rect 8343 35037 8355 35071
rect 8297 35031 8355 35037
rect 8389 35071 8447 35077
rect 8389 35037 8401 35071
rect 8435 35037 8447 35071
rect 8389 35031 8447 35037
rect 7984 35028 7990 35031
rect 7668 35000 7696 35028
rect 6472 34972 7696 35000
rect 8021 35003 8079 35009
rect 6472 34932 6500 34972
rect 8021 34969 8033 35003
rect 8067 35000 8079 35003
rect 8312 35000 8340 35031
rect 8067 34972 8340 35000
rect 8067 34969 8079 34972
rect 8021 34963 8079 34969
rect 6012 34904 6500 34932
rect 6917 34935 6975 34941
rect 6917 34901 6929 34935
rect 6963 34932 6975 34935
rect 7006 34932 7012 34944
rect 6963 34904 7012 34932
rect 6963 34901 6975 34904
rect 6917 34895 6975 34901
rect 7006 34892 7012 34904
rect 7064 34932 7070 34944
rect 8404 34932 8432 35031
rect 8570 35028 8576 35080
rect 8628 35028 8634 35080
rect 8938 35028 8944 35080
rect 8996 35028 9002 35080
rect 9125 35071 9183 35077
rect 9125 35037 9137 35071
rect 9171 35037 9183 35071
rect 9125 35031 9183 35037
rect 9493 35071 9551 35077
rect 9493 35037 9505 35071
rect 9539 35068 9551 35071
rect 9582 35068 9588 35080
rect 9539 35040 9588 35068
rect 9539 35037 9551 35040
rect 9493 35031 9551 35037
rect 8846 34960 8852 35012
rect 8904 35000 8910 35012
rect 9140 35000 9168 35031
rect 9582 35028 9588 35040
rect 9640 35028 9646 35080
rect 10226 35028 10232 35080
rect 10284 35028 10290 35080
rect 10686 35028 10692 35080
rect 10744 35068 10750 35080
rect 10781 35071 10839 35077
rect 10781 35068 10793 35071
rect 10744 35040 10793 35068
rect 10744 35028 10750 35040
rect 10781 35037 10793 35040
rect 10827 35037 10839 35071
rect 10781 35031 10839 35037
rect 10962 35028 10968 35080
rect 11020 35068 11026 35080
rect 11422 35068 11428 35080
rect 11020 35040 11428 35068
rect 11020 35028 11026 35040
rect 11422 35028 11428 35040
rect 11480 35028 11486 35080
rect 11514 35028 11520 35080
rect 11572 35028 11578 35080
rect 11606 35028 11612 35080
rect 11664 35028 11670 35080
rect 12268 35077 12296 35176
rect 13265 35173 13277 35207
rect 13311 35204 13323 35207
rect 13630 35204 13636 35216
rect 13311 35176 13636 35204
rect 13311 35173 13323 35176
rect 13265 35167 13323 35173
rect 13630 35164 13636 35176
rect 13688 35164 13694 35216
rect 13725 35207 13783 35213
rect 13725 35173 13737 35207
rect 13771 35204 13783 35207
rect 14182 35204 14188 35216
rect 13771 35176 14188 35204
rect 13771 35173 13783 35176
rect 13725 35167 13783 35173
rect 14182 35164 14188 35176
rect 14240 35164 14246 35216
rect 14918 35164 14924 35216
rect 14976 35204 14982 35216
rect 16853 35207 16911 35213
rect 16853 35204 16865 35207
rect 14976 35176 16865 35204
rect 14976 35164 14982 35176
rect 16853 35173 16865 35176
rect 16899 35204 16911 35207
rect 17586 35204 17592 35216
rect 16899 35176 17592 35204
rect 16899 35173 16911 35176
rect 16853 35167 16911 35173
rect 17586 35164 17592 35176
rect 17644 35204 17650 35216
rect 18690 35204 18696 35216
rect 17644 35176 18696 35204
rect 17644 35164 17650 35176
rect 18690 35164 18696 35176
rect 18748 35164 18754 35216
rect 12894 35096 12900 35148
rect 12952 35136 12958 35148
rect 13081 35139 13139 35145
rect 13081 35136 13093 35139
rect 12952 35108 13093 35136
rect 12952 35096 12958 35108
rect 13081 35105 13093 35108
rect 13127 35105 13139 35139
rect 13081 35099 13139 35105
rect 13170 35096 13176 35148
rect 13228 35136 13234 35148
rect 13228 35108 13492 35136
rect 13228 35096 13234 35108
rect 13464 35077 13492 35108
rect 13998 35096 14004 35148
rect 14056 35136 14062 35148
rect 14550 35136 14556 35148
rect 14056 35108 14556 35136
rect 14056 35096 14062 35108
rect 14550 35096 14556 35108
rect 14608 35096 14614 35148
rect 15105 35139 15163 35145
rect 14660 35108 14964 35136
rect 12069 35071 12127 35077
rect 12069 35037 12081 35071
rect 12115 35037 12127 35071
rect 12069 35031 12127 35037
rect 12253 35071 12311 35077
rect 12253 35037 12265 35071
rect 12299 35037 12311 35071
rect 12253 35031 12311 35037
rect 12437 35071 12495 35077
rect 12437 35037 12449 35071
rect 12483 35068 12495 35071
rect 13357 35071 13415 35077
rect 13357 35068 13369 35071
rect 12483 35040 13369 35068
rect 12483 35037 12495 35040
rect 12437 35031 12495 35037
rect 13357 35037 13369 35040
rect 13403 35037 13415 35071
rect 13357 35031 13415 35037
rect 13449 35071 13507 35077
rect 13449 35037 13461 35071
rect 13495 35037 13507 35071
rect 13449 35031 13507 35037
rect 13541 35071 13599 35077
rect 13541 35037 13553 35071
rect 13587 35068 13599 35071
rect 13906 35068 13912 35080
rect 13587 35040 13912 35068
rect 13587 35037 13599 35040
rect 13541 35031 13599 35037
rect 8904 34972 9168 35000
rect 9677 35003 9735 35009
rect 8904 34960 8910 34972
rect 9677 34969 9689 35003
rect 9723 35000 9735 35003
rect 9858 35000 9864 35012
rect 9723 34972 9864 35000
rect 9723 34969 9735 34972
rect 9677 34963 9735 34969
rect 9858 34960 9864 34972
rect 9916 35000 9922 35012
rect 10505 35003 10563 35009
rect 10505 35000 10517 35003
rect 9916 34972 10517 35000
rect 9916 34960 9922 34972
rect 10505 34969 10517 34972
rect 10551 35000 10563 35003
rect 12084 35000 12112 35031
rect 10551 34972 12112 35000
rect 13372 35000 13400 35031
rect 13556 35000 13584 35031
rect 13906 35028 13912 35040
rect 13964 35028 13970 35080
rect 14660 35077 14688 35108
rect 14936 35077 14964 35108
rect 15105 35105 15117 35139
rect 15151 35136 15163 35139
rect 15473 35139 15531 35145
rect 15473 35136 15485 35139
rect 15151 35108 15485 35136
rect 15151 35105 15163 35108
rect 15105 35099 15163 35105
rect 15473 35105 15485 35108
rect 15519 35105 15531 35139
rect 15473 35099 15531 35105
rect 17310 35096 17316 35148
rect 17368 35136 17374 35148
rect 17405 35139 17463 35145
rect 17405 35136 17417 35139
rect 17368 35108 17417 35136
rect 17368 35096 17374 35108
rect 17405 35105 17417 35108
rect 17451 35105 17463 35139
rect 17405 35099 17463 35105
rect 18325 35139 18383 35145
rect 18325 35105 18337 35139
rect 18371 35136 18383 35139
rect 18414 35136 18420 35148
rect 18371 35108 18420 35136
rect 18371 35105 18383 35108
rect 18325 35099 18383 35105
rect 18414 35096 18420 35108
rect 18472 35096 18478 35148
rect 19610 35096 19616 35148
rect 19668 35136 19674 35148
rect 20993 35139 21051 35145
rect 19668 35108 20300 35136
rect 19668 35096 19674 35108
rect 14645 35071 14703 35077
rect 14645 35037 14657 35071
rect 14691 35037 14703 35071
rect 14645 35031 14703 35037
rect 14829 35071 14887 35077
rect 14829 35037 14841 35071
rect 14875 35037 14887 35071
rect 14829 35031 14887 35037
rect 14921 35071 14979 35077
rect 14921 35037 14933 35071
rect 14967 35068 14979 35071
rect 15010 35068 15016 35080
rect 14967 35040 15016 35068
rect 14967 35037 14979 35040
rect 14921 35031 14979 35037
rect 13372 34972 13584 35000
rect 13725 35003 13783 35009
rect 10551 34969 10563 34972
rect 10505 34963 10563 34969
rect 13725 34969 13737 35003
rect 13771 35000 13783 35003
rect 14090 35000 14096 35012
rect 13771 34972 14096 35000
rect 13771 34969 13783 34972
rect 13725 34963 13783 34969
rect 14090 34960 14096 34972
rect 14148 34960 14154 35012
rect 14844 35000 14872 35031
rect 15010 35028 15016 35040
rect 15068 35028 15074 35080
rect 15378 35028 15384 35080
rect 15436 35068 15442 35080
rect 15657 35071 15715 35077
rect 15657 35068 15669 35071
rect 15436 35040 15669 35068
rect 15436 35028 15442 35040
rect 15657 35037 15669 35040
rect 15703 35037 15715 35071
rect 15657 35031 15715 35037
rect 15749 35071 15807 35077
rect 15749 35037 15761 35071
rect 15795 35068 15807 35071
rect 16209 35071 16267 35077
rect 15795 35040 16160 35068
rect 15795 35037 15807 35040
rect 15749 35031 15807 35037
rect 16025 35003 16083 35009
rect 16025 35000 16037 35003
rect 14844 34972 16037 35000
rect 16025 34969 16037 34972
rect 16071 34969 16083 35003
rect 16025 34963 16083 34969
rect 7064 34904 8432 34932
rect 7064 34892 7070 34904
rect 8754 34892 8760 34944
rect 8812 34892 8818 34944
rect 10321 34935 10379 34941
rect 10321 34901 10333 34935
rect 10367 34932 10379 34935
rect 11054 34932 11060 34944
rect 10367 34904 11060 34932
rect 10367 34901 10379 34904
rect 10321 34895 10379 34901
rect 11054 34892 11060 34904
rect 11112 34932 11118 34944
rect 12158 34932 12164 34944
rect 11112 34904 12164 34932
rect 11112 34892 11118 34904
rect 12158 34892 12164 34904
rect 12216 34932 12222 34944
rect 13998 34932 14004 34944
rect 12216 34904 14004 34932
rect 12216 34892 12222 34904
rect 13998 34892 14004 34904
rect 14056 34892 14062 34944
rect 14182 34892 14188 34944
rect 14240 34932 14246 34944
rect 14642 34932 14648 34944
rect 14240 34904 14648 34932
rect 14240 34892 14246 34904
rect 14642 34892 14648 34904
rect 14700 34892 14706 34944
rect 14734 34892 14740 34944
rect 14792 34892 14798 34944
rect 15286 34892 15292 34944
rect 15344 34932 15350 34944
rect 16132 34932 16160 35040
rect 16209 35037 16221 35071
rect 16255 35068 16267 35071
rect 16298 35068 16304 35080
rect 16255 35040 16304 35068
rect 16255 35037 16267 35040
rect 16209 35031 16267 35037
rect 16298 35028 16304 35040
rect 16356 35028 16362 35080
rect 16482 35028 16488 35080
rect 16540 35028 16546 35080
rect 16850 35028 16856 35080
rect 16908 35068 16914 35080
rect 17129 35071 17187 35077
rect 17129 35068 17141 35071
rect 16908 35040 17141 35068
rect 16908 35028 16914 35040
rect 17129 35037 17141 35040
rect 17175 35037 17187 35071
rect 17129 35031 17187 35037
rect 17497 35071 17555 35077
rect 17497 35037 17509 35071
rect 17543 35068 17555 35071
rect 17862 35068 17868 35080
rect 17543 35040 17868 35068
rect 17543 35037 17555 35040
rect 17497 35031 17555 35037
rect 16758 34960 16764 35012
rect 16816 35000 16822 35012
rect 17512 35000 17540 35031
rect 17862 35028 17868 35040
rect 17920 35028 17926 35080
rect 20272 35077 20300 35108
rect 20993 35105 21005 35139
rect 21039 35136 21051 35139
rect 22278 35136 22284 35148
rect 21039 35108 22284 35136
rect 21039 35105 21051 35108
rect 20993 35099 21051 35105
rect 22278 35096 22284 35108
rect 22336 35136 22342 35148
rect 23293 35139 23351 35145
rect 23293 35136 23305 35139
rect 22336 35108 23305 35136
rect 22336 35096 22342 35108
rect 23293 35105 23305 35108
rect 23339 35136 23351 35139
rect 23842 35136 23848 35148
rect 23339 35108 23848 35136
rect 23339 35105 23351 35108
rect 23293 35099 23351 35105
rect 23842 35096 23848 35108
rect 23900 35096 23906 35148
rect 19061 35071 19119 35077
rect 19061 35037 19073 35071
rect 19107 35068 19119 35071
rect 20257 35071 20315 35077
rect 19107 35040 20208 35068
rect 19107 35037 19119 35040
rect 19061 35031 19119 35037
rect 20180 35012 20208 35040
rect 20257 35037 20269 35071
rect 20303 35037 20315 35071
rect 20257 35031 20315 35037
rect 23014 35028 23020 35080
rect 23072 35028 23078 35080
rect 27249 35071 27307 35077
rect 27249 35037 27261 35071
rect 27295 35037 27307 35071
rect 27249 35031 27307 35037
rect 16816 34972 17540 35000
rect 19429 35003 19487 35009
rect 16816 34960 16822 34972
rect 19429 34969 19441 35003
rect 19475 35000 19487 35003
rect 19610 35000 19616 35012
rect 19475 34972 19616 35000
rect 19475 34969 19487 34972
rect 19429 34963 19487 34969
rect 19610 34960 19616 34972
rect 19668 34960 19674 35012
rect 20162 34960 20168 35012
rect 20220 34960 20226 35012
rect 21269 35003 21327 35009
rect 21269 34969 21281 35003
rect 21315 35000 21327 35003
rect 21542 35000 21548 35012
rect 21315 34972 21548 35000
rect 21315 34969 21327 34972
rect 21269 34963 21327 34969
rect 21542 34960 21548 34972
rect 21600 34960 21606 35012
rect 22554 35000 22560 35012
rect 22494 34972 22560 35000
rect 22554 34960 22560 34972
rect 22612 34960 22618 35012
rect 24029 35003 24087 35009
rect 24029 34969 24041 35003
rect 24075 34969 24087 35003
rect 24029 34963 24087 34969
rect 25133 35003 25191 35009
rect 25133 34969 25145 35003
rect 25179 35000 25191 35003
rect 25314 35000 25320 35012
rect 25179 34972 25320 35000
rect 25179 34969 25191 34972
rect 25133 34963 25191 34969
rect 15344 34904 16160 34932
rect 15344 34892 15350 34904
rect 16390 34892 16396 34944
rect 16448 34892 16454 34944
rect 20180 34932 20208 34960
rect 24044 34932 24072 34963
rect 25314 34960 25320 34972
rect 25372 34960 25378 35012
rect 25869 35003 25927 35009
rect 25869 34969 25881 35003
rect 25915 34969 25927 35003
rect 27264 35000 27292 35031
rect 27522 35028 27528 35080
rect 27580 35028 27586 35080
rect 27798 35000 27804 35012
rect 27264 34972 27804 35000
rect 25869 34963 25927 34969
rect 25884 34932 25912 34963
rect 27798 34960 27804 34972
rect 27856 34960 27862 35012
rect 20180 34904 25912 34932
rect 26602 34892 26608 34944
rect 26660 34932 26666 34944
rect 27065 34935 27123 34941
rect 27065 34932 27077 34935
rect 26660 34904 27077 34932
rect 26660 34892 26666 34904
rect 27065 34901 27077 34904
rect 27111 34901 27123 34935
rect 27065 34895 27123 34901
rect 27338 34892 27344 34944
rect 27396 34932 27402 34944
rect 27433 34935 27491 34941
rect 27433 34932 27445 34935
rect 27396 34904 27445 34932
rect 27396 34892 27402 34904
rect 27433 34901 27445 34904
rect 27479 34901 27491 34935
rect 27433 34895 27491 34901
rect 1104 34842 36432 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 36432 34842
rect 1104 34768 36432 34790
rect 6086 34688 6092 34740
rect 6144 34688 6150 34740
rect 6270 34688 6276 34740
rect 6328 34728 6334 34740
rect 6733 34731 6791 34737
rect 6733 34728 6745 34731
rect 6328 34700 6745 34728
rect 6328 34688 6334 34700
rect 6733 34697 6745 34700
rect 6779 34697 6791 34731
rect 7377 34731 7435 34737
rect 7377 34728 7389 34731
rect 6733 34691 6791 34697
rect 6932 34700 7389 34728
rect 5997 34595 6055 34601
rect 5997 34561 6009 34595
rect 6043 34561 6055 34595
rect 5997 34555 6055 34561
rect 5442 34484 5448 34536
rect 5500 34524 5506 34536
rect 6012 34524 6040 34555
rect 6178 34552 6184 34604
rect 6236 34552 6242 34604
rect 6825 34595 6883 34601
rect 6825 34561 6837 34595
rect 6871 34592 6883 34595
rect 6932 34592 6960 34700
rect 7377 34697 7389 34700
rect 7423 34697 7435 34731
rect 7377 34691 7435 34697
rect 7484 34700 8248 34728
rect 7098 34620 7104 34672
rect 7156 34620 7162 34672
rect 7484 34660 7512 34700
rect 7208 34632 7512 34660
rect 7561 34663 7619 34669
rect 6871 34564 6960 34592
rect 6871 34561 6883 34564
rect 6825 34555 6883 34561
rect 7006 34552 7012 34604
rect 7064 34592 7070 34604
rect 7208 34592 7236 34632
rect 7561 34629 7573 34663
rect 7607 34660 7619 34663
rect 8220 34660 8248 34700
rect 9030 34688 9036 34740
rect 9088 34728 9094 34740
rect 9217 34731 9275 34737
rect 9217 34728 9229 34731
rect 9088 34700 9229 34728
rect 9088 34688 9094 34700
rect 9217 34697 9229 34700
rect 9263 34697 9275 34731
rect 9217 34691 9275 34697
rect 9766 34688 9772 34740
rect 9824 34728 9830 34740
rect 9953 34731 10011 34737
rect 9953 34728 9965 34731
rect 9824 34700 9965 34728
rect 9824 34688 9830 34700
rect 9953 34697 9965 34700
rect 9999 34697 10011 34731
rect 9953 34691 10011 34697
rect 10686 34688 10692 34740
rect 10744 34728 10750 34740
rect 12434 34728 12440 34740
rect 10744 34700 12440 34728
rect 10744 34688 10750 34700
rect 12406 34688 12440 34700
rect 12492 34688 12498 34740
rect 12618 34688 12624 34740
rect 12676 34728 12682 34740
rect 12713 34731 12771 34737
rect 12713 34728 12725 34731
rect 12676 34700 12725 34728
rect 12676 34688 12682 34700
rect 12713 34697 12725 34700
rect 12759 34697 12771 34731
rect 12713 34691 12771 34697
rect 12802 34688 12808 34740
rect 12860 34728 12866 34740
rect 12897 34731 12955 34737
rect 12897 34728 12909 34731
rect 12860 34700 12909 34728
rect 12860 34688 12866 34700
rect 12897 34697 12909 34700
rect 12943 34728 12955 34731
rect 13906 34728 13912 34740
rect 12943 34700 13912 34728
rect 12943 34697 12955 34700
rect 12897 34691 12955 34697
rect 13906 34688 13912 34700
rect 13964 34688 13970 34740
rect 15197 34731 15255 34737
rect 15197 34697 15209 34731
rect 15243 34728 15255 34731
rect 15286 34728 15292 34740
rect 15243 34700 15292 34728
rect 15243 34697 15255 34700
rect 15197 34691 15255 34697
rect 15286 34688 15292 34700
rect 15344 34688 15350 34740
rect 16206 34688 16212 34740
rect 16264 34728 16270 34740
rect 16485 34731 16543 34737
rect 16485 34728 16497 34731
rect 16264 34700 16497 34728
rect 16264 34688 16270 34700
rect 16485 34697 16497 34700
rect 16531 34697 16543 34731
rect 16485 34691 16543 34697
rect 16666 34688 16672 34740
rect 16724 34688 16730 34740
rect 17402 34688 17408 34740
rect 17460 34688 17466 34740
rect 18233 34731 18291 34737
rect 18233 34697 18245 34731
rect 18279 34728 18291 34731
rect 19242 34728 19248 34740
rect 18279 34700 19248 34728
rect 18279 34697 18291 34700
rect 18233 34691 18291 34697
rect 19242 34688 19248 34700
rect 19300 34688 19306 34740
rect 22094 34728 22100 34740
rect 20272 34700 22100 34728
rect 8665 34663 8723 34669
rect 7607 34632 7788 34660
rect 8220 34632 8340 34660
rect 7607 34629 7619 34632
rect 7561 34623 7619 34629
rect 7064 34564 7236 34592
rect 7064 34552 7070 34564
rect 7282 34552 7288 34604
rect 7340 34552 7346 34604
rect 7374 34552 7380 34604
rect 7432 34552 7438 34604
rect 7466 34552 7472 34604
rect 7524 34552 7530 34604
rect 7650 34552 7656 34604
rect 7708 34552 7714 34604
rect 7760 34601 7788 34632
rect 7745 34595 7803 34601
rect 7745 34561 7757 34595
rect 7791 34561 7803 34595
rect 7745 34555 7803 34561
rect 7929 34595 7987 34601
rect 7929 34561 7941 34595
rect 7975 34561 7987 34595
rect 7929 34555 7987 34561
rect 7098 34524 7104 34536
rect 5500 34496 7104 34524
rect 5500 34484 5506 34496
rect 7098 34484 7104 34496
rect 7156 34484 7162 34536
rect 7300 34524 7328 34552
rect 7834 34524 7840 34536
rect 7300 34496 7840 34524
rect 7834 34484 7840 34496
rect 7892 34524 7898 34536
rect 7944 34524 7972 34555
rect 8202 34552 8208 34604
rect 8260 34552 8266 34604
rect 8312 34601 8340 34632
rect 8665 34629 8677 34663
rect 8711 34660 8723 34663
rect 9306 34660 9312 34672
rect 8711 34632 9312 34660
rect 8711 34629 8723 34632
rect 8665 34623 8723 34629
rect 9306 34620 9312 34632
rect 9364 34620 9370 34672
rect 9398 34620 9404 34672
rect 9456 34660 9462 34672
rect 12406 34660 12434 34688
rect 13081 34663 13139 34669
rect 9456 34632 10088 34660
rect 12406 34632 12940 34660
rect 9456 34620 9462 34632
rect 8297 34595 8355 34601
rect 8297 34561 8309 34595
rect 8343 34561 8355 34595
rect 8297 34555 8355 34561
rect 8481 34595 8539 34601
rect 8481 34561 8493 34595
rect 8527 34592 8539 34595
rect 8570 34592 8576 34604
rect 8527 34564 8576 34592
rect 8527 34561 8539 34564
rect 8481 34555 8539 34561
rect 8570 34552 8576 34564
rect 8628 34552 8634 34604
rect 8938 34552 8944 34604
rect 8996 34592 9002 34604
rect 9033 34595 9091 34601
rect 9033 34592 9045 34595
rect 8996 34564 9045 34592
rect 8996 34552 9002 34564
rect 9033 34561 9045 34564
rect 9079 34561 9091 34595
rect 9033 34555 9091 34561
rect 9858 34552 9864 34604
rect 9916 34552 9922 34604
rect 10060 34601 10088 34632
rect 10045 34595 10103 34601
rect 10045 34561 10057 34595
rect 10091 34592 10103 34595
rect 11330 34592 11336 34604
rect 10091 34564 11336 34592
rect 10091 34561 10103 34564
rect 10045 34555 10103 34561
rect 11330 34552 11336 34564
rect 11388 34552 11394 34604
rect 12158 34552 12164 34604
rect 12216 34592 12222 34604
rect 12253 34595 12311 34601
rect 12253 34592 12265 34595
rect 12216 34564 12265 34592
rect 12216 34552 12222 34564
rect 12253 34561 12265 34564
rect 12299 34561 12311 34595
rect 12253 34555 12311 34561
rect 12345 34595 12403 34601
rect 12345 34561 12357 34595
rect 12391 34592 12403 34595
rect 12434 34592 12440 34604
rect 12391 34564 12440 34592
rect 12391 34561 12403 34564
rect 12345 34555 12403 34561
rect 12434 34552 12440 34564
rect 12492 34552 12498 34604
rect 12526 34552 12532 34604
rect 12584 34552 12590 34604
rect 12805 34595 12863 34601
rect 12805 34561 12817 34595
rect 12851 34561 12863 34595
rect 12912 34592 12940 34632
rect 13081 34629 13093 34663
rect 13127 34660 13139 34663
rect 14274 34660 14280 34672
rect 13127 34632 14280 34660
rect 13127 34629 13139 34632
rect 13081 34623 13139 34629
rect 14274 34620 14280 34632
rect 14332 34620 14338 34672
rect 14734 34620 14740 34672
rect 14792 34660 14798 34672
rect 19337 34663 19395 34669
rect 19337 34660 19349 34663
rect 14792 34632 15976 34660
rect 14792 34620 14798 34632
rect 13262 34592 13268 34604
rect 12912 34564 13268 34592
rect 12805 34555 12863 34561
rect 7892 34496 7972 34524
rect 7892 34484 7898 34496
rect 8846 34484 8852 34536
rect 8904 34484 8910 34536
rect 11974 34484 11980 34536
rect 12032 34524 12038 34536
rect 12820 34524 12848 34555
rect 13262 34552 13268 34564
rect 13320 34592 13326 34604
rect 13630 34592 13636 34604
rect 13320 34564 13636 34592
rect 13320 34552 13326 34564
rect 13630 34552 13636 34564
rect 13688 34552 13694 34604
rect 15194 34552 15200 34604
rect 15252 34592 15258 34604
rect 15473 34595 15531 34601
rect 15473 34592 15485 34595
rect 15252 34564 15485 34592
rect 15252 34552 15258 34564
rect 15473 34561 15485 34564
rect 15519 34592 15531 34595
rect 15838 34592 15844 34604
rect 15519 34564 15844 34592
rect 15519 34561 15531 34564
rect 15473 34555 15531 34561
rect 15838 34552 15844 34564
rect 15896 34552 15902 34604
rect 15948 34592 15976 34632
rect 18064 34632 19349 34660
rect 18064 34604 18092 34632
rect 19337 34629 19349 34632
rect 19383 34629 19395 34663
rect 19337 34623 19395 34629
rect 19886 34620 19892 34672
rect 19944 34620 19950 34672
rect 20272 34660 20300 34700
rect 22094 34688 22100 34700
rect 22152 34728 22158 34740
rect 22281 34731 22339 34737
rect 22281 34728 22293 34731
rect 22152 34700 22293 34728
rect 22152 34688 22158 34700
rect 22281 34697 22293 34700
rect 22327 34728 22339 34731
rect 22554 34728 22560 34740
rect 22327 34700 22560 34728
rect 22327 34697 22339 34700
rect 22281 34691 22339 34697
rect 22554 34688 22560 34700
rect 22612 34688 22618 34740
rect 23566 34728 23572 34740
rect 23216 34700 23572 34728
rect 20346 34660 20352 34672
rect 20272 34632 20352 34660
rect 20346 34620 20352 34632
rect 20404 34620 20410 34672
rect 21634 34620 21640 34672
rect 21692 34620 21698 34672
rect 22373 34663 22431 34669
rect 22373 34629 22385 34663
rect 22419 34660 22431 34663
rect 23216 34660 23244 34700
rect 23566 34688 23572 34700
rect 23624 34728 23630 34740
rect 23842 34728 23848 34740
rect 23624 34700 23848 34728
rect 23624 34688 23630 34700
rect 23842 34688 23848 34700
rect 23900 34688 23906 34740
rect 25406 34688 25412 34740
rect 25464 34728 25470 34740
rect 25501 34731 25559 34737
rect 25501 34728 25513 34731
rect 25464 34700 25513 34728
rect 25464 34688 25470 34700
rect 25501 34697 25513 34700
rect 25547 34697 25559 34731
rect 25501 34691 25559 34697
rect 27430 34688 27436 34740
rect 27488 34728 27494 34740
rect 27488 34700 29960 34728
rect 27488 34688 27494 34700
rect 22419 34632 23244 34660
rect 22419 34629 22431 34632
rect 22373 34623 22431 34629
rect 24118 34620 24124 34672
rect 24176 34660 24182 34672
rect 24581 34663 24639 34669
rect 24581 34660 24593 34663
rect 24176 34632 24593 34660
rect 24176 34620 24182 34632
rect 24581 34629 24593 34632
rect 24627 34660 24639 34663
rect 25130 34660 25136 34672
rect 24627 34632 25136 34660
rect 24627 34629 24639 34632
rect 24581 34623 24639 34629
rect 25130 34620 25136 34632
rect 25188 34620 25194 34672
rect 28994 34620 29000 34672
rect 29052 34620 29058 34672
rect 17129 34595 17187 34601
rect 17129 34592 17141 34595
rect 15948 34590 16712 34592
rect 16868 34590 17141 34592
rect 15948 34564 17141 34590
rect 16684 34562 16896 34564
rect 17129 34561 17141 34564
rect 17175 34561 17187 34595
rect 17129 34555 17187 34561
rect 17218 34552 17224 34604
rect 17276 34592 17282 34604
rect 17313 34595 17371 34601
rect 17313 34592 17325 34595
rect 17276 34564 17325 34592
rect 17276 34552 17282 34564
rect 17313 34561 17325 34564
rect 17359 34561 17371 34595
rect 17313 34555 17371 34561
rect 17494 34552 17500 34604
rect 17552 34552 17558 34604
rect 17589 34595 17647 34601
rect 17589 34561 17601 34595
rect 17635 34561 17647 34595
rect 17589 34555 17647 34561
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34561 17831 34595
rect 17773 34555 17831 34561
rect 13538 34524 13544 34536
rect 12032 34496 13544 34524
rect 12032 34484 12038 34496
rect 13538 34484 13544 34496
rect 13596 34524 13602 34536
rect 14366 34524 14372 34536
rect 13596 34496 14372 34524
rect 13596 34484 13602 34496
rect 14366 34484 14372 34496
rect 14424 34524 14430 34536
rect 14918 34524 14924 34536
rect 14424 34496 14924 34524
rect 14424 34484 14430 34496
rect 14918 34484 14924 34496
rect 14976 34484 14982 34536
rect 15381 34527 15439 34533
rect 15381 34493 15393 34527
rect 15427 34493 15439 34527
rect 15381 34487 15439 34493
rect 6549 34459 6607 34465
rect 6549 34425 6561 34459
rect 6595 34456 6607 34459
rect 7926 34456 7932 34468
rect 6595 34428 7932 34456
rect 6595 34425 6607 34428
rect 6549 34419 6607 34425
rect 7926 34416 7932 34428
rect 7984 34416 7990 34468
rect 13998 34416 14004 34468
rect 14056 34456 14062 34468
rect 15010 34456 15016 34468
rect 14056 34428 15016 34456
rect 14056 34416 14062 34428
rect 15010 34416 15016 34428
rect 15068 34416 15074 34468
rect 15396 34456 15424 34487
rect 15562 34484 15568 34536
rect 15620 34484 15626 34536
rect 15654 34484 15660 34536
rect 15712 34484 15718 34536
rect 15746 34484 15752 34536
rect 15804 34524 15810 34536
rect 16025 34527 16083 34533
rect 16025 34524 16037 34527
rect 15804 34496 16037 34524
rect 15804 34484 15810 34496
rect 16025 34493 16037 34496
rect 16071 34524 16083 34527
rect 16482 34524 16488 34536
rect 16071 34496 16488 34524
rect 16071 34493 16083 34496
rect 16025 34487 16083 34493
rect 16482 34484 16488 34496
rect 16540 34524 16546 34536
rect 16853 34527 16911 34533
rect 16853 34524 16865 34527
rect 16540 34496 16865 34524
rect 16540 34484 16546 34496
rect 16853 34493 16865 34496
rect 16899 34493 16911 34527
rect 16853 34487 16911 34493
rect 16945 34527 17003 34533
rect 16945 34493 16957 34527
rect 16991 34493 17003 34527
rect 16945 34487 17003 34493
rect 16206 34456 16212 34468
rect 15396 34428 16212 34456
rect 16206 34416 16212 34428
rect 16264 34416 16270 34468
rect 16298 34416 16304 34468
rect 16356 34416 16362 34468
rect 16390 34416 16396 34468
rect 16448 34456 16454 34468
rect 16960 34456 16988 34487
rect 17034 34484 17040 34536
rect 17092 34524 17098 34536
rect 17604 34524 17632 34555
rect 17092 34496 17632 34524
rect 17788 34524 17816 34555
rect 18046 34552 18052 34604
rect 18104 34552 18110 34604
rect 18414 34552 18420 34604
rect 18472 34552 18478 34604
rect 19150 34552 19156 34604
rect 19208 34552 19214 34604
rect 19426 34592 19432 34604
rect 19306 34564 19432 34592
rect 18874 34524 18880 34536
rect 17788 34496 18880 34524
rect 17092 34484 17098 34496
rect 17788 34456 17816 34496
rect 18874 34484 18880 34496
rect 18932 34484 18938 34536
rect 16448 34428 17816 34456
rect 16448 34416 16454 34428
rect 18598 34416 18604 34468
rect 18656 34456 18662 34468
rect 19306 34456 19334 34564
rect 19426 34552 19432 34564
rect 19484 34552 19490 34604
rect 23934 34552 23940 34604
rect 23992 34592 23998 34604
rect 25038 34592 25044 34604
rect 23992 34564 25044 34592
rect 23992 34552 23998 34564
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 26237 34595 26295 34601
rect 26237 34592 26249 34595
rect 25608 34564 26249 34592
rect 19613 34527 19671 34533
rect 19613 34524 19625 34527
rect 19536 34496 19625 34524
rect 19536 34468 19564 34496
rect 19613 34493 19625 34496
rect 19659 34493 19671 34527
rect 19613 34487 19671 34493
rect 22278 34484 22284 34536
rect 22336 34524 22342 34536
rect 22557 34527 22615 34533
rect 22557 34524 22569 34527
rect 22336 34496 22569 34524
rect 22336 34484 22342 34496
rect 22557 34493 22569 34496
rect 22603 34493 22615 34527
rect 22557 34487 22615 34493
rect 22830 34484 22836 34536
rect 22888 34484 22894 34536
rect 24486 34484 24492 34536
rect 24544 34524 24550 34536
rect 25608 34524 25636 34564
rect 26237 34561 26249 34564
rect 26283 34561 26295 34595
rect 26237 34555 26295 34561
rect 26418 34552 26424 34604
rect 26476 34552 26482 34604
rect 27338 34552 27344 34604
rect 27396 34592 27402 34604
rect 27433 34595 27491 34601
rect 27433 34592 27445 34595
rect 27396 34564 27445 34592
rect 27396 34552 27402 34564
rect 27433 34561 27445 34564
rect 27479 34561 27491 34595
rect 27433 34555 27491 34561
rect 24544 34496 25636 34524
rect 24544 34484 24550 34496
rect 26142 34484 26148 34536
rect 26200 34484 26206 34536
rect 27982 34484 27988 34536
rect 28040 34484 28046 34536
rect 29932 34533 29960 34700
rect 29917 34527 29975 34533
rect 29917 34493 29929 34527
rect 29963 34524 29975 34527
rect 31662 34524 31668 34536
rect 29963 34496 31668 34524
rect 29963 34493 29975 34496
rect 29917 34487 29975 34493
rect 31662 34484 31668 34496
rect 31720 34484 31726 34536
rect 18656 34428 19334 34456
rect 18656 34416 18662 34428
rect 19518 34416 19524 34468
rect 19576 34416 19582 34468
rect 22066 34428 22232 34456
rect 7190 34348 7196 34400
rect 7248 34388 7254 34400
rect 7745 34391 7803 34397
rect 7745 34388 7757 34391
rect 7248 34360 7757 34388
rect 7248 34348 7254 34360
rect 7745 34357 7757 34360
rect 7791 34357 7803 34391
rect 7745 34351 7803 34357
rect 13078 34348 13084 34400
rect 13136 34348 13142 34400
rect 13630 34348 13636 34400
rect 13688 34388 13694 34400
rect 14642 34388 14648 34400
rect 13688 34360 14648 34388
rect 13688 34348 13694 34360
rect 14642 34348 14648 34360
rect 14700 34348 14706 34400
rect 16316 34388 16344 34416
rect 16482 34388 16488 34400
rect 16316 34360 16488 34388
rect 16482 34348 16488 34360
rect 16540 34348 16546 34400
rect 18966 34348 18972 34400
rect 19024 34388 19030 34400
rect 19153 34391 19211 34397
rect 19153 34388 19165 34391
rect 19024 34360 19165 34388
rect 19024 34348 19030 34360
rect 19153 34357 19165 34360
rect 19199 34357 19211 34391
rect 19153 34351 19211 34357
rect 19242 34348 19248 34400
rect 19300 34388 19306 34400
rect 22066 34388 22094 34428
rect 19300 34360 22094 34388
rect 22204 34388 22232 34428
rect 23842 34416 23848 34468
rect 23900 34456 23906 34468
rect 27614 34456 27620 34468
rect 23900 34428 27620 34456
rect 23900 34416 23906 34428
rect 27614 34416 27620 34428
rect 27672 34416 27678 34468
rect 24854 34388 24860 34400
rect 22204 34360 24860 34388
rect 19300 34348 19306 34360
rect 24854 34348 24860 34360
rect 24912 34348 24918 34400
rect 28166 34348 28172 34400
rect 28224 34348 28230 34400
rect 28258 34348 28264 34400
rect 28316 34388 28322 34400
rect 29653 34391 29711 34397
rect 29653 34388 29665 34391
rect 28316 34360 29665 34388
rect 28316 34348 28322 34360
rect 29653 34357 29665 34360
rect 29699 34357 29711 34391
rect 29653 34351 29711 34357
rect 1104 34298 36432 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 36432 34298
rect 1104 34224 36432 34246
rect 5534 34144 5540 34196
rect 5592 34184 5598 34196
rect 5994 34184 6000 34196
rect 5592 34156 6000 34184
rect 5592 34144 5598 34156
rect 5994 34144 6000 34156
rect 6052 34184 6058 34196
rect 6362 34184 6368 34196
rect 6052 34156 6368 34184
rect 6052 34144 6058 34156
rect 6362 34144 6368 34156
rect 6420 34144 6426 34196
rect 7834 34144 7840 34196
rect 7892 34144 7898 34196
rect 9490 34144 9496 34196
rect 9548 34184 9554 34196
rect 9548 34156 9812 34184
rect 9548 34144 9554 34156
rect 6086 34076 6092 34128
rect 6144 34116 6150 34128
rect 7006 34116 7012 34128
rect 6144 34088 7012 34116
rect 6144 34076 6150 34088
rect 7006 34076 7012 34088
rect 7064 34076 7070 34128
rect 7098 34076 7104 34128
rect 7156 34116 7162 34128
rect 7156 34088 8340 34116
rect 7156 34076 7162 34088
rect 5350 34008 5356 34060
rect 5408 34048 5414 34060
rect 6457 34051 6515 34057
rect 6457 34048 6469 34051
rect 5408 34020 6469 34048
rect 5408 34008 5414 34020
rect 6457 34017 6469 34020
rect 6503 34048 6515 34051
rect 7466 34048 7472 34060
rect 6503 34020 7472 34048
rect 6503 34017 6515 34020
rect 6457 34011 6515 34017
rect 7466 34008 7472 34020
rect 7524 34048 7530 34060
rect 8202 34048 8208 34060
rect 7524 34020 8208 34048
rect 7524 34008 7530 34020
rect 8202 34008 8208 34020
rect 8260 34008 8266 34060
rect 8312 34057 8340 34088
rect 8386 34076 8392 34128
rect 8444 34076 8450 34128
rect 8938 34076 8944 34128
rect 8996 34116 9002 34128
rect 9122 34116 9128 34128
rect 8996 34088 9128 34116
rect 8996 34076 9002 34088
rect 9122 34076 9128 34088
rect 9180 34116 9186 34128
rect 9784 34116 9812 34156
rect 9858 34144 9864 34196
rect 9916 34144 9922 34196
rect 11514 34144 11520 34196
rect 11572 34184 11578 34196
rect 11793 34187 11851 34193
rect 11793 34184 11805 34187
rect 11572 34156 11805 34184
rect 11572 34144 11578 34156
rect 11793 34153 11805 34156
rect 11839 34153 11851 34187
rect 11793 34147 11851 34153
rect 12434 34144 12440 34196
rect 12492 34184 12498 34196
rect 12897 34187 12955 34193
rect 12897 34184 12909 34187
rect 12492 34156 12909 34184
rect 12492 34144 12498 34156
rect 12897 34153 12909 34156
rect 12943 34153 12955 34187
rect 12897 34147 12955 34153
rect 10137 34119 10195 34125
rect 10137 34116 10149 34119
rect 9180 34088 9674 34116
rect 9784 34088 10149 34116
rect 9180 34076 9186 34088
rect 8297 34051 8355 34057
rect 8297 34017 8309 34051
rect 8343 34048 8355 34051
rect 8478 34048 8484 34060
rect 8343 34020 8484 34048
rect 8343 34017 8355 34020
rect 8297 34011 8355 34017
rect 8478 34008 8484 34020
rect 8536 34048 8542 34060
rect 9398 34048 9404 34060
rect 8536 34020 9404 34048
rect 8536 34008 8542 34020
rect 9398 34008 9404 34020
rect 9456 34008 9462 34060
rect 9490 34008 9496 34060
rect 9548 34008 9554 34060
rect 9646 34048 9674 34088
rect 10137 34085 10149 34088
rect 10183 34085 10195 34119
rect 12158 34116 12164 34128
rect 10137 34079 10195 34085
rect 11072 34088 12164 34116
rect 9646 34020 9812 34048
rect 4706 33940 4712 33992
rect 4764 33940 4770 33992
rect 6270 33940 6276 33992
rect 6328 33980 6334 33992
rect 6641 33983 6699 33989
rect 6641 33980 6653 33983
rect 6328 33952 6653 33980
rect 6328 33940 6334 33952
rect 6641 33949 6653 33952
rect 6687 33949 6699 33983
rect 6641 33943 6699 33949
rect 6822 33940 6828 33992
rect 6880 33940 6886 33992
rect 6914 33940 6920 33992
rect 6972 33940 6978 33992
rect 7190 33940 7196 33992
rect 7248 33940 7254 33992
rect 7282 33940 7288 33992
rect 7340 33980 7346 33992
rect 7653 33983 7711 33989
rect 7653 33980 7665 33983
rect 7340 33952 7665 33980
rect 7340 33940 7346 33952
rect 7653 33949 7665 33952
rect 7699 33949 7711 33983
rect 7653 33943 7711 33949
rect 7742 33940 7748 33992
rect 7800 33980 7806 33992
rect 8021 33983 8079 33989
rect 8021 33980 8033 33983
rect 7800 33952 8033 33980
rect 7800 33940 7806 33952
rect 8021 33949 8033 33952
rect 8067 33949 8079 33983
rect 8021 33943 8079 33949
rect 4985 33915 5043 33921
rect 4985 33881 4997 33915
rect 5031 33912 5043 33915
rect 5258 33912 5264 33924
rect 5031 33884 5264 33912
rect 5031 33881 5043 33884
rect 4985 33875 5043 33881
rect 5258 33872 5264 33884
rect 5316 33872 5322 33924
rect 6210 33884 6316 33912
rect 4614 33804 4620 33856
rect 4672 33844 4678 33856
rect 6288 33844 6316 33884
rect 6546 33844 6552 33856
rect 4672 33816 6552 33844
rect 4672 33804 4678 33816
rect 6546 33804 6552 33816
rect 6604 33804 6610 33856
rect 6638 33804 6644 33856
rect 6696 33804 6702 33856
rect 7098 33804 7104 33856
rect 7156 33844 7162 33856
rect 7374 33844 7380 33856
rect 7156 33816 7380 33844
rect 7156 33804 7162 33816
rect 7374 33804 7380 33816
rect 7432 33804 7438 33856
rect 8036 33844 8064 33943
rect 8110 33940 8116 33992
rect 8168 33980 8174 33992
rect 8665 33983 8723 33989
rect 8665 33980 8677 33983
rect 8168 33952 8677 33980
rect 8168 33940 8174 33952
rect 8665 33949 8677 33952
rect 8711 33949 8723 33983
rect 9610 33983 9668 33989
rect 9610 33980 9622 33983
rect 8665 33943 8723 33949
rect 9600 33949 9622 33980
rect 9656 33949 9668 33983
rect 9784 33980 9812 34020
rect 9950 34008 9956 34060
rect 10008 34048 10014 34060
rect 10045 34051 10103 34057
rect 10045 34048 10057 34051
rect 10008 34020 10057 34048
rect 10008 34008 10014 34020
rect 10045 34017 10057 34020
rect 10091 34017 10103 34051
rect 10045 34011 10103 34017
rect 10152 34020 10364 34048
rect 10152 33980 10180 34020
rect 9784 33952 10180 33980
rect 9600 33943 9668 33949
rect 8297 33915 8355 33921
rect 8297 33881 8309 33915
rect 8343 33912 8355 33915
rect 8389 33915 8447 33921
rect 8389 33912 8401 33915
rect 8343 33884 8401 33912
rect 8343 33881 8355 33884
rect 8297 33875 8355 33881
rect 8389 33881 8401 33884
rect 8435 33881 8447 33915
rect 9600 33912 9628 33943
rect 10226 33940 10232 33992
rect 10284 33940 10290 33992
rect 10336 33989 10364 34020
rect 10686 34008 10692 34060
rect 10744 34048 10750 34060
rect 11072 34048 11100 34088
rect 12158 34076 12164 34088
rect 12216 34076 12222 34128
rect 12912 34116 12940 34147
rect 13814 34144 13820 34196
rect 13872 34144 13878 34196
rect 14090 34144 14096 34196
rect 14148 34144 14154 34196
rect 15289 34187 15347 34193
rect 15289 34184 15301 34187
rect 14200 34156 15301 34184
rect 12912 34088 13676 34116
rect 10744 34020 11100 34048
rect 10744 34008 10750 34020
rect 10980 33989 11008 34020
rect 11422 34008 11428 34060
rect 11480 34008 11486 34060
rect 12342 34048 12348 34060
rect 11532 34020 12348 34048
rect 11532 33989 11560 34020
rect 12342 34008 12348 34020
rect 12400 34048 12406 34060
rect 12400 34020 12480 34048
rect 12400 34008 12406 34020
rect 10321 33983 10379 33989
rect 10321 33949 10333 33983
rect 10367 33949 10379 33983
rect 10321 33943 10379 33949
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33949 10839 33983
rect 10781 33943 10839 33949
rect 10873 33983 10931 33989
rect 10873 33949 10885 33983
rect 10919 33949 10931 33983
rect 10873 33943 10931 33949
rect 10965 33983 11023 33989
rect 10965 33949 10977 33983
rect 11011 33949 11023 33983
rect 11517 33983 11575 33989
rect 11517 33980 11529 33983
rect 10965 33943 11023 33949
rect 11072 33952 11529 33980
rect 10244 33912 10272 33940
rect 10796 33912 10824 33943
rect 9600 33884 9720 33912
rect 10244 33884 10824 33912
rect 8389 33875 8447 33881
rect 8573 33847 8631 33853
rect 8573 33844 8585 33847
rect 8036 33816 8585 33844
rect 8573 33813 8585 33816
rect 8619 33844 8631 33847
rect 9490 33844 9496 33856
rect 8619 33816 9496 33844
rect 8619 33813 8631 33816
rect 8573 33807 8631 33813
rect 9490 33804 9496 33816
rect 9548 33804 9554 33856
rect 9692 33844 9720 33884
rect 10410 33844 10416 33856
rect 9692 33816 10416 33844
rect 10410 33804 10416 33816
rect 10468 33844 10474 33856
rect 10888 33844 10916 33943
rect 11072 33924 11100 33952
rect 11517 33949 11529 33952
rect 11563 33949 11575 33983
rect 11517 33943 11575 33949
rect 12250 33940 12256 33992
rect 12308 33940 12314 33992
rect 12452 33989 12480 34020
rect 13078 34008 13084 34060
rect 13136 34008 13142 34060
rect 12437 33983 12495 33989
rect 12437 33949 12449 33983
rect 12483 33949 12495 33983
rect 12437 33943 12495 33949
rect 12710 33940 12716 33992
rect 12768 33940 12774 33992
rect 12986 33940 12992 33992
rect 13044 33980 13050 33992
rect 13648 33989 13676 34088
rect 13909 34051 13967 34057
rect 13909 34017 13921 34051
rect 13955 34048 13967 34051
rect 13998 34048 14004 34060
rect 13955 34020 14004 34048
rect 13955 34017 13967 34020
rect 13909 34011 13967 34017
rect 13998 34008 14004 34020
rect 14056 34008 14062 34060
rect 13173 33983 13231 33989
rect 13173 33980 13185 33983
rect 13044 33952 13185 33980
rect 13044 33940 13050 33952
rect 13173 33949 13185 33952
rect 13219 33949 13231 33983
rect 13173 33943 13231 33949
rect 13633 33983 13691 33989
rect 13633 33949 13645 33983
rect 13679 33949 13691 33983
rect 13633 33943 13691 33949
rect 13722 33940 13728 33992
rect 13780 33940 13786 33992
rect 11054 33872 11060 33924
rect 11112 33872 11118 33924
rect 14200 33912 14228 34156
rect 15289 34153 15301 34156
rect 15335 34153 15347 34187
rect 15289 34147 15347 34153
rect 15654 34144 15660 34196
rect 15712 34184 15718 34196
rect 16114 34184 16120 34196
rect 15712 34156 16120 34184
rect 15712 34144 15718 34156
rect 16114 34144 16120 34156
rect 16172 34184 16178 34196
rect 16209 34187 16267 34193
rect 16209 34184 16221 34187
rect 16172 34156 16221 34184
rect 16172 34144 16178 34156
rect 16209 34153 16221 34156
rect 16255 34153 16267 34187
rect 17310 34184 17316 34196
rect 16209 34147 16267 34153
rect 16684 34156 17316 34184
rect 14274 34076 14280 34128
rect 14332 34076 14338 34128
rect 14461 34119 14519 34125
rect 14461 34085 14473 34119
rect 14507 34116 14519 34119
rect 14550 34116 14556 34128
rect 14507 34088 14556 34116
rect 14507 34085 14519 34088
rect 14461 34079 14519 34085
rect 14550 34076 14556 34088
rect 14608 34076 14614 34128
rect 14642 34076 14648 34128
rect 14700 34076 14706 34128
rect 14734 34076 14740 34128
rect 14792 34116 14798 34128
rect 15197 34119 15255 34125
rect 15197 34116 15209 34119
rect 14792 34088 15209 34116
rect 14792 34076 14798 34088
rect 15197 34085 15209 34088
rect 15243 34116 15255 34119
rect 15243 34088 15884 34116
rect 15243 34085 15255 34088
rect 15197 34079 15255 34085
rect 14292 34048 14320 34076
rect 14292 34020 14872 34048
rect 14366 33940 14372 33992
rect 14424 33940 14430 33992
rect 14844 33989 14872 34020
rect 14918 34008 14924 34060
rect 14976 34048 14982 34060
rect 15856 34057 15884 34088
rect 16684 34060 16712 34156
rect 17310 34144 17316 34156
rect 17368 34144 17374 34196
rect 17420 34156 22094 34184
rect 16853 34119 16911 34125
rect 16853 34085 16865 34119
rect 16899 34085 16911 34119
rect 16853 34079 16911 34085
rect 15105 34051 15163 34057
rect 15105 34048 15117 34051
rect 14976 34020 15117 34048
rect 14976 34008 14982 34020
rect 15105 34017 15117 34020
rect 15151 34017 15163 34051
rect 15105 34011 15163 34017
rect 15841 34051 15899 34057
rect 15841 34017 15853 34051
rect 15887 34017 15899 34051
rect 16577 34051 16635 34057
rect 16577 34048 16589 34051
rect 15841 34011 15899 34017
rect 15948 34020 16589 34048
rect 14553 33983 14611 33989
rect 14553 33949 14565 33983
rect 14599 33949 14611 33983
rect 14553 33943 14611 33949
rect 14829 33983 14887 33989
rect 14829 33949 14841 33983
rect 14875 33949 14887 33983
rect 14829 33943 14887 33949
rect 14568 33912 14596 33943
rect 15194 33940 15200 33992
rect 15252 33940 15258 33992
rect 15286 33940 15292 33992
rect 15344 33940 15350 33992
rect 15473 33983 15531 33989
rect 15473 33949 15485 33983
rect 15519 33949 15531 33983
rect 15473 33943 15531 33949
rect 15565 33983 15623 33989
rect 15565 33949 15577 33983
rect 15611 33980 15623 33983
rect 15948 33980 15976 34020
rect 16577 34017 16589 34020
rect 16623 34048 16635 34051
rect 16666 34048 16672 34060
rect 16623 34020 16672 34048
rect 16623 34017 16635 34020
rect 16577 34011 16635 34017
rect 16666 34008 16672 34020
rect 16724 34008 16730 34060
rect 16868 34048 16896 34079
rect 17037 34051 17095 34057
rect 17037 34048 17049 34051
rect 16868 34020 17049 34048
rect 17037 34017 17049 34020
rect 17083 34017 17095 34051
rect 17037 34011 17095 34017
rect 15611 33952 15976 33980
rect 16025 33983 16083 33989
rect 15611 33949 15623 33952
rect 15565 33943 15623 33949
rect 16025 33949 16037 33983
rect 16071 33949 16083 33983
rect 16485 33983 16543 33989
rect 16485 33980 16497 33983
rect 16025 33943 16083 33949
rect 16224 33952 16497 33980
rect 11256 33884 14228 33912
rect 14384 33884 14596 33912
rect 11256 33853 11284 33884
rect 10468 33816 10916 33844
rect 11241 33847 11299 33853
rect 10468 33804 10474 33816
rect 11241 33813 11253 33847
rect 11287 33813 11299 33847
rect 11241 33807 11299 33813
rect 13541 33847 13599 33853
rect 13541 33813 13553 33847
rect 13587 33844 13599 33847
rect 13814 33844 13820 33856
rect 13587 33816 13820 33844
rect 13587 33813 13599 33816
rect 13541 33807 13599 33813
rect 13814 33804 13820 33816
rect 13872 33804 13878 33856
rect 13906 33804 13912 33856
rect 13964 33844 13970 33856
rect 14384 33844 14412 33884
rect 14918 33872 14924 33924
rect 14976 33872 14982 33924
rect 15488 33912 15516 33943
rect 15838 33912 15844 33924
rect 15488 33884 15844 33912
rect 13964 33816 14412 33844
rect 13964 33804 13970 33816
rect 14642 33804 14648 33856
rect 14700 33844 14706 33856
rect 15488 33844 15516 33884
rect 15838 33872 15844 33884
rect 15896 33912 15902 33924
rect 16040 33912 16068 33943
rect 15896 33884 16068 33912
rect 15896 33872 15902 33884
rect 14700 33816 15516 33844
rect 14700 33804 14706 33816
rect 15746 33804 15752 33856
rect 15804 33804 15810 33856
rect 16022 33804 16028 33856
rect 16080 33844 16086 33856
rect 16224 33844 16252 33952
rect 16485 33949 16497 33952
rect 16531 33949 16543 33983
rect 16485 33943 16543 33949
rect 17126 33940 17132 33992
rect 17184 33940 17190 33992
rect 16298 33872 16304 33924
rect 16356 33912 16362 33924
rect 17420 33912 17448 34156
rect 17497 34119 17555 34125
rect 17497 34085 17509 34119
rect 17543 34085 17555 34119
rect 18785 34119 18843 34125
rect 18785 34116 18797 34119
rect 17497 34079 17555 34085
rect 17972 34088 18797 34116
rect 16356 33884 17448 33912
rect 17512 33912 17540 34079
rect 17865 33983 17923 33989
rect 17865 33949 17877 33983
rect 17911 33980 17923 33983
rect 17972 33980 18000 34088
rect 18785 34085 18797 34088
rect 18831 34085 18843 34119
rect 18785 34079 18843 34085
rect 18322 34008 18328 34060
rect 18380 34048 18386 34060
rect 18693 34051 18751 34057
rect 18693 34048 18705 34051
rect 18380 34020 18705 34048
rect 18380 34008 18386 34020
rect 18693 34017 18705 34020
rect 18739 34017 18751 34051
rect 18693 34011 18751 34017
rect 19245 34051 19303 34057
rect 19245 34017 19257 34051
rect 19291 34048 19303 34051
rect 19518 34048 19524 34060
rect 19291 34020 19524 34048
rect 19291 34017 19303 34020
rect 19245 34011 19303 34017
rect 19518 34008 19524 34020
rect 19576 34008 19582 34060
rect 22066 34048 22094 34156
rect 22830 34144 22836 34196
rect 22888 34184 22894 34196
rect 23109 34187 23167 34193
rect 23109 34184 23121 34187
rect 22888 34156 23121 34184
rect 22888 34144 22894 34156
rect 23109 34153 23121 34156
rect 23155 34153 23167 34187
rect 23109 34147 23167 34153
rect 24762 34144 24768 34196
rect 24820 34184 24826 34196
rect 29362 34184 29368 34196
rect 24820 34156 25544 34184
rect 24820 34144 24826 34156
rect 22646 34076 22652 34128
rect 22704 34116 22710 34128
rect 25516 34116 25544 34156
rect 26344 34156 29368 34184
rect 26344 34116 26372 34156
rect 29362 34144 29368 34156
rect 29420 34144 29426 34196
rect 22704 34088 24348 34116
rect 25516 34088 26372 34116
rect 22704 34076 22710 34088
rect 22066 34020 23520 34048
rect 17911 33952 18000 33980
rect 18049 33983 18107 33989
rect 17911 33949 17923 33952
rect 17865 33943 17923 33949
rect 18049 33949 18061 33983
rect 18095 33949 18107 33983
rect 18049 33943 18107 33949
rect 18064 33912 18092 33943
rect 18138 33940 18144 33992
rect 18196 33940 18202 33992
rect 18230 33940 18236 33992
rect 18288 33940 18294 33992
rect 18417 33983 18475 33989
rect 18417 33949 18429 33983
rect 18463 33949 18475 33983
rect 18417 33943 18475 33949
rect 17512 33884 18092 33912
rect 16356 33872 16362 33884
rect 18432 33844 18460 33943
rect 18506 33940 18512 33992
rect 18564 33980 18570 33992
rect 18877 33983 18935 33989
rect 18877 33980 18889 33983
rect 18564 33952 18889 33980
rect 18564 33940 18570 33952
rect 18877 33949 18889 33952
rect 18923 33949 18935 33983
rect 18877 33943 18935 33949
rect 18966 33940 18972 33992
rect 19024 33940 19030 33992
rect 21634 33940 21640 33992
rect 21692 33940 21698 33992
rect 22002 33940 22008 33992
rect 22060 33940 22066 33992
rect 22278 33940 22284 33992
rect 22336 33980 22342 33992
rect 22373 33983 22431 33989
rect 22373 33980 22385 33983
rect 22336 33952 22385 33980
rect 22336 33940 22342 33952
rect 22373 33949 22385 33952
rect 22419 33980 22431 33983
rect 23198 33980 23204 33992
rect 22419 33952 23204 33980
rect 22419 33949 22431 33952
rect 22373 33943 22431 33949
rect 23198 33940 23204 33952
rect 23256 33940 23262 33992
rect 23492 33989 23520 34020
rect 23658 34008 23664 34060
rect 23716 34008 23722 34060
rect 23477 33983 23535 33989
rect 23477 33949 23489 33983
rect 23523 33949 23535 33983
rect 23477 33943 23535 33949
rect 23569 33983 23627 33989
rect 23569 33949 23581 33983
rect 23615 33980 23627 33983
rect 24118 33980 24124 33992
rect 23615 33952 24124 33980
rect 23615 33949 23627 33952
rect 23569 33943 23627 33949
rect 24118 33940 24124 33952
rect 24176 33940 24182 33992
rect 24213 33983 24271 33989
rect 24213 33949 24225 33983
rect 24259 33949 24271 33983
rect 24213 33943 24271 33949
rect 18601 33915 18659 33921
rect 18601 33881 18613 33915
rect 18647 33912 18659 33915
rect 19521 33915 19579 33921
rect 19521 33912 19533 33915
rect 18647 33884 19533 33912
rect 18647 33881 18659 33884
rect 18601 33875 18659 33881
rect 19521 33881 19533 33884
rect 19567 33881 19579 33915
rect 19521 33875 19579 33881
rect 20254 33872 20260 33924
rect 20312 33872 20318 33924
rect 21821 33915 21879 33921
rect 21821 33881 21833 33915
rect 21867 33881 21879 33915
rect 21821 33875 21879 33881
rect 21913 33915 21971 33921
rect 21913 33881 21925 33915
rect 21959 33912 21971 33915
rect 21959 33884 23520 33912
rect 21959 33881 21971 33884
rect 21913 33875 21971 33881
rect 20993 33847 21051 33853
rect 20993 33844 21005 33847
rect 16080 33816 21005 33844
rect 16080 33804 16086 33816
rect 20993 33813 21005 33816
rect 21039 33813 21051 33847
rect 21836 33844 21864 33875
rect 23492 33856 23520 33884
rect 23934 33872 23940 33924
rect 23992 33912 23998 33924
rect 24228 33912 24256 33943
rect 23992 33884 24256 33912
rect 23992 33872 23998 33884
rect 22002 33844 22008 33856
rect 21836 33816 22008 33844
rect 20993 33807 21051 33813
rect 22002 33804 22008 33816
rect 22060 33804 22066 33856
rect 22189 33847 22247 33853
rect 22189 33813 22201 33847
rect 22235 33844 22247 33847
rect 22370 33844 22376 33856
rect 22235 33816 22376 33844
rect 22235 33813 22247 33816
rect 22189 33807 22247 33813
rect 22370 33804 22376 33816
rect 22428 33804 22434 33856
rect 23474 33804 23480 33856
rect 23532 33804 23538 33856
rect 24026 33804 24032 33856
rect 24084 33804 24090 33856
rect 24320 33844 24348 34088
rect 27614 34076 27620 34128
rect 27672 34116 27678 34128
rect 29454 34116 29460 34128
rect 27672 34088 29460 34116
rect 27672 34076 27678 34088
rect 29454 34076 29460 34088
rect 29512 34076 29518 34128
rect 24397 34051 24455 34057
rect 24397 34017 24409 34051
rect 24443 34048 24455 34051
rect 25314 34048 25320 34060
rect 24443 34020 25320 34048
rect 24443 34017 24455 34020
rect 24397 34011 24455 34017
rect 25314 34008 25320 34020
rect 25372 34048 25378 34060
rect 25498 34048 25504 34060
rect 25372 34020 25504 34048
rect 25372 34008 25378 34020
rect 25498 34008 25504 34020
rect 25556 34048 25562 34060
rect 26329 34051 26387 34057
rect 26329 34048 26341 34051
rect 25556 34020 26341 34048
rect 25556 34008 25562 34020
rect 26329 34017 26341 34020
rect 26375 34048 26387 34051
rect 27338 34048 27344 34060
rect 26375 34020 27344 34048
rect 26375 34017 26387 34020
rect 26329 34011 26387 34017
rect 27338 34008 27344 34020
rect 27396 34008 27402 34060
rect 28166 34008 28172 34060
rect 28224 34048 28230 34060
rect 28353 34051 28411 34057
rect 28353 34048 28365 34051
rect 28224 34020 28365 34048
rect 28224 34008 28230 34020
rect 28353 34017 28365 34020
rect 28399 34017 28411 34051
rect 28353 34011 28411 34017
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33980 24823 33983
rect 24854 33980 24860 33992
rect 24811 33952 24860 33980
rect 24811 33949 24823 33952
rect 24765 33943 24823 33949
rect 24854 33940 24860 33952
rect 24912 33940 24918 33992
rect 27908 33952 29224 33980
rect 25774 33872 25780 33924
rect 25832 33872 25838 33924
rect 26142 33872 26148 33924
rect 26200 33921 26206 33924
rect 26200 33915 26249 33921
rect 26200 33881 26203 33915
rect 26237 33881 26249 33915
rect 26200 33875 26249 33881
rect 26200 33872 26206 33875
rect 26602 33872 26608 33924
rect 26660 33872 26666 33924
rect 26878 33872 26884 33924
rect 26936 33912 26942 33924
rect 26936 33884 27094 33912
rect 26936 33872 26942 33884
rect 27908 33844 27936 33952
rect 29196 33924 29224 33952
rect 30190 33940 30196 33992
rect 30248 33980 30254 33992
rect 30377 33983 30435 33989
rect 30377 33980 30389 33983
rect 30248 33952 30389 33980
rect 30248 33940 30254 33952
rect 30377 33949 30389 33952
rect 30423 33949 30435 33983
rect 30377 33943 30435 33949
rect 32490 33940 32496 33992
rect 32548 33980 32554 33992
rect 32769 33983 32827 33989
rect 32769 33980 32781 33983
rect 32548 33952 32781 33980
rect 32548 33940 32554 33952
rect 32769 33949 32781 33952
rect 32815 33949 32827 33983
rect 32769 33943 32827 33949
rect 28902 33872 28908 33924
rect 28960 33912 28966 33924
rect 28960 33884 29132 33912
rect 28960 33872 28966 33884
rect 24320 33816 27936 33844
rect 27982 33804 27988 33856
rect 28040 33844 28046 33856
rect 28077 33847 28135 33853
rect 28077 33844 28089 33847
rect 28040 33816 28089 33844
rect 28040 33804 28046 33816
rect 28077 33813 28089 33816
rect 28123 33813 28135 33847
rect 28077 33807 28135 33813
rect 28534 33804 28540 33856
rect 28592 33844 28598 33856
rect 28997 33847 29055 33853
rect 28997 33844 29009 33847
rect 28592 33816 29009 33844
rect 28592 33804 28598 33816
rect 28997 33813 29009 33816
rect 29043 33813 29055 33847
rect 29104 33844 29132 33884
rect 29178 33872 29184 33924
rect 29236 33912 29242 33924
rect 29641 33915 29699 33921
rect 29641 33912 29653 33915
rect 29236 33884 29653 33912
rect 29236 33872 29242 33884
rect 29641 33881 29653 33884
rect 29687 33881 29699 33915
rect 29641 33875 29699 33881
rect 29914 33872 29920 33924
rect 29972 33912 29978 33924
rect 29972 33884 31754 33912
rect 29972 33872 29978 33884
rect 29733 33847 29791 33853
rect 29733 33844 29745 33847
rect 29104 33816 29745 33844
rect 28997 33807 29055 33813
rect 29733 33813 29745 33816
rect 29779 33813 29791 33847
rect 29733 33807 29791 33813
rect 30193 33847 30251 33853
rect 30193 33813 30205 33847
rect 30239 33844 30251 33847
rect 31570 33844 31576 33856
rect 30239 33816 31576 33844
rect 30239 33813 30251 33816
rect 30193 33807 30251 33813
rect 31570 33804 31576 33816
rect 31628 33804 31634 33856
rect 31726 33844 31754 33884
rect 32585 33847 32643 33853
rect 32585 33844 32597 33847
rect 31726 33816 32597 33844
rect 32585 33813 32597 33816
rect 32631 33844 32643 33847
rect 32858 33844 32864 33856
rect 32631 33816 32864 33844
rect 32631 33813 32643 33816
rect 32585 33807 32643 33813
rect 32858 33804 32864 33816
rect 32916 33804 32922 33856
rect 1104 33754 36432 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 36432 33754
rect 1104 33680 36432 33702
rect 5077 33643 5135 33649
rect 5077 33609 5089 33643
rect 5123 33640 5135 33643
rect 5258 33640 5264 33652
rect 5123 33612 5264 33640
rect 5123 33609 5135 33612
rect 5077 33603 5135 33609
rect 5258 33600 5264 33612
rect 5316 33600 5322 33652
rect 6178 33600 6184 33652
rect 6236 33640 6242 33652
rect 6365 33643 6423 33649
rect 6365 33640 6377 33643
rect 6236 33612 6377 33640
rect 6236 33600 6242 33612
rect 6365 33609 6377 33612
rect 6411 33609 6423 33643
rect 7190 33640 7196 33652
rect 6365 33603 6423 33609
rect 6564 33612 7196 33640
rect 5534 33572 5540 33584
rect 5460 33544 5540 33572
rect 5261 33507 5319 33513
rect 5261 33473 5273 33507
rect 5307 33504 5319 33507
rect 5350 33504 5356 33516
rect 5307 33476 5356 33504
rect 5307 33473 5319 33476
rect 5261 33467 5319 33473
rect 5350 33464 5356 33476
rect 5408 33464 5414 33516
rect 5460 33513 5488 33544
rect 5534 33532 5540 33544
rect 5592 33532 5598 33584
rect 5905 33575 5963 33581
rect 5905 33541 5917 33575
rect 5951 33572 5963 33575
rect 6564 33572 6592 33612
rect 7190 33600 7196 33612
rect 7248 33600 7254 33652
rect 7745 33643 7803 33649
rect 7745 33609 7757 33643
rect 7791 33640 7803 33643
rect 8110 33640 8116 33652
rect 7791 33612 8116 33640
rect 7791 33609 7803 33612
rect 7745 33603 7803 33609
rect 8110 33600 8116 33612
rect 8168 33600 8174 33652
rect 8294 33600 8300 33652
rect 8352 33600 8358 33652
rect 9398 33600 9404 33652
rect 9456 33640 9462 33652
rect 10686 33640 10692 33652
rect 9456 33612 10692 33640
rect 9456 33600 9462 33612
rect 10686 33600 10692 33612
rect 10744 33600 10750 33652
rect 11422 33600 11428 33652
rect 11480 33640 11486 33652
rect 11517 33643 11575 33649
rect 11517 33640 11529 33643
rect 11480 33612 11529 33640
rect 11480 33600 11486 33612
rect 11517 33609 11529 33612
rect 11563 33609 11575 33643
rect 11517 33603 11575 33609
rect 12250 33600 12256 33652
rect 12308 33640 12314 33652
rect 14918 33640 14924 33652
rect 12308 33612 14924 33640
rect 12308 33600 12314 33612
rect 14918 33600 14924 33612
rect 14976 33600 14982 33652
rect 15378 33600 15384 33652
rect 15436 33640 15442 33652
rect 16117 33643 16175 33649
rect 15436 33612 15700 33640
rect 15436 33600 15442 33612
rect 5951 33544 6592 33572
rect 5951 33541 5963 33544
rect 5905 33535 5963 33541
rect 6638 33532 6644 33584
rect 6696 33532 6702 33584
rect 8312 33572 8340 33600
rect 9582 33572 9588 33584
rect 6932 33544 7696 33572
rect 5445 33507 5503 33513
rect 5445 33473 5457 33507
rect 5491 33473 5503 33507
rect 5445 33467 5503 33473
rect 5629 33507 5687 33513
rect 5629 33473 5641 33507
rect 5675 33473 5687 33507
rect 5629 33467 5687 33473
rect 5813 33507 5871 33513
rect 5813 33473 5825 33507
rect 5859 33504 5871 33507
rect 5859 33476 6132 33504
rect 5859 33473 5871 33476
rect 5813 33467 5871 33473
rect 5534 33396 5540 33448
rect 5592 33396 5598 33448
rect 5258 33328 5264 33380
rect 5316 33368 5322 33380
rect 5644 33368 5672 33467
rect 6104 33436 6132 33476
rect 6178 33464 6184 33516
rect 6236 33464 6242 33516
rect 6549 33507 6607 33513
rect 6549 33473 6561 33507
rect 6595 33473 6607 33507
rect 6549 33467 6607 33473
rect 6104 33408 6408 33436
rect 5316 33340 5672 33368
rect 6089 33371 6147 33377
rect 5316 33328 5322 33340
rect 6089 33337 6101 33371
rect 6135 33368 6147 33371
rect 6380 33368 6408 33408
rect 6454 33396 6460 33448
rect 6512 33436 6518 33448
rect 6564 33436 6592 33467
rect 6730 33464 6736 33516
rect 6788 33464 6794 33516
rect 6932 33513 6960 33544
rect 6917 33507 6975 33513
rect 6917 33473 6929 33507
rect 6963 33473 6975 33507
rect 6917 33467 6975 33473
rect 7101 33507 7159 33513
rect 7101 33473 7113 33507
rect 7147 33504 7159 33507
rect 7190 33504 7196 33516
rect 7147 33476 7196 33504
rect 7147 33473 7159 33476
rect 7101 33467 7159 33473
rect 7190 33464 7196 33476
rect 7248 33464 7254 33516
rect 7285 33507 7343 33513
rect 7285 33473 7297 33507
rect 7331 33504 7343 33507
rect 7374 33504 7380 33516
rect 7331 33476 7380 33504
rect 7331 33473 7343 33476
rect 7285 33467 7343 33473
rect 7374 33464 7380 33476
rect 7432 33464 7438 33516
rect 7561 33507 7619 33513
rect 7561 33473 7573 33507
rect 7607 33473 7619 33507
rect 7561 33467 7619 33473
rect 7576 33436 7604 33467
rect 6512 33408 7604 33436
rect 6512 33396 6518 33408
rect 7282 33368 7288 33380
rect 6135 33340 6316 33368
rect 6380 33340 7288 33368
rect 6135 33337 6147 33340
rect 6089 33331 6147 33337
rect 6178 33260 6184 33312
rect 6236 33260 6242 33312
rect 6288 33300 6316 33340
rect 7282 33328 7288 33340
rect 7340 33328 7346 33380
rect 6914 33300 6920 33312
rect 6288 33272 6920 33300
rect 6914 33260 6920 33272
rect 6972 33260 6978 33312
rect 7190 33260 7196 33312
rect 7248 33300 7254 33312
rect 7668 33300 7696 33544
rect 7852 33544 8340 33572
rect 9338 33544 9588 33572
rect 7852 33513 7880 33544
rect 9582 33532 9588 33544
rect 9640 33532 9646 33584
rect 9674 33532 9680 33584
rect 9732 33572 9738 33584
rect 10321 33575 10379 33581
rect 10321 33572 10333 33575
rect 9732 33544 10333 33572
rect 9732 33532 9738 33544
rect 10321 33541 10333 33544
rect 10367 33541 10379 33575
rect 10321 33535 10379 33541
rect 11333 33575 11391 33581
rect 11333 33541 11345 33575
rect 11379 33572 11391 33575
rect 12710 33572 12716 33584
rect 11379 33544 12716 33572
rect 11379 33541 11391 33544
rect 11333 33535 11391 33541
rect 12710 33532 12716 33544
rect 12768 33532 12774 33584
rect 13173 33575 13231 33581
rect 13173 33541 13185 33575
rect 13219 33572 13231 33575
rect 15562 33572 15568 33584
rect 13219 33544 14964 33572
rect 13219 33541 13231 33544
rect 13173 33535 13231 33541
rect 7837 33507 7895 33513
rect 7837 33473 7849 33507
rect 7883 33473 7895 33507
rect 10137 33507 10195 33513
rect 10137 33504 10149 33507
rect 7837 33467 7895 33473
rect 9324 33476 10149 33504
rect 8110 33396 8116 33448
rect 8168 33396 8174 33448
rect 8570 33300 8576 33312
rect 7248 33272 8576 33300
rect 7248 33260 7254 33272
rect 8570 33260 8576 33272
rect 8628 33300 8634 33312
rect 9324 33300 9352 33476
rect 10137 33473 10149 33476
rect 10183 33473 10195 33507
rect 10137 33467 10195 33473
rect 10229 33507 10287 33513
rect 10229 33473 10241 33507
rect 10275 33504 10287 33507
rect 10410 33504 10416 33516
rect 10275 33476 10416 33504
rect 10275 33473 10287 33476
rect 10229 33467 10287 33473
rect 10410 33464 10416 33476
rect 10468 33464 10474 33516
rect 10505 33507 10563 33513
rect 10505 33473 10517 33507
rect 10551 33504 10563 33507
rect 11149 33507 11207 33513
rect 11149 33504 11161 33507
rect 10551 33476 11161 33504
rect 10551 33473 10563 33476
rect 10505 33467 10563 33473
rect 11149 33473 11161 33476
rect 11195 33504 11207 33507
rect 11701 33507 11759 33513
rect 11701 33504 11713 33507
rect 11195 33476 11713 33504
rect 11195 33473 11207 33476
rect 11149 33467 11207 33473
rect 11701 33473 11713 33476
rect 11747 33473 11759 33507
rect 11977 33507 12035 33513
rect 11977 33504 11989 33507
rect 11701 33467 11759 33473
rect 11808 33476 11989 33504
rect 9398 33396 9404 33448
rect 9456 33436 9462 33448
rect 9861 33439 9919 33445
rect 9861 33436 9873 33439
rect 9456 33408 9873 33436
rect 9456 33396 9462 33408
rect 9861 33405 9873 33408
rect 9907 33405 9919 33439
rect 9861 33399 9919 33405
rect 10965 33439 11023 33445
rect 10965 33405 10977 33439
rect 11011 33436 11023 33439
rect 11054 33436 11060 33448
rect 11011 33408 11060 33436
rect 11011 33405 11023 33408
rect 10965 33399 11023 33405
rect 11054 33396 11060 33408
rect 11112 33436 11118 33448
rect 11514 33436 11520 33448
rect 11112 33408 11520 33436
rect 11112 33396 11118 33408
rect 11514 33396 11520 33408
rect 11572 33396 11578 33448
rect 9490 33328 9496 33380
rect 9548 33368 9554 33380
rect 9953 33371 10011 33377
rect 9953 33368 9965 33371
rect 9548 33340 9965 33368
rect 9548 33328 9554 33340
rect 9953 33337 9965 33340
rect 9999 33337 10011 33371
rect 9953 33331 10011 33337
rect 10410 33328 10416 33380
rect 10468 33368 10474 33380
rect 11808 33368 11836 33476
rect 11977 33473 11989 33476
rect 12023 33473 12035 33507
rect 11977 33467 12035 33473
rect 12158 33464 12164 33516
rect 12216 33464 12222 33516
rect 12434 33464 12440 33516
rect 12492 33464 12498 33516
rect 13081 33507 13139 33513
rect 13081 33473 13093 33507
rect 13127 33473 13139 33507
rect 13081 33467 13139 33473
rect 12345 33439 12403 33445
rect 12345 33436 12357 33439
rect 11992 33408 12357 33436
rect 11992 33380 12020 33408
rect 12345 33405 12357 33408
rect 12391 33405 12403 33439
rect 12345 33399 12403 33405
rect 12805 33439 12863 33445
rect 12805 33405 12817 33439
rect 12851 33436 12863 33439
rect 12986 33436 12992 33448
rect 12851 33408 12992 33436
rect 12851 33405 12863 33408
rect 12805 33399 12863 33405
rect 12986 33396 12992 33408
rect 13044 33396 13050 33448
rect 13096 33436 13124 33467
rect 13354 33464 13360 33516
rect 13412 33464 13418 33516
rect 13541 33507 13599 33513
rect 13541 33473 13553 33507
rect 13587 33504 13599 33507
rect 13633 33507 13691 33513
rect 13633 33504 13645 33507
rect 13587 33476 13645 33504
rect 13587 33473 13599 33476
rect 13541 33467 13599 33473
rect 13633 33473 13645 33476
rect 13679 33473 13691 33507
rect 13633 33467 13691 33473
rect 13814 33464 13820 33516
rect 13872 33464 13878 33516
rect 13998 33464 14004 33516
rect 14056 33464 14062 33516
rect 14182 33464 14188 33516
rect 14240 33464 14246 33516
rect 14366 33464 14372 33516
rect 14424 33464 14430 33516
rect 14458 33464 14464 33516
rect 14516 33464 14522 33516
rect 14553 33507 14611 33513
rect 14553 33473 14565 33507
rect 14599 33473 14611 33507
rect 14553 33467 14611 33473
rect 13722 33436 13728 33448
rect 13096 33408 13728 33436
rect 10468 33340 11836 33368
rect 10468 33328 10474 33340
rect 11974 33328 11980 33380
rect 12032 33328 12038 33380
rect 13096 33368 13124 33408
rect 13722 33396 13728 33408
rect 13780 33396 13786 33448
rect 13906 33396 13912 33448
rect 13964 33396 13970 33448
rect 14274 33396 14280 33448
rect 14332 33436 14338 33448
rect 14568 33436 14596 33467
rect 14734 33464 14740 33516
rect 14792 33464 14798 33516
rect 14936 33513 14964 33544
rect 15120 33544 15568 33572
rect 14921 33507 14979 33513
rect 14921 33473 14933 33507
rect 14967 33504 14979 33507
rect 15013 33507 15071 33513
rect 15013 33504 15025 33507
rect 14967 33476 15025 33504
rect 14967 33473 14979 33476
rect 14921 33467 14979 33473
rect 15013 33473 15025 33476
rect 15059 33473 15071 33507
rect 15013 33467 15071 33473
rect 15120 33436 15148 33544
rect 15562 33532 15568 33544
rect 15620 33532 15626 33584
rect 15194 33464 15200 33516
rect 15252 33504 15258 33516
rect 15381 33507 15439 33513
rect 15381 33504 15393 33507
rect 15252 33476 15393 33504
rect 15252 33464 15258 33476
rect 15381 33473 15393 33476
rect 15427 33473 15439 33507
rect 15672 33504 15700 33612
rect 16117 33609 16129 33643
rect 16163 33640 16175 33643
rect 16390 33640 16396 33652
rect 16163 33612 16396 33640
rect 16163 33609 16175 33612
rect 16117 33603 16175 33609
rect 16390 33600 16396 33612
rect 16448 33600 16454 33652
rect 18049 33643 18107 33649
rect 18049 33609 18061 33643
rect 18095 33640 18107 33643
rect 18322 33640 18328 33652
rect 18095 33612 18328 33640
rect 18095 33609 18107 33612
rect 18049 33603 18107 33609
rect 18322 33600 18328 33612
rect 18380 33600 18386 33652
rect 18506 33600 18512 33652
rect 18564 33640 18570 33652
rect 19242 33640 19248 33652
rect 18564 33612 19248 33640
rect 18564 33600 18570 33612
rect 19242 33600 19248 33612
rect 19300 33600 19306 33652
rect 20254 33600 20260 33652
rect 20312 33640 20318 33652
rect 20312 33612 20484 33640
rect 20312 33600 20318 33612
rect 15838 33532 15844 33584
rect 15896 33572 15902 33584
rect 15896 33544 16252 33572
rect 15896 33532 15902 33544
rect 15933 33507 15991 33513
rect 15933 33504 15945 33507
rect 15672 33476 15945 33504
rect 15381 33467 15439 33473
rect 15933 33473 15945 33476
rect 15979 33473 15991 33507
rect 15933 33467 15991 33473
rect 16114 33464 16120 33516
rect 16172 33464 16178 33516
rect 16224 33513 16252 33544
rect 16298 33532 16304 33584
rect 16356 33532 16362 33584
rect 16666 33532 16672 33584
rect 16724 33532 16730 33584
rect 18141 33575 18199 33581
rect 18141 33541 18153 33575
rect 18187 33572 18199 33575
rect 18966 33572 18972 33584
rect 18187 33544 18972 33572
rect 18187 33541 18199 33544
rect 18141 33535 18199 33541
rect 18966 33532 18972 33544
rect 19024 33532 19030 33584
rect 19061 33575 19119 33581
rect 19061 33541 19073 33575
rect 19107 33572 19119 33575
rect 19150 33572 19156 33584
rect 19107 33544 19156 33572
rect 19107 33541 19119 33544
rect 19061 33535 19119 33541
rect 19150 33532 19156 33544
rect 19208 33532 19214 33584
rect 20456 33572 20484 33612
rect 21818 33600 21824 33652
rect 21876 33640 21882 33652
rect 23014 33640 23020 33652
rect 21876 33612 23020 33640
rect 21876 33600 21882 33612
rect 23014 33600 23020 33612
rect 23072 33640 23078 33652
rect 23072 33612 23520 33640
rect 23072 33600 23078 33612
rect 20456 33544 20562 33572
rect 22554 33532 22560 33584
rect 22612 33532 22618 33584
rect 23492 33572 23520 33612
rect 24670 33600 24676 33652
rect 24728 33640 24734 33652
rect 25038 33640 25044 33652
rect 24728 33612 25044 33640
rect 24728 33600 24734 33612
rect 25038 33600 25044 33612
rect 25096 33640 25102 33652
rect 25774 33640 25780 33652
rect 25096 33612 25780 33640
rect 25096 33600 25102 33612
rect 25774 33600 25780 33612
rect 25832 33640 25838 33652
rect 26694 33640 26700 33652
rect 25832 33612 26700 33640
rect 25832 33600 25838 33612
rect 23492 33544 24256 33572
rect 16209 33507 16267 33513
rect 16209 33473 16221 33507
rect 16255 33473 16267 33507
rect 16209 33467 16267 33473
rect 16850 33464 16856 33516
rect 16908 33464 16914 33516
rect 18046 33464 18052 33516
rect 18104 33504 18110 33516
rect 18233 33507 18291 33513
rect 18233 33504 18245 33507
rect 18104 33476 18245 33504
rect 18104 33464 18110 33476
rect 18233 33473 18245 33476
rect 18279 33504 18291 33507
rect 18506 33504 18512 33516
rect 18279 33476 18512 33504
rect 18279 33473 18291 33476
rect 18233 33467 18291 33473
rect 18506 33464 18512 33476
rect 18564 33464 18570 33516
rect 18598 33464 18604 33516
rect 18656 33464 18662 33516
rect 18690 33464 18696 33516
rect 18748 33464 18754 33516
rect 18874 33464 18880 33516
rect 18932 33464 18938 33516
rect 24228 33513 24256 33544
rect 24394 33532 24400 33584
rect 24452 33572 24458 33584
rect 24765 33575 24823 33581
rect 24765 33572 24777 33575
rect 24452 33544 24777 33572
rect 24452 33532 24458 33544
rect 24765 33541 24777 33544
rect 24811 33541 24823 33575
rect 26252 33572 26280 33612
rect 26694 33600 26700 33612
rect 26752 33640 26758 33652
rect 29365 33643 29423 33649
rect 29365 33640 29377 33643
rect 26752 33612 29377 33640
rect 26752 33600 26758 33612
rect 29365 33609 29377 33612
rect 29411 33609 29423 33643
rect 29365 33603 29423 33609
rect 32306 33600 32312 33652
rect 32364 33640 32370 33652
rect 33873 33643 33931 33649
rect 33873 33640 33885 33643
rect 32364 33612 33885 33640
rect 32364 33600 32370 33612
rect 33873 33609 33885 33612
rect 33919 33609 33931 33643
rect 33873 33603 33931 33609
rect 25990 33544 26280 33572
rect 27157 33575 27215 33581
rect 24765 33535 24823 33541
rect 27157 33541 27169 33575
rect 27203 33572 27215 33575
rect 27982 33572 27988 33584
rect 27203 33544 27988 33572
rect 27203 33541 27215 33544
rect 27157 33535 27215 33541
rect 27982 33532 27988 33544
rect 28040 33532 28046 33584
rect 29914 33572 29920 33584
rect 29012 33544 29920 33572
rect 29012 33516 29040 33544
rect 29914 33532 29920 33544
rect 29972 33572 29978 33584
rect 29972 33544 30222 33572
rect 29972 33532 29978 33544
rect 32858 33532 32864 33584
rect 32916 33532 32922 33584
rect 19521 33507 19579 33513
rect 19521 33504 19533 33507
rect 19168 33476 19533 33504
rect 19168 33448 19196 33476
rect 19521 33473 19533 33476
rect 19567 33473 19579 33507
rect 19521 33467 19579 33473
rect 19705 33507 19763 33513
rect 19705 33473 19717 33507
rect 19751 33504 19763 33507
rect 20165 33507 20223 33513
rect 20165 33504 20177 33507
rect 19751 33476 20177 33504
rect 19751 33473 19763 33476
rect 19705 33467 19763 33473
rect 20165 33473 20177 33476
rect 20211 33473 20223 33507
rect 20165 33467 20223 33473
rect 23569 33507 23627 33513
rect 23569 33473 23581 33507
rect 23615 33473 23627 33507
rect 23569 33467 23627 33473
rect 24213 33507 24271 33513
rect 24213 33473 24225 33507
rect 24259 33473 24271 33507
rect 24213 33467 24271 33473
rect 14332 33408 15148 33436
rect 14332 33396 14338 33408
rect 15286 33396 15292 33448
rect 15344 33436 15350 33448
rect 17773 33439 17831 33445
rect 17773 33436 17785 33439
rect 15344 33408 17785 33436
rect 15344 33396 15350 33408
rect 17773 33405 17785 33408
rect 17819 33436 17831 33439
rect 18414 33436 18420 33448
rect 17819 33408 18420 33436
rect 17819 33405 17831 33408
rect 17773 33399 17831 33405
rect 18414 33396 18420 33408
rect 18472 33396 18478 33448
rect 18782 33396 18788 33448
rect 18840 33436 18846 33448
rect 18969 33439 19027 33445
rect 18969 33436 18981 33439
rect 18840 33408 18981 33436
rect 18840 33396 18846 33408
rect 18969 33405 18981 33408
rect 19015 33405 19027 33439
rect 18969 33399 19027 33405
rect 19150 33396 19156 33448
rect 19208 33396 19214 33448
rect 19337 33439 19395 33445
rect 19337 33405 19349 33439
rect 19383 33436 19395 33439
rect 19426 33436 19432 33448
rect 19383 33408 19432 33436
rect 19383 33405 19395 33408
rect 19337 33399 19395 33405
rect 19426 33396 19432 33408
rect 19484 33396 19490 33448
rect 19797 33439 19855 33445
rect 19797 33405 19809 33439
rect 19843 33405 19855 33439
rect 19797 33399 19855 33405
rect 12406 33340 13124 33368
rect 8628 33272 9352 33300
rect 8628 33260 8634 33272
rect 9398 33260 9404 33312
rect 9456 33300 9462 33312
rect 12406 33300 12434 33340
rect 13262 33328 13268 33380
rect 13320 33368 13326 33380
rect 13924 33368 13952 33396
rect 13320 33340 13952 33368
rect 13320 33328 13326 33340
rect 14090 33328 14096 33380
rect 14148 33368 14154 33380
rect 15197 33371 15255 33377
rect 15197 33368 15209 33371
rect 14148 33340 15209 33368
rect 14148 33328 14154 33340
rect 15197 33337 15209 33340
rect 15243 33337 15255 33371
rect 15197 33331 15255 33337
rect 15562 33328 15568 33380
rect 15620 33328 15626 33380
rect 18690 33328 18696 33380
rect 18748 33368 18754 33380
rect 19518 33368 19524 33380
rect 18748 33340 19524 33368
rect 18748 33328 18754 33340
rect 19518 33328 19524 33340
rect 19576 33368 19582 33380
rect 19812 33368 19840 33399
rect 22738 33396 22744 33448
rect 22796 33436 22802 33448
rect 23293 33439 23351 33445
rect 23293 33436 23305 33439
rect 22796 33408 23305 33436
rect 22796 33396 22802 33408
rect 23293 33405 23305 33408
rect 23339 33405 23351 33439
rect 23584 33436 23612 33467
rect 26050 33464 26056 33516
rect 26108 33504 26114 33516
rect 26329 33507 26387 33513
rect 26329 33504 26341 33507
rect 26108 33476 26341 33504
rect 26108 33464 26114 33476
rect 26329 33473 26341 33476
rect 26375 33473 26387 33507
rect 27341 33507 27399 33513
rect 27341 33504 27353 33507
rect 26329 33467 26387 33473
rect 27172 33476 27353 33504
rect 27172 33448 27200 33476
rect 27341 33473 27353 33476
rect 27387 33473 27399 33507
rect 27341 33467 27399 33473
rect 27430 33464 27436 33516
rect 27488 33464 27494 33516
rect 28994 33504 29000 33516
rect 28842 33490 29000 33504
rect 28828 33476 29000 33490
rect 23293 33399 23351 33405
rect 23492 33408 23612 33436
rect 24489 33439 24547 33445
rect 19576 33340 19840 33368
rect 19576 33328 19582 33340
rect 9456 33272 12434 33300
rect 9456 33260 9462 33272
rect 13906 33260 13912 33312
rect 13964 33300 13970 33312
rect 14642 33300 14648 33312
rect 13964 33272 14648 33300
rect 13964 33260 13970 33272
rect 14642 33260 14648 33272
rect 14700 33300 14706 33312
rect 15105 33303 15163 33309
rect 15105 33300 15117 33303
rect 14700 33272 15117 33300
rect 14700 33260 14706 33272
rect 15105 33269 15117 33272
rect 15151 33269 15163 33303
rect 15105 33263 15163 33269
rect 19426 33260 19432 33312
rect 19484 33300 19490 33312
rect 21591 33303 21649 33309
rect 21591 33300 21603 33303
rect 19484 33272 21603 33300
rect 19484 33260 19490 33272
rect 21591 33269 21603 33272
rect 21637 33300 21649 33303
rect 22278 33300 22284 33312
rect 21637 33272 22284 33300
rect 21637 33269 21649 33272
rect 21591 33263 21649 33269
rect 22278 33260 22284 33272
rect 22336 33260 22342 33312
rect 23198 33260 23204 33312
rect 23256 33300 23262 33312
rect 23492 33300 23520 33408
rect 24489 33405 24501 33439
rect 24535 33436 24547 33439
rect 25498 33436 25504 33448
rect 24535 33408 25504 33436
rect 24535 33405 24547 33408
rect 24489 33399 24547 33405
rect 25498 33396 25504 33408
rect 25556 33396 25562 33448
rect 25958 33396 25964 33448
rect 26016 33436 26022 33448
rect 26418 33436 26424 33448
rect 26016 33408 26424 33436
rect 26016 33396 26022 33408
rect 26418 33396 26424 33408
rect 26476 33436 26482 33448
rect 26513 33439 26571 33445
rect 26513 33436 26525 33439
rect 26476 33408 26525 33436
rect 26476 33396 26482 33408
rect 26513 33405 26525 33408
rect 26559 33405 26571 33439
rect 26513 33399 26571 33405
rect 27154 33396 27160 33448
rect 27212 33396 27218 33448
rect 27706 33396 27712 33448
rect 27764 33396 27770 33448
rect 26878 33328 26884 33380
rect 26936 33368 26942 33380
rect 26936 33340 27568 33368
rect 26936 33328 26942 33340
rect 23256 33272 23520 33300
rect 23256 33260 23262 33272
rect 23658 33260 23664 33312
rect 23716 33260 23722 33312
rect 26234 33260 26240 33312
rect 26292 33260 26298 33312
rect 26602 33260 26608 33312
rect 26660 33300 26666 33312
rect 26973 33303 27031 33309
rect 26973 33300 26985 33303
rect 26660 33272 26985 33300
rect 26660 33260 26666 33272
rect 26973 33269 26985 33272
rect 27019 33269 27031 33303
rect 27540 33300 27568 33340
rect 28828 33300 28856 33476
rect 28994 33464 29000 33476
rect 29052 33464 29058 33516
rect 29454 33464 29460 33516
rect 29512 33464 29518 33516
rect 31662 33464 31668 33516
rect 31720 33504 31726 33516
rect 32125 33507 32183 33513
rect 32125 33504 32137 33507
rect 31720 33476 32137 33504
rect 31720 33464 31726 33476
rect 32125 33473 32137 33476
rect 32171 33473 32183 33507
rect 32125 33467 32183 33473
rect 29178 33396 29184 33448
rect 29236 33396 29242 33448
rect 29638 33396 29644 33448
rect 29696 33396 29702 33448
rect 31386 33396 31392 33448
rect 31444 33396 31450 33448
rect 32398 33396 32404 33448
rect 32456 33396 32462 33448
rect 27540 33272 28856 33300
rect 26973 33263 27031 33269
rect 29362 33260 29368 33312
rect 29420 33300 29426 33312
rect 32214 33300 32220 33312
rect 29420 33272 32220 33300
rect 29420 33260 29426 33272
rect 32214 33260 32220 33272
rect 32272 33260 32278 33312
rect 1104 33210 36432 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 36432 33210
rect 1104 33136 36432 33158
rect 4525 33099 4583 33105
rect 4525 33065 4537 33099
rect 4571 33096 4583 33099
rect 5074 33096 5080 33108
rect 4571 33068 5080 33096
rect 4571 33065 4583 33068
rect 4525 33059 4583 33065
rect 3973 33031 4031 33037
rect 3973 32997 3985 33031
rect 4019 33028 4031 33031
rect 4430 33028 4436 33040
rect 4019 33000 4436 33028
rect 4019 32997 4031 33000
rect 3973 32991 4031 32997
rect 4430 32988 4436 33000
rect 4488 32988 4494 33040
rect 4540 32960 4568 33059
rect 5074 33056 5080 33068
rect 5132 33056 5138 33108
rect 5258 33056 5264 33108
rect 5316 33056 5322 33108
rect 5445 33099 5503 33105
rect 5445 33065 5457 33099
rect 5491 33096 5503 33099
rect 5534 33096 5540 33108
rect 5491 33068 5540 33096
rect 5491 33065 5503 33068
rect 5445 33059 5503 33065
rect 5534 33056 5540 33068
rect 5592 33056 5598 33108
rect 6178 33056 6184 33108
rect 6236 33096 6242 33108
rect 6236 33068 6408 33096
rect 6236 33056 6242 33068
rect 4709 33031 4767 33037
rect 4709 32997 4721 33031
rect 4755 33028 4767 33031
rect 5166 33028 5172 33040
rect 4755 33000 5172 33028
rect 4755 32997 4767 33000
rect 4709 32991 4767 32997
rect 5166 32988 5172 33000
rect 5224 32988 5230 33040
rect 5675 33031 5733 33037
rect 5675 32997 5687 33031
rect 5721 32997 5733 33031
rect 6380 33028 6408 33068
rect 6454 33056 6460 33108
rect 6512 33056 6518 33108
rect 6546 33056 6552 33108
rect 6604 33056 6610 33108
rect 6638 33056 6644 33108
rect 6696 33096 6702 33108
rect 7190 33096 7196 33108
rect 6696 33068 7196 33096
rect 6696 33056 6702 33068
rect 7190 33056 7196 33068
rect 7248 33056 7254 33108
rect 7282 33056 7288 33108
rect 7340 33056 7346 33108
rect 7837 33099 7895 33105
rect 7837 33065 7849 33099
rect 7883 33096 7895 33099
rect 8110 33096 8116 33108
rect 7883 33068 8116 33096
rect 7883 33065 7895 33068
rect 7837 33059 7895 33065
rect 8110 33056 8116 33068
rect 8168 33056 8174 33108
rect 9401 33099 9459 33105
rect 9401 33065 9413 33099
rect 9447 33096 9459 33099
rect 10226 33096 10232 33108
rect 9447 33068 10232 33096
rect 9447 33065 9459 33068
rect 9401 33059 9459 33065
rect 10226 33056 10232 33068
rect 10284 33056 10290 33108
rect 10962 33056 10968 33108
rect 11020 33096 11026 33108
rect 12161 33099 12219 33105
rect 11020 33068 12112 33096
rect 11020 33056 11026 33068
rect 6380 33000 7236 33028
rect 5675 32991 5733 32997
rect 4172 32932 4568 32960
rect 3326 32852 3332 32904
rect 3384 32892 3390 32904
rect 4172 32901 4200 32932
rect 4798 32920 4804 32972
rect 4856 32920 4862 32972
rect 4893 32963 4951 32969
rect 4893 32929 4905 32963
rect 4939 32960 4951 32963
rect 5537 32963 5595 32969
rect 5537 32960 5549 32963
rect 4939 32932 5549 32960
rect 4939 32929 4951 32932
rect 4893 32923 4951 32929
rect 5276 32904 5304 32932
rect 5537 32929 5549 32932
rect 5583 32929 5595 32963
rect 5690 32960 5718 32991
rect 6546 32960 6552 32972
rect 5537 32923 5595 32929
rect 5644 32932 5718 32960
rect 6012 32932 6552 32960
rect 5644 32904 5672 32932
rect 4157 32895 4215 32901
rect 4157 32892 4169 32895
rect 3384 32864 4169 32892
rect 3384 32852 3390 32864
rect 4157 32861 4169 32864
rect 4203 32861 4215 32895
rect 4157 32855 4215 32861
rect 4249 32895 4307 32901
rect 4249 32861 4261 32895
rect 4295 32892 4307 32895
rect 4295 32864 4568 32892
rect 4295 32861 4307 32864
rect 4249 32855 4307 32861
rect 2958 32784 2964 32836
rect 3016 32824 3022 32836
rect 3973 32827 4031 32833
rect 3973 32824 3985 32827
rect 3016 32796 3985 32824
rect 3016 32784 3022 32796
rect 3973 32793 3985 32796
rect 4019 32824 4031 32827
rect 4338 32824 4344 32836
rect 4019 32796 4344 32824
rect 4019 32793 4031 32796
rect 3973 32787 4031 32793
rect 4338 32784 4344 32796
rect 4396 32784 4402 32836
rect 4540 32833 4568 32864
rect 5074 32852 5080 32904
rect 5132 32852 5138 32904
rect 5258 32852 5264 32904
rect 5316 32852 5322 32904
rect 5353 32895 5411 32901
rect 5353 32861 5365 32895
rect 5399 32892 5411 32895
rect 5442 32892 5448 32904
rect 5399 32864 5448 32892
rect 5399 32861 5411 32864
rect 5353 32855 5411 32861
rect 5442 32852 5448 32864
rect 5500 32852 5506 32904
rect 5626 32852 5632 32904
rect 5684 32852 5690 32904
rect 5810 32852 5816 32904
rect 5868 32852 5874 32904
rect 5902 32852 5908 32904
rect 5960 32892 5966 32904
rect 6012 32901 6040 32932
rect 6546 32920 6552 32932
rect 6604 32920 6610 32972
rect 6638 32920 6644 32972
rect 6696 32920 6702 32972
rect 6730 32920 6736 32972
rect 6788 32920 6794 32972
rect 5997 32895 6055 32901
rect 5997 32892 6009 32895
rect 5960 32864 6009 32892
rect 5960 32852 5966 32864
rect 5997 32861 6009 32864
rect 6043 32861 6055 32895
rect 5997 32855 6055 32861
rect 6086 32852 6092 32904
rect 6144 32852 6150 32904
rect 6178 32852 6184 32904
rect 6236 32892 6242 32904
rect 6273 32895 6331 32901
rect 6273 32892 6285 32895
rect 6236 32864 6285 32892
rect 6236 32852 6242 32864
rect 6273 32861 6285 32864
rect 6319 32861 6331 32895
rect 6273 32855 6331 32861
rect 4540 32827 4615 32833
rect 4540 32796 4569 32827
rect 4557 32793 4569 32796
rect 4603 32824 4615 32827
rect 6549 32827 6607 32833
rect 4603 32796 4844 32824
rect 4603 32793 4615 32796
rect 4557 32787 4615 32793
rect 4816 32768 4844 32796
rect 6549 32793 6561 32827
rect 6595 32824 6607 32827
rect 6638 32824 6644 32836
rect 6595 32796 6644 32824
rect 6595 32793 6607 32796
rect 6549 32787 6607 32793
rect 4798 32716 4804 32768
rect 4856 32716 4862 32768
rect 5074 32716 5080 32768
rect 5132 32756 5138 32768
rect 5810 32756 5816 32768
rect 5132 32728 5816 32756
rect 5132 32716 5138 32728
rect 5810 32716 5816 32728
rect 5868 32716 5874 32768
rect 6086 32716 6092 32768
rect 6144 32756 6150 32768
rect 6564 32756 6592 32787
rect 6638 32784 6644 32796
rect 6696 32784 6702 32836
rect 6748 32768 6776 32920
rect 6825 32895 6883 32901
rect 6825 32861 6837 32895
rect 6871 32861 6883 32895
rect 6825 32855 6883 32861
rect 6840 32824 6868 32855
rect 7098 32852 7104 32904
rect 7156 32852 7162 32904
rect 7208 32892 7236 33000
rect 7374 32988 7380 33040
rect 7432 33028 7438 33040
rect 9953 33031 10011 33037
rect 7432 33000 9352 33028
rect 7432 32988 7438 33000
rect 8754 32960 8760 32972
rect 8312 32932 8760 32960
rect 7285 32895 7343 32901
rect 7285 32892 7297 32895
rect 7208 32864 7297 32892
rect 7285 32861 7297 32864
rect 7331 32861 7343 32895
rect 7285 32855 7343 32861
rect 7561 32895 7619 32901
rect 7561 32861 7573 32895
rect 7607 32892 7619 32895
rect 7926 32892 7932 32904
rect 7607 32864 7932 32892
rect 7607 32861 7619 32864
rect 7561 32855 7619 32861
rect 7926 32852 7932 32864
rect 7984 32852 7990 32904
rect 8018 32852 8024 32904
rect 8076 32852 8082 32904
rect 8312 32901 8340 32932
rect 8754 32920 8760 32932
rect 8812 32920 8818 32972
rect 9324 32960 9352 33000
rect 9953 32997 9965 33031
rect 9999 33028 10011 33031
rect 10042 33028 10048 33040
rect 9999 33000 10048 33028
rect 9999 32997 10011 33000
rect 9953 32991 10011 32997
rect 10042 32988 10048 33000
rect 10100 32988 10106 33040
rect 10134 32988 10140 33040
rect 10192 33028 10198 33040
rect 12084 33028 12112 33068
rect 12161 33065 12173 33099
rect 12207 33096 12219 33099
rect 12250 33096 12256 33108
rect 12207 33068 12256 33096
rect 12207 33065 12219 33068
rect 12161 33059 12219 33065
rect 12250 33056 12256 33068
rect 12308 33056 12314 33108
rect 18230 33096 18236 33108
rect 12406 33068 18236 33096
rect 12406 33028 12434 33068
rect 18230 33056 18236 33068
rect 18288 33056 18294 33108
rect 18322 33056 18328 33108
rect 18380 33096 18386 33108
rect 19521 33099 19579 33105
rect 19521 33096 19533 33099
rect 18380 33068 19533 33096
rect 18380 33056 18386 33068
rect 19521 33065 19533 33068
rect 19567 33065 19579 33099
rect 19521 33059 19579 33065
rect 22094 33056 22100 33108
rect 22152 33096 22158 33108
rect 22152 33068 22232 33096
rect 22152 33056 22158 33068
rect 10192 33000 11468 33028
rect 12084 33000 12434 33028
rect 10192 32988 10198 33000
rect 9674 32960 9680 32972
rect 9324 32932 9680 32960
rect 8113 32895 8171 32901
rect 8113 32861 8125 32895
rect 8159 32861 8171 32895
rect 8113 32855 8171 32861
rect 8297 32895 8355 32901
rect 8297 32861 8309 32895
rect 8343 32861 8355 32895
rect 8297 32855 8355 32861
rect 7742 32824 7748 32836
rect 6840 32796 7748 32824
rect 6840 32768 6868 32796
rect 7742 32784 7748 32796
rect 7800 32784 7806 32836
rect 8128 32824 8156 32855
rect 8386 32852 8392 32904
rect 8444 32852 8450 32904
rect 9324 32901 9352 32932
rect 9674 32920 9680 32932
rect 9732 32920 9738 32972
rect 10226 32960 10232 32972
rect 10060 32932 10232 32960
rect 9309 32895 9367 32901
rect 9309 32861 9321 32895
rect 9355 32861 9367 32895
rect 9309 32855 9367 32861
rect 9490 32852 9496 32904
rect 9548 32852 9554 32904
rect 10060 32901 10088 32932
rect 10226 32920 10232 32932
rect 10284 32960 10290 32972
rect 11330 32960 11336 32972
rect 10284 32932 11336 32960
rect 10284 32920 10290 32932
rect 11330 32920 11336 32932
rect 11388 32920 11394 32972
rect 10045 32895 10103 32901
rect 10045 32861 10057 32895
rect 10091 32861 10103 32895
rect 10045 32855 10103 32861
rect 10137 32895 10195 32901
rect 10137 32861 10149 32895
rect 10183 32861 10195 32895
rect 10137 32855 10195 32861
rect 8754 32824 8760 32836
rect 8128 32796 8760 32824
rect 8754 32784 8760 32796
rect 8812 32784 8818 32836
rect 9766 32784 9772 32836
rect 9824 32784 9830 32836
rect 10152 32824 10180 32855
rect 10318 32852 10324 32904
rect 10376 32852 10382 32904
rect 10502 32852 10508 32904
rect 10560 32892 10566 32904
rect 10962 32892 10968 32904
rect 10560 32864 10968 32892
rect 10560 32852 10566 32864
rect 10962 32852 10968 32864
rect 11020 32892 11026 32904
rect 11241 32895 11299 32901
rect 11241 32892 11253 32895
rect 11020 32864 11253 32892
rect 11020 32852 11026 32864
rect 11241 32861 11253 32864
rect 11287 32861 11299 32895
rect 11440 32892 11468 33000
rect 15838 32988 15844 33040
rect 15896 33028 15902 33040
rect 15896 33000 20299 33028
rect 15896 32988 15902 33000
rect 13832 32932 15608 32960
rect 11977 32895 12035 32901
rect 11977 32892 11989 32895
rect 11440 32864 11989 32892
rect 11241 32855 11299 32861
rect 11977 32861 11989 32864
rect 12023 32892 12035 32895
rect 12158 32892 12164 32904
rect 12023 32864 12164 32892
rect 12023 32861 12035 32864
rect 11977 32855 12035 32861
rect 12158 32852 12164 32864
rect 12216 32852 12222 32904
rect 10060 32796 10180 32824
rect 6144 32728 6592 32756
rect 6144 32716 6150 32728
rect 6730 32716 6736 32768
rect 6788 32716 6794 32768
rect 6822 32716 6828 32768
rect 6880 32716 6886 32768
rect 7009 32759 7067 32765
rect 7009 32725 7021 32759
rect 7055 32756 7067 32759
rect 9950 32756 9956 32768
rect 7055 32728 9956 32756
rect 7055 32725 7067 32728
rect 7009 32719 7067 32725
rect 9950 32716 9956 32728
rect 10008 32716 10014 32768
rect 10060 32765 10088 32796
rect 10410 32784 10416 32836
rect 10468 32824 10474 32836
rect 11793 32827 11851 32833
rect 11793 32824 11805 32827
rect 10468 32796 11805 32824
rect 10468 32784 10474 32796
rect 11793 32793 11805 32796
rect 11839 32793 11851 32827
rect 11793 32787 11851 32793
rect 10045 32759 10103 32765
rect 10045 32725 10057 32759
rect 10091 32725 10103 32759
rect 10045 32719 10103 32725
rect 10226 32716 10232 32768
rect 10284 32716 10290 32768
rect 10962 32716 10968 32768
rect 11020 32756 11026 32768
rect 11149 32759 11207 32765
rect 11149 32756 11161 32759
rect 11020 32728 11161 32756
rect 11020 32716 11026 32728
rect 11149 32725 11161 32728
rect 11195 32725 11207 32759
rect 11808 32756 11836 32787
rect 13832 32756 13860 32932
rect 14090 32852 14096 32904
rect 14148 32852 14154 32904
rect 15580 32892 15608 32932
rect 16114 32920 16120 32972
rect 16172 32960 16178 32972
rect 19886 32960 19892 32972
rect 16172 32932 19892 32960
rect 16172 32920 16178 32932
rect 19886 32920 19892 32932
rect 19944 32920 19950 32972
rect 20271 32904 20299 33000
rect 22104 32963 22162 32969
rect 22104 32929 22116 32963
rect 22150 32960 22162 32963
rect 22204 32960 22232 33068
rect 22462 33056 22468 33108
rect 22520 33096 22526 33108
rect 24486 33096 24492 33108
rect 22520 33068 24492 33096
rect 22520 33056 22526 33068
rect 24486 33056 24492 33068
rect 24544 33056 24550 33108
rect 24854 33056 24860 33108
rect 24912 33096 24918 33108
rect 25225 33099 25283 33105
rect 25225 33096 25237 33099
rect 24912 33068 25237 33096
rect 24912 33056 24918 33068
rect 25225 33065 25237 33068
rect 25271 33065 25283 33099
rect 29638 33096 29644 33108
rect 25225 33059 25283 33065
rect 25332 33068 29644 33096
rect 24029 33031 24087 33037
rect 24029 32997 24041 33031
rect 24075 33028 24087 33031
rect 24118 33028 24124 33040
rect 24075 33000 24124 33028
rect 24075 32997 24087 33000
rect 24029 32991 24087 32997
rect 24118 32988 24124 33000
rect 24176 32988 24182 33040
rect 24578 32988 24584 33040
rect 24636 33028 24642 33040
rect 25332 33028 25360 33068
rect 29638 33056 29644 33068
rect 29696 33096 29702 33108
rect 29696 33068 31248 33096
rect 29696 33056 29702 33068
rect 24636 33000 25360 33028
rect 27617 33031 27675 33037
rect 24636 32988 24642 33000
rect 27617 32997 27629 33031
rect 27663 32997 27675 33031
rect 27617 32991 27675 32997
rect 22150 32932 22232 32960
rect 22150 32929 22162 32932
rect 22104 32923 22162 32929
rect 22370 32920 22376 32972
rect 22428 32920 22434 32972
rect 23382 32920 23388 32972
rect 23440 32960 23446 32972
rect 23658 32960 23664 32972
rect 23440 32932 23664 32960
rect 23440 32920 23446 32932
rect 23658 32920 23664 32932
rect 23716 32920 23722 32972
rect 25133 32968 25191 32969
rect 25133 32963 25268 32968
rect 25133 32929 25145 32963
rect 25179 32940 25268 32963
rect 25179 32929 25191 32940
rect 25133 32923 25191 32929
rect 16574 32892 16580 32904
rect 15580 32864 16580 32892
rect 16574 32852 16580 32864
rect 16632 32852 16638 32904
rect 19429 32895 19487 32901
rect 19429 32861 19441 32895
rect 19475 32892 19487 32895
rect 20070 32892 20076 32904
rect 19475 32864 20076 32892
rect 19475 32861 19487 32864
rect 19429 32855 19487 32861
rect 20070 32852 20076 32864
rect 20128 32852 20134 32904
rect 20254 32892 20260 32904
rect 20215 32864 20260 32892
rect 20254 32852 20260 32864
rect 20312 32852 20318 32904
rect 20349 32895 20407 32901
rect 20349 32861 20361 32895
rect 20395 32861 20407 32895
rect 20349 32855 20407 32861
rect 14366 32784 14372 32836
rect 14424 32784 14430 32836
rect 14918 32784 14924 32836
rect 14976 32784 14982 32836
rect 16117 32827 16175 32833
rect 16117 32793 16129 32827
rect 16163 32793 16175 32827
rect 16117 32787 16175 32793
rect 11808 32728 13860 32756
rect 11149 32719 11207 32725
rect 14182 32716 14188 32768
rect 14240 32756 14246 32768
rect 16132 32756 16160 32787
rect 19242 32784 19248 32836
rect 19300 32824 19306 32836
rect 19705 32827 19763 32833
rect 19705 32824 19717 32827
rect 19300 32796 19717 32824
rect 19300 32784 19306 32796
rect 19705 32793 19717 32796
rect 19751 32793 19763 32827
rect 19705 32787 19763 32793
rect 19889 32827 19947 32833
rect 19889 32793 19901 32827
rect 19935 32793 19947 32827
rect 20364 32824 20392 32855
rect 21818 32852 21824 32904
rect 21876 32852 21882 32904
rect 24026 32852 24032 32904
rect 24084 32892 24090 32904
rect 24213 32895 24271 32901
rect 24213 32892 24225 32895
rect 24084 32864 24225 32892
rect 24084 32852 24090 32864
rect 24213 32861 24225 32864
rect 24259 32861 24271 32895
rect 24213 32855 24271 32861
rect 24394 32852 24400 32904
rect 24452 32852 24458 32904
rect 24670 32852 24676 32904
rect 24728 32852 24734 32904
rect 24854 32852 24860 32904
rect 24912 32901 24918 32904
rect 24912 32895 24974 32901
rect 24912 32861 24928 32895
rect 24962 32892 24974 32895
rect 25038 32892 25044 32904
rect 24962 32864 25044 32892
rect 24962 32861 24974 32864
rect 24912 32855 24974 32861
rect 24912 32852 24918 32855
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 20714 32824 20720 32836
rect 20364 32796 20720 32824
rect 19889 32787 19947 32793
rect 14240 32728 16160 32756
rect 14240 32716 14246 32728
rect 19334 32716 19340 32768
rect 19392 32716 19398 32768
rect 19904 32756 19932 32787
rect 20714 32784 20720 32796
rect 20772 32824 20778 32836
rect 21910 32824 21916 32836
rect 20772 32796 21916 32824
rect 20772 32784 20778 32796
rect 21910 32784 21916 32796
rect 21968 32784 21974 32836
rect 22005 32827 22063 32833
rect 22005 32793 22017 32827
rect 22051 32793 22063 32827
rect 24688 32824 24716 32852
rect 25240 32824 25268 32940
rect 25314 32920 25320 32972
rect 25372 32960 25378 32972
rect 27632 32960 27660 32991
rect 28258 32988 28264 33040
rect 28316 32988 28322 33040
rect 28350 32988 28356 33040
rect 28408 33028 28414 33040
rect 29549 33031 29607 33037
rect 29549 33028 29561 33031
rect 28408 33000 29561 33028
rect 28408 32988 28414 33000
rect 29549 32997 29561 33000
rect 29595 33028 29607 33031
rect 30006 33028 30012 33040
rect 29595 33000 30012 33028
rect 29595 32997 29607 33000
rect 29549 32991 29607 32997
rect 30006 32988 30012 33000
rect 30064 32988 30070 33040
rect 31220 33028 31248 33068
rect 31386 33056 31392 33108
rect 31444 33056 31450 33108
rect 32033 33099 32091 33105
rect 32033 33065 32045 33099
rect 32079 33096 32091 33099
rect 32398 33096 32404 33108
rect 32079 33068 32404 33096
rect 32079 33065 32091 33068
rect 32033 33059 32091 33065
rect 32398 33056 32404 33068
rect 32456 33056 32462 33108
rect 31220 33000 31784 33028
rect 27706 32960 27712 32972
rect 25372 32932 27568 32960
rect 27632 32932 27712 32960
rect 25372 32920 25378 32932
rect 27540 32904 27568 32932
rect 27706 32920 27712 32932
rect 27764 32920 27770 32972
rect 29178 32960 29184 32972
rect 28000 32932 29184 32960
rect 25406 32852 25412 32904
rect 25464 32852 25470 32904
rect 25498 32852 25504 32904
rect 25556 32852 25562 32904
rect 25774 32852 25780 32904
rect 25832 32892 25838 32904
rect 25869 32895 25927 32901
rect 25869 32892 25881 32895
rect 25832 32864 25881 32892
rect 25832 32852 25838 32864
rect 25869 32861 25881 32864
rect 25915 32861 25927 32895
rect 25869 32855 25927 32861
rect 27522 32852 27528 32904
rect 27580 32892 27586 32904
rect 27801 32895 27859 32901
rect 27801 32892 27813 32895
rect 27580 32864 27813 32892
rect 27580 32852 27586 32864
rect 27801 32861 27813 32864
rect 27847 32861 27859 32895
rect 27801 32855 27859 32861
rect 23598 32796 24716 32824
rect 25056 32796 25268 32824
rect 22005 32787 22063 32793
rect 19978 32756 19984 32768
rect 19904 32728 19984 32756
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 21637 32759 21695 32765
rect 21637 32725 21649 32759
rect 21683 32756 21695 32759
rect 21726 32756 21732 32768
rect 21683 32728 21732 32756
rect 21683 32725 21695 32728
rect 21637 32719 21695 32725
rect 21726 32716 21732 32728
rect 21784 32716 21790 32768
rect 22020 32756 22048 32787
rect 23658 32756 23664 32768
rect 22020 32728 23664 32756
rect 23658 32716 23664 32728
rect 23716 32716 23722 32768
rect 23845 32759 23903 32765
rect 23845 32725 23857 32759
rect 23891 32756 23903 32759
rect 24026 32756 24032 32768
rect 23891 32728 24032 32756
rect 23891 32725 23903 32728
rect 23845 32719 23903 32725
rect 24026 32716 24032 32728
rect 24084 32716 24090 32768
rect 24857 32759 24915 32765
rect 24857 32725 24869 32759
rect 24903 32756 24915 32759
rect 24946 32756 24952 32768
rect 24903 32728 24952 32756
rect 24903 32725 24915 32728
rect 24857 32719 24915 32725
rect 24946 32716 24952 32728
rect 25004 32716 25010 32768
rect 25056 32765 25084 32796
rect 26694 32784 26700 32836
rect 26752 32784 26758 32836
rect 27816 32824 27844 32855
rect 27890 32852 27896 32904
rect 27948 32852 27954 32904
rect 28000 32901 28028 32932
rect 29178 32920 29184 32932
rect 29236 32920 29242 32972
rect 29270 32920 29276 32972
rect 29328 32920 29334 32972
rect 31297 32963 31355 32969
rect 31297 32929 31309 32963
rect 31343 32960 31355 32963
rect 31662 32960 31668 32972
rect 31343 32932 31668 32960
rect 31343 32929 31355 32932
rect 31297 32923 31355 32929
rect 31662 32920 31668 32932
rect 31720 32920 31726 32972
rect 27985 32895 28043 32901
rect 27985 32861 27997 32895
rect 28031 32861 28043 32895
rect 27985 32855 28043 32861
rect 28074 32852 28080 32904
rect 28132 32892 28138 32904
rect 28169 32895 28227 32901
rect 28169 32892 28181 32895
rect 28132 32864 28181 32892
rect 28132 32852 28138 32864
rect 28169 32861 28181 32864
rect 28215 32861 28227 32895
rect 28169 32855 28227 32861
rect 28445 32895 28503 32901
rect 28445 32861 28457 32895
rect 28491 32861 28503 32895
rect 28445 32855 28503 32861
rect 28460 32824 28488 32855
rect 28534 32852 28540 32904
rect 28592 32852 28598 32904
rect 28810 32852 28816 32904
rect 28868 32852 28874 32904
rect 28994 32852 29000 32904
rect 29052 32892 29058 32904
rect 29089 32895 29147 32901
rect 29089 32892 29101 32895
rect 29052 32864 29101 32892
rect 29052 32852 29058 32864
rect 29089 32861 29101 32864
rect 29135 32861 29147 32895
rect 29089 32855 29147 32861
rect 29914 32852 29920 32904
rect 29972 32852 29978 32904
rect 31570 32852 31576 32904
rect 31628 32852 31634 32904
rect 31756 32892 31784 33000
rect 32122 32920 32128 32972
rect 32180 32960 32186 32972
rect 32309 32963 32367 32969
rect 32309 32960 32321 32963
rect 32180 32932 32321 32960
rect 32180 32920 32186 32932
rect 32309 32929 32321 32932
rect 32355 32960 32367 32963
rect 33045 32963 33103 32969
rect 33045 32960 33057 32963
rect 32355 32932 33057 32960
rect 32355 32929 32367 32932
rect 32309 32923 32367 32929
rect 33045 32929 33057 32932
rect 33091 32929 33103 32963
rect 33045 32923 33103 32929
rect 31680 32864 31784 32892
rect 27816 32796 28488 32824
rect 28626 32784 28632 32836
rect 28684 32784 28690 32836
rect 28828 32824 28856 32852
rect 31680 32833 31708 32864
rect 31938 32852 31944 32904
rect 31996 32852 32002 32904
rect 32214 32852 32220 32904
rect 32272 32852 32278 32904
rect 32398 32852 32404 32904
rect 32456 32852 32462 32904
rect 32493 32895 32551 32901
rect 32493 32861 32505 32895
rect 32539 32892 32551 32895
rect 33410 32892 33416 32904
rect 32539 32864 33416 32892
rect 32539 32861 32551 32864
rect 32493 32855 32551 32861
rect 33410 32852 33416 32864
rect 33468 32852 33474 32904
rect 28905 32827 28963 32833
rect 28905 32824 28917 32827
rect 28828 32796 28917 32824
rect 28905 32793 28917 32796
rect 28951 32793 28963 32827
rect 28905 32787 28963 32793
rect 31021 32827 31079 32833
rect 31021 32793 31033 32827
rect 31067 32793 31079 32827
rect 31021 32787 31079 32793
rect 31665 32827 31723 32833
rect 31665 32793 31677 32827
rect 31711 32793 31723 32827
rect 31665 32787 31723 32793
rect 31757 32827 31815 32833
rect 31757 32793 31769 32827
rect 31803 32824 31815 32827
rect 32769 32827 32827 32833
rect 32769 32824 32781 32827
rect 31803 32796 32781 32824
rect 31803 32793 31815 32796
rect 31757 32787 31815 32793
rect 32769 32793 32781 32796
rect 32815 32793 32827 32827
rect 32769 32787 32827 32793
rect 25041 32759 25099 32765
rect 25041 32725 25053 32759
rect 25087 32725 25099 32759
rect 25041 32719 25099 32725
rect 25222 32716 25228 32768
rect 25280 32756 25286 32768
rect 26142 32756 26148 32768
rect 25280 32728 26148 32756
rect 25280 32716 25286 32728
rect 26142 32716 26148 32728
rect 26200 32716 26206 32768
rect 27154 32716 27160 32768
rect 27212 32756 27218 32768
rect 27295 32759 27353 32765
rect 27295 32756 27307 32759
rect 27212 32728 27307 32756
rect 27212 32716 27218 32728
rect 27295 32725 27307 32728
rect 27341 32725 27353 32759
rect 27295 32719 27353 32725
rect 30374 32716 30380 32768
rect 30432 32756 30438 32768
rect 31036 32756 31064 32787
rect 30432 32728 31064 32756
rect 30432 32716 30438 32728
rect 31110 32716 31116 32768
rect 31168 32756 31174 32768
rect 31772 32756 31800 32787
rect 31168 32728 31800 32756
rect 31168 32716 31174 32728
rect 1104 32666 36432 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 36432 32666
rect 1104 32592 36432 32614
rect 4614 32552 4620 32564
rect 3988 32524 4620 32552
rect 1302 32444 1308 32496
rect 1360 32484 1366 32496
rect 1489 32487 1547 32493
rect 1489 32484 1501 32487
rect 1360 32456 1501 32484
rect 1360 32444 1366 32456
rect 1489 32453 1501 32456
rect 1535 32453 1547 32487
rect 3988 32484 4016 32524
rect 4614 32512 4620 32524
rect 4672 32512 4678 32564
rect 4893 32555 4951 32561
rect 4893 32521 4905 32555
rect 4939 32552 4951 32555
rect 5258 32552 5264 32564
rect 4939 32524 5264 32552
rect 4939 32521 4951 32524
rect 4893 32515 4951 32521
rect 5258 32512 5264 32524
rect 5316 32512 5322 32564
rect 5997 32555 6055 32561
rect 5997 32521 6009 32555
rect 6043 32552 6055 32555
rect 6086 32552 6092 32564
rect 6043 32524 6092 32552
rect 6043 32521 6055 32524
rect 5997 32515 6055 32521
rect 6086 32512 6092 32524
rect 6144 32512 6150 32564
rect 6730 32512 6736 32564
rect 6788 32512 6794 32564
rect 6825 32555 6883 32561
rect 6825 32521 6837 32555
rect 6871 32552 6883 32555
rect 6914 32552 6920 32564
rect 6871 32524 6920 32552
rect 6871 32521 6883 32524
rect 6825 32515 6883 32521
rect 6914 32512 6920 32524
rect 6972 32552 6978 32564
rect 6972 32524 8064 32552
rect 6972 32512 6978 32524
rect 2806 32456 4016 32484
rect 1489 32447 1547 32453
rect 4430 32444 4436 32496
rect 4488 32484 4494 32496
rect 4488 32456 5856 32484
rect 4488 32444 4494 32456
rect 3513 32419 3571 32425
rect 3513 32385 3525 32419
rect 3559 32416 3571 32419
rect 4706 32416 4712 32428
rect 3559 32388 4712 32416
rect 3559 32385 3571 32388
rect 3513 32379 3571 32385
rect 4706 32376 4712 32388
rect 4764 32376 4770 32428
rect 4798 32376 4804 32428
rect 4856 32376 4862 32428
rect 4985 32419 5043 32425
rect 4985 32385 4997 32419
rect 5031 32416 5043 32419
rect 5258 32416 5264 32428
rect 5031 32388 5264 32416
rect 5031 32385 5043 32388
rect 4985 32379 5043 32385
rect 2498 32308 2504 32360
rect 2556 32348 2562 32360
rect 3237 32351 3295 32357
rect 3237 32348 3249 32351
rect 2556 32320 3249 32348
rect 2556 32308 2562 32320
rect 3237 32317 3249 32320
rect 3283 32317 3295 32351
rect 3237 32311 3295 32317
rect 4614 32308 4620 32360
rect 4672 32348 4678 32360
rect 5000 32348 5028 32379
rect 5258 32376 5264 32388
rect 5316 32376 5322 32428
rect 5442 32376 5448 32428
rect 5500 32416 5506 32428
rect 5629 32419 5687 32425
rect 5629 32416 5641 32419
rect 5500 32388 5641 32416
rect 5500 32376 5506 32388
rect 5629 32385 5641 32388
rect 5675 32385 5687 32419
rect 5828 32416 5856 32456
rect 6454 32444 6460 32496
rect 6512 32484 6518 32496
rect 6549 32487 6607 32493
rect 6549 32484 6561 32487
rect 6512 32456 6561 32484
rect 6512 32444 6518 32456
rect 6549 32453 6561 32456
rect 6595 32453 6607 32487
rect 6549 32447 6607 32453
rect 7377 32487 7435 32493
rect 7377 32453 7389 32487
rect 7423 32484 7435 32487
rect 7423 32456 7880 32484
rect 7423 32453 7435 32456
rect 7377 32447 7435 32453
rect 6365 32419 6423 32425
rect 6365 32416 6377 32419
rect 5828 32388 6377 32416
rect 5629 32379 5687 32385
rect 6365 32385 6377 32388
rect 6411 32385 6423 32419
rect 7009 32419 7067 32425
rect 7009 32416 7021 32419
rect 6365 32379 6423 32385
rect 6472 32388 7021 32416
rect 4672 32320 5028 32348
rect 5537 32351 5595 32357
rect 4672 32308 4678 32320
rect 5537 32317 5549 32351
rect 5583 32317 5595 32351
rect 5537 32311 5595 32317
rect 4522 32240 4528 32292
rect 4580 32280 4586 32292
rect 4890 32280 4896 32292
rect 4580 32252 4896 32280
rect 4580 32240 4586 32252
rect 4890 32240 4896 32252
rect 4948 32240 4954 32292
rect 5552 32280 5580 32311
rect 5718 32308 5724 32360
rect 5776 32308 5782 32360
rect 6178 32308 6184 32360
rect 6236 32348 6242 32360
rect 6472 32348 6500 32388
rect 7009 32385 7021 32388
rect 7055 32416 7067 32419
rect 7098 32416 7104 32428
rect 7055 32388 7104 32416
rect 7055 32385 7067 32388
rect 7009 32379 7067 32385
rect 7098 32376 7104 32388
rect 7156 32376 7162 32428
rect 7285 32419 7343 32425
rect 7285 32416 7297 32419
rect 7208 32388 7297 32416
rect 6236 32320 6500 32348
rect 6236 32308 6242 32320
rect 6546 32308 6552 32360
rect 6604 32348 6610 32360
rect 7208 32357 7236 32388
rect 7285 32385 7297 32388
rect 7331 32385 7343 32419
rect 7285 32379 7343 32385
rect 7466 32376 7472 32428
rect 7524 32376 7530 32428
rect 7558 32376 7564 32428
rect 7616 32376 7622 32428
rect 7852 32425 7880 32456
rect 8036 32425 8064 32524
rect 9858 32512 9864 32564
rect 9916 32552 9922 32564
rect 9916 32524 11008 32552
rect 9916 32512 9922 32524
rect 9030 32444 9036 32496
rect 9088 32444 9094 32496
rect 10594 32484 10600 32496
rect 10258 32456 10600 32484
rect 10594 32444 10600 32456
rect 10652 32444 10658 32496
rect 10980 32493 11008 32524
rect 12894 32512 12900 32564
rect 12952 32552 12958 32564
rect 16758 32552 16764 32564
rect 12952 32524 16764 32552
rect 12952 32512 12958 32524
rect 16758 32512 16764 32524
rect 16816 32512 16822 32564
rect 18233 32555 18291 32561
rect 18233 32552 18245 32555
rect 17604 32524 18245 32552
rect 10965 32487 11023 32493
rect 10965 32453 10977 32487
rect 11011 32484 11023 32487
rect 13906 32484 13912 32496
rect 11011 32456 13912 32484
rect 11011 32453 11023 32456
rect 10965 32447 11023 32453
rect 13906 32444 13912 32456
rect 13964 32444 13970 32496
rect 16301 32487 16359 32493
rect 15580 32456 16252 32484
rect 7745 32419 7803 32425
rect 7745 32385 7757 32419
rect 7791 32385 7803 32419
rect 7745 32379 7803 32385
rect 7837 32419 7895 32425
rect 7837 32385 7849 32419
rect 7883 32385 7895 32419
rect 7837 32379 7895 32385
rect 8021 32419 8079 32425
rect 8021 32385 8033 32419
rect 8067 32385 8079 32419
rect 8021 32379 8079 32385
rect 7193 32351 7251 32357
rect 7193 32348 7205 32351
rect 6604 32320 7205 32348
rect 6604 32308 6610 32320
rect 7193 32317 7205 32320
rect 7239 32317 7251 32351
rect 7193 32311 7251 32317
rect 7760 32348 7788 32379
rect 8294 32376 8300 32428
rect 8352 32416 8358 32428
rect 8757 32419 8815 32425
rect 8757 32416 8769 32419
rect 8352 32388 8769 32416
rect 8352 32376 8358 32388
rect 8757 32385 8769 32388
rect 8803 32385 8815 32419
rect 8757 32379 8815 32385
rect 11790 32376 11796 32428
rect 11848 32376 11854 32428
rect 12437 32419 12495 32425
rect 12437 32385 12449 32419
rect 12483 32416 12495 32419
rect 14642 32416 14648 32428
rect 12483 32388 14648 32416
rect 12483 32385 12495 32388
rect 12437 32379 12495 32385
rect 14642 32376 14648 32388
rect 14700 32376 14706 32428
rect 15580 32425 15608 32456
rect 16224 32428 16252 32456
rect 16301 32453 16313 32487
rect 16347 32484 16359 32487
rect 16574 32484 16580 32496
rect 16347 32456 16580 32484
rect 16347 32453 16359 32456
rect 16301 32447 16359 32453
rect 16574 32444 16580 32456
rect 16632 32484 16638 32496
rect 17494 32484 17500 32496
rect 16632 32456 17500 32484
rect 16632 32444 16638 32456
rect 17494 32444 17500 32456
rect 17552 32444 17558 32496
rect 15565 32419 15623 32425
rect 15565 32385 15577 32419
rect 15611 32385 15623 32419
rect 15565 32379 15623 32385
rect 15838 32376 15844 32428
rect 15896 32376 15902 32428
rect 16117 32419 16175 32425
rect 16117 32385 16129 32419
rect 16163 32385 16175 32419
rect 16117 32379 16175 32385
rect 8478 32348 8484 32360
rect 7760 32320 8484 32348
rect 6086 32280 6092 32292
rect 5552 32252 6092 32280
rect 2590 32172 2596 32224
rect 2648 32212 2654 32224
rect 4982 32212 4988 32224
rect 2648 32184 4988 32212
rect 2648 32172 2654 32184
rect 4982 32172 4988 32184
rect 5040 32172 5046 32224
rect 5074 32172 5080 32224
rect 5132 32172 5138 32224
rect 5442 32172 5448 32224
rect 5500 32172 5506 32224
rect 5828 32221 5856 32252
rect 6086 32240 6092 32252
rect 6144 32240 6150 32292
rect 7466 32240 7472 32292
rect 7524 32280 7530 32292
rect 7760 32280 7788 32320
rect 8478 32308 8484 32320
rect 8536 32348 8542 32360
rect 9490 32348 9496 32360
rect 8536 32320 9496 32348
rect 8536 32308 8542 32320
rect 9490 32308 9496 32320
rect 9548 32308 9554 32360
rect 9582 32308 9588 32360
rect 9640 32348 9646 32360
rect 10318 32348 10324 32360
rect 9640 32320 10324 32348
rect 9640 32308 9646 32320
rect 10318 32308 10324 32320
rect 10376 32308 10382 32360
rect 12069 32351 12127 32357
rect 12069 32317 12081 32351
rect 12115 32348 12127 32351
rect 12342 32348 12348 32360
rect 12115 32320 12348 32348
rect 12115 32317 12127 32320
rect 12069 32311 12127 32317
rect 12342 32308 12348 32320
rect 12400 32308 12406 32360
rect 13906 32308 13912 32360
rect 13964 32348 13970 32360
rect 14918 32348 14924 32360
rect 13964 32320 14924 32348
rect 13964 32308 13970 32320
rect 14918 32308 14924 32320
rect 14976 32308 14982 32360
rect 16132 32348 16160 32379
rect 16206 32376 16212 32428
rect 16264 32376 16270 32428
rect 16390 32376 16396 32428
rect 16448 32416 16454 32428
rect 16485 32419 16543 32425
rect 16485 32416 16497 32419
rect 16448 32388 16497 32416
rect 16448 32376 16454 32388
rect 16485 32385 16497 32388
rect 16531 32385 16543 32419
rect 16485 32379 16543 32385
rect 17604 32348 17632 32524
rect 18233 32521 18245 32524
rect 18279 32552 18291 32555
rect 18874 32552 18880 32564
rect 18279 32524 18880 32552
rect 18279 32521 18291 32524
rect 18233 32515 18291 32521
rect 18874 32512 18880 32524
rect 18932 32512 18938 32564
rect 19705 32555 19763 32561
rect 19705 32552 19717 32555
rect 18984 32524 19717 32552
rect 18322 32484 18328 32496
rect 17788 32456 18328 32484
rect 17788 32425 17816 32456
rect 18322 32444 18328 32456
rect 18380 32444 18386 32496
rect 17773 32419 17831 32425
rect 17773 32385 17785 32419
rect 17819 32385 17831 32419
rect 17773 32379 17831 32385
rect 18046 32376 18052 32428
rect 18104 32416 18110 32428
rect 18141 32419 18199 32425
rect 18141 32416 18153 32419
rect 18104 32388 18153 32416
rect 18104 32376 18110 32388
rect 18141 32385 18153 32388
rect 18187 32385 18199 32419
rect 18141 32379 18199 32385
rect 16132 32320 17632 32348
rect 17678 32308 17684 32360
rect 17736 32308 17742 32360
rect 17865 32351 17923 32357
rect 17865 32317 17877 32351
rect 17911 32317 17923 32351
rect 17865 32311 17923 32317
rect 7524 32252 7788 32280
rect 7524 32240 7530 32252
rect 7926 32240 7932 32292
rect 7984 32280 7990 32292
rect 8386 32280 8392 32292
rect 7984 32252 8392 32280
rect 7984 32240 7990 32252
rect 8386 32240 8392 32252
rect 8444 32240 8450 32292
rect 11238 32240 11244 32292
rect 11296 32280 11302 32292
rect 12253 32283 12311 32289
rect 12253 32280 12265 32283
rect 11296 32252 12265 32280
rect 11296 32240 11302 32252
rect 12253 32249 12265 32252
rect 12299 32249 12311 32283
rect 12253 32243 12311 32249
rect 15749 32283 15807 32289
rect 15749 32249 15761 32283
rect 15795 32280 15807 32283
rect 16114 32280 16120 32292
rect 15795 32252 16120 32280
rect 15795 32249 15807 32252
rect 15749 32243 15807 32249
rect 16114 32240 16120 32252
rect 16172 32240 16178 32292
rect 17880 32280 17908 32311
rect 17954 32308 17960 32360
rect 18012 32308 18018 32360
rect 18156 32348 18184 32379
rect 18414 32376 18420 32428
rect 18472 32376 18478 32428
rect 18984 32425 19012 32524
rect 19705 32521 19717 32524
rect 19751 32552 19763 32555
rect 19794 32552 19800 32564
rect 19751 32524 19800 32552
rect 19751 32521 19763 32524
rect 19705 32515 19763 32521
rect 19794 32512 19800 32524
rect 19852 32512 19858 32564
rect 19886 32512 19892 32564
rect 19944 32512 19950 32564
rect 21545 32555 21603 32561
rect 21545 32521 21557 32555
rect 21591 32552 21603 32555
rect 21634 32552 21640 32564
rect 21591 32524 21640 32552
rect 21591 32521 21603 32524
rect 21545 32515 21603 32521
rect 21634 32512 21640 32524
rect 21692 32512 21698 32564
rect 21726 32512 21732 32564
rect 21784 32552 21790 32564
rect 21784 32524 21956 32552
rect 21784 32512 21790 32524
rect 21266 32484 21272 32496
rect 19076 32456 21272 32484
rect 18969 32419 19027 32425
rect 18969 32385 18981 32419
rect 19015 32385 19027 32419
rect 18969 32379 19027 32385
rect 19076 32348 19104 32456
rect 19153 32419 19211 32425
rect 19153 32385 19165 32419
rect 19199 32385 19211 32419
rect 19153 32379 19211 32385
rect 18156 32320 19104 32348
rect 18417 32283 18475 32289
rect 18417 32280 18429 32283
rect 17880 32252 18429 32280
rect 18417 32249 18429 32252
rect 18463 32280 18475 32283
rect 19168 32280 19196 32379
rect 19242 32376 19248 32428
rect 19300 32376 19306 32428
rect 19334 32376 19340 32428
rect 19392 32376 19398 32428
rect 19426 32376 19432 32428
rect 19484 32376 19490 32428
rect 19845 32425 19873 32456
rect 21266 32444 21272 32456
rect 21324 32484 21330 32496
rect 21928 32484 21956 32524
rect 22002 32512 22008 32564
rect 22060 32552 22066 32564
rect 22060 32524 22692 32552
rect 22060 32512 22066 32524
rect 22097 32487 22155 32493
rect 22097 32484 22109 32487
rect 21324 32456 21772 32484
rect 21928 32456 22109 32484
rect 21324 32444 21330 32456
rect 19830 32419 19888 32425
rect 19830 32385 19842 32419
rect 19876 32385 19888 32419
rect 19830 32379 19888 32385
rect 19978 32376 19984 32428
rect 20036 32416 20042 32428
rect 20349 32419 20407 32425
rect 20349 32416 20361 32419
rect 20036 32388 20361 32416
rect 20036 32376 20042 32388
rect 20349 32385 20361 32388
rect 20395 32385 20407 32419
rect 20349 32379 20407 32385
rect 21453 32419 21511 32425
rect 21453 32385 21465 32419
rect 21499 32385 21511 32419
rect 21453 32379 21511 32385
rect 21468 32348 21496 32379
rect 21634 32376 21640 32428
rect 21692 32376 21698 32428
rect 19352 32320 21496 32348
rect 21744 32348 21772 32456
rect 22097 32453 22109 32456
rect 22143 32453 22155 32487
rect 22097 32447 22155 32453
rect 22189 32487 22247 32493
rect 22189 32453 22201 32487
rect 22235 32484 22247 32487
rect 22554 32484 22560 32496
rect 22235 32456 22560 32484
rect 22235 32453 22247 32456
rect 22189 32447 22247 32453
rect 22554 32444 22560 32456
rect 22612 32444 22618 32496
rect 22664 32484 22692 32524
rect 22738 32512 22744 32564
rect 22796 32512 22802 32564
rect 22922 32512 22928 32564
rect 22980 32552 22986 32564
rect 22980 32524 23060 32552
rect 22980 32512 22986 32524
rect 22664 32456 22876 32484
rect 22848 32428 22876 32456
rect 21818 32376 21824 32428
rect 21876 32376 21882 32428
rect 21910 32376 21916 32428
rect 21968 32416 21974 32428
rect 22286 32419 22344 32425
rect 22286 32416 22298 32419
rect 21968 32388 22013 32416
rect 22066 32388 22298 32416
rect 21968 32376 21974 32388
rect 22066 32348 22094 32388
rect 22286 32385 22298 32388
rect 22332 32385 22344 32419
rect 22286 32379 22344 32385
rect 22830 32376 22836 32428
rect 22888 32416 22894 32428
rect 23032 32425 23060 32524
rect 23474 32512 23480 32564
rect 23532 32512 23538 32564
rect 24118 32512 24124 32564
rect 24176 32552 24182 32564
rect 25314 32552 25320 32564
rect 24176 32524 25320 32552
rect 24176 32512 24182 32524
rect 25314 32512 25320 32524
rect 25372 32512 25378 32564
rect 25409 32555 25467 32561
rect 25409 32521 25421 32555
rect 25455 32552 25467 32555
rect 26050 32552 26056 32564
rect 25455 32524 26056 32552
rect 25455 32521 25467 32524
rect 25409 32515 25467 32521
rect 26050 32512 26056 32524
rect 26108 32512 26114 32564
rect 26234 32512 26240 32564
rect 26292 32552 26298 32564
rect 26510 32552 26516 32564
rect 26292 32524 26516 32552
rect 26292 32512 26298 32524
rect 26510 32512 26516 32524
rect 26568 32512 26574 32564
rect 27617 32555 27675 32561
rect 27617 32521 27629 32555
rect 27663 32552 27675 32555
rect 27985 32555 28043 32561
rect 27985 32552 27997 32555
rect 27663 32524 27997 32552
rect 27663 32521 27675 32524
rect 27617 32515 27675 32521
rect 27985 32521 27997 32524
rect 28031 32552 28043 32555
rect 28074 32552 28080 32564
rect 28031 32524 28080 32552
rect 28031 32521 28043 32524
rect 27985 32515 28043 32521
rect 28074 32512 28080 32524
rect 28132 32512 28138 32564
rect 29178 32512 29184 32564
rect 29236 32512 29242 32564
rect 29365 32555 29423 32561
rect 29365 32521 29377 32555
rect 29411 32552 29423 32555
rect 30282 32552 30288 32564
rect 29411 32524 30288 32552
rect 29411 32521 29423 32524
rect 29365 32515 29423 32521
rect 30282 32512 30288 32524
rect 30340 32512 30346 32564
rect 30374 32512 30380 32564
rect 30432 32512 30438 32564
rect 30742 32512 30748 32564
rect 30800 32512 30806 32564
rect 31205 32555 31263 32561
rect 31205 32521 31217 32555
rect 31251 32552 31263 32555
rect 31294 32552 31300 32564
rect 31251 32524 31300 32552
rect 31251 32521 31263 32524
rect 31205 32515 31263 32521
rect 31294 32512 31300 32524
rect 31352 32512 31358 32564
rect 31573 32555 31631 32561
rect 31573 32552 31585 32555
rect 31496 32524 31585 32552
rect 23198 32444 23204 32496
rect 23256 32493 23262 32496
rect 23256 32487 23305 32493
rect 23256 32453 23259 32487
rect 23293 32484 23305 32487
rect 24136 32484 24164 32512
rect 23293 32456 24164 32484
rect 24765 32487 24823 32493
rect 23293 32453 23305 32456
rect 23256 32447 23305 32453
rect 24765 32453 24777 32487
rect 24811 32484 24823 32487
rect 24854 32484 24860 32496
rect 24811 32456 24860 32484
rect 24811 32453 24823 32456
rect 24765 32447 24823 32453
rect 23256 32444 23262 32447
rect 24854 32444 24860 32456
rect 24912 32444 24918 32496
rect 26418 32484 26424 32496
rect 25240 32456 26424 32484
rect 22925 32419 22983 32425
rect 22925 32416 22937 32419
rect 22888 32388 22937 32416
rect 22888 32376 22894 32388
rect 22925 32385 22937 32388
rect 22971 32385 22983 32419
rect 22925 32379 22983 32385
rect 23017 32419 23075 32425
rect 23017 32385 23029 32419
rect 23063 32385 23075 32419
rect 23017 32379 23075 32385
rect 23109 32419 23167 32425
rect 23109 32385 23121 32419
rect 23155 32385 23167 32419
rect 23109 32379 23167 32385
rect 23124 32348 23152 32379
rect 23382 32376 23388 32428
rect 23440 32376 23446 32428
rect 23750 32376 23756 32428
rect 23808 32416 23814 32428
rect 24213 32419 24271 32425
rect 24213 32416 24225 32419
rect 23808 32388 24225 32416
rect 23808 32376 23814 32388
rect 24213 32385 24225 32388
rect 24259 32385 24271 32419
rect 24213 32379 24271 32385
rect 24302 32376 24308 32428
rect 24360 32416 24366 32428
rect 25240 32425 25268 32456
rect 26418 32444 26424 32456
rect 26476 32444 26482 32496
rect 27341 32487 27399 32493
rect 27341 32453 27353 32487
rect 27387 32484 27399 32487
rect 27522 32484 27528 32496
rect 27387 32456 27528 32484
rect 27387 32453 27399 32456
rect 27341 32447 27399 32453
rect 27522 32444 27528 32456
rect 27580 32444 27586 32496
rect 27706 32444 27712 32496
rect 27764 32484 27770 32496
rect 27764 32456 28120 32484
rect 27764 32444 27770 32456
rect 24397 32419 24455 32425
rect 24397 32416 24409 32419
rect 24360 32388 24409 32416
rect 24360 32376 24366 32388
rect 24397 32385 24409 32388
rect 24443 32385 24455 32419
rect 24397 32379 24455 32385
rect 25225 32419 25283 32425
rect 26602 32422 26608 32428
rect 25225 32385 25237 32419
rect 25271 32385 25283 32419
rect 26528 32416 26608 32422
rect 25225 32379 25283 32385
rect 26068 32394 26608 32416
rect 26068 32388 26556 32394
rect 23474 32348 23480 32360
rect 21744 32320 22094 32348
rect 23032 32320 23480 32348
rect 19352 32292 19380 32320
rect 18463 32252 19196 32280
rect 18463 32249 18475 32252
rect 18417 32243 18475 32249
rect 19334 32240 19340 32292
rect 19392 32240 19398 32292
rect 19613 32283 19671 32289
rect 19613 32249 19625 32283
rect 19659 32280 19671 32283
rect 19886 32280 19892 32292
rect 19659 32252 19892 32280
rect 19659 32249 19671 32252
rect 19613 32243 19671 32249
rect 19886 32240 19892 32252
rect 19944 32240 19950 32292
rect 21468 32280 21496 32320
rect 23032 32280 23060 32320
rect 23474 32308 23480 32320
rect 23532 32308 23538 32360
rect 24026 32308 24032 32360
rect 24084 32308 24090 32360
rect 25133 32351 25191 32357
rect 25133 32317 25145 32351
rect 25179 32348 25191 32351
rect 26068 32348 26096 32388
rect 26602 32376 26608 32394
rect 26660 32376 26666 32428
rect 27249 32419 27307 32425
rect 27249 32385 27261 32419
rect 27295 32416 27307 32419
rect 27982 32416 27988 32428
rect 27295 32388 27988 32416
rect 27295 32385 27307 32388
rect 27249 32379 27307 32385
rect 27982 32376 27988 32388
rect 28040 32376 28046 32428
rect 28092 32416 28120 32456
rect 28166 32444 28172 32496
rect 28224 32444 28230 32496
rect 29196 32484 29224 32512
rect 29914 32484 29920 32496
rect 29196 32456 29920 32484
rect 29914 32444 29920 32456
rect 29972 32444 29978 32496
rect 30006 32444 30012 32496
rect 30064 32444 30070 32496
rect 31018 32484 31024 32496
rect 30392 32456 31024 32484
rect 28445 32419 28503 32425
rect 28445 32416 28457 32419
rect 28092 32388 28457 32416
rect 28445 32385 28457 32388
rect 28491 32416 28503 32419
rect 29086 32416 29092 32428
rect 28491 32388 29092 32416
rect 28491 32385 28503 32388
rect 28445 32379 28503 32385
rect 29086 32376 29092 32388
rect 29144 32376 29150 32428
rect 29181 32419 29239 32425
rect 29181 32385 29193 32419
rect 29227 32385 29239 32419
rect 29181 32379 29239 32385
rect 25179 32320 26096 32348
rect 26145 32351 26203 32357
rect 25179 32317 25191 32320
rect 25133 32311 25191 32317
rect 26145 32317 26157 32351
rect 26191 32348 26203 32351
rect 26234 32348 26240 32360
rect 26191 32320 26240 32348
rect 26191 32317 26203 32320
rect 26145 32311 26203 32317
rect 26160 32280 26188 32311
rect 26234 32308 26240 32320
rect 26292 32308 26298 32360
rect 26329 32351 26387 32357
rect 26329 32317 26341 32351
rect 26375 32317 26387 32351
rect 26329 32311 26387 32317
rect 21468 32252 23060 32280
rect 25240 32252 26188 32280
rect 5813 32215 5871 32221
rect 5813 32181 5825 32215
rect 5859 32181 5871 32215
rect 5813 32175 5871 32181
rect 7374 32172 7380 32224
rect 7432 32212 7438 32224
rect 7561 32215 7619 32221
rect 7561 32212 7573 32215
rect 7432 32184 7573 32212
rect 7432 32172 7438 32184
rect 7561 32181 7573 32184
rect 7607 32181 7619 32215
rect 7561 32175 7619 32181
rect 7650 32172 7656 32224
rect 7708 32212 7714 32224
rect 7837 32215 7895 32221
rect 7837 32212 7849 32215
rect 7708 32184 7849 32212
rect 7708 32172 7714 32184
rect 7837 32181 7849 32184
rect 7883 32181 7895 32215
rect 7837 32175 7895 32181
rect 8846 32172 8852 32224
rect 8904 32212 8910 32224
rect 10505 32215 10563 32221
rect 10505 32212 10517 32215
rect 8904 32184 10517 32212
rect 8904 32172 8910 32184
rect 10505 32181 10517 32184
rect 10551 32181 10563 32215
rect 10505 32175 10563 32181
rect 11422 32172 11428 32224
rect 11480 32212 11486 32224
rect 11609 32215 11667 32221
rect 11609 32212 11621 32215
rect 11480 32184 11621 32212
rect 11480 32172 11486 32184
rect 11609 32181 11621 32184
rect 11655 32181 11667 32215
rect 11609 32175 11667 32181
rect 11882 32172 11888 32224
rect 11940 32212 11946 32224
rect 11977 32215 12035 32221
rect 11977 32212 11989 32215
rect 11940 32184 11989 32212
rect 11940 32172 11946 32184
rect 11977 32181 11989 32184
rect 12023 32181 12035 32215
rect 11977 32175 12035 32181
rect 15381 32215 15439 32221
rect 15381 32181 15393 32215
rect 15427 32212 15439 32215
rect 15470 32212 15476 32224
rect 15427 32184 15476 32212
rect 15427 32181 15439 32184
rect 15381 32175 15439 32181
rect 15470 32172 15476 32184
rect 15528 32172 15534 32224
rect 15930 32172 15936 32224
rect 15988 32172 15994 32224
rect 17494 32172 17500 32224
rect 17552 32172 17558 32224
rect 20257 32215 20315 32221
rect 20257 32181 20269 32215
rect 20303 32212 20315 32215
rect 20438 32212 20444 32224
rect 20303 32184 20444 32212
rect 20303 32181 20315 32184
rect 20257 32175 20315 32181
rect 20438 32172 20444 32184
rect 20496 32172 20502 32224
rect 22465 32215 22523 32221
rect 22465 32181 22477 32215
rect 22511 32212 22523 32215
rect 23106 32212 23112 32224
rect 22511 32184 23112 32212
rect 22511 32181 22523 32184
rect 22465 32175 22523 32181
rect 23106 32172 23112 32184
rect 23164 32172 23170 32224
rect 24302 32172 24308 32224
rect 24360 32212 24366 32224
rect 24581 32215 24639 32221
rect 24581 32212 24593 32215
rect 24360 32184 24593 32212
rect 24360 32172 24366 32184
rect 24581 32181 24593 32184
rect 24627 32212 24639 32215
rect 25130 32212 25136 32224
rect 24627 32184 25136 32212
rect 24627 32181 24639 32184
rect 24581 32175 24639 32181
rect 25130 32172 25136 32184
rect 25188 32172 25194 32224
rect 25240 32221 25268 32252
rect 25225 32215 25283 32221
rect 25225 32181 25237 32215
rect 25271 32181 25283 32215
rect 25225 32175 25283 32181
rect 25501 32215 25559 32221
rect 25501 32181 25513 32215
rect 25547 32212 25559 32215
rect 25682 32212 25688 32224
rect 25547 32184 25688 32212
rect 25547 32181 25559 32184
rect 25501 32175 25559 32181
rect 25682 32172 25688 32184
rect 25740 32172 25746 32224
rect 26142 32172 26148 32224
rect 26200 32212 26206 32224
rect 26344 32212 26372 32311
rect 26418 32308 26424 32360
rect 26476 32308 26482 32360
rect 26510 32308 26516 32360
rect 26568 32308 26574 32360
rect 26970 32308 26976 32360
rect 27028 32308 27034 32360
rect 27458 32351 27516 32357
rect 27458 32317 27470 32351
rect 27504 32348 27516 32351
rect 27706 32348 27712 32360
rect 27504 32320 27712 32348
rect 27504 32317 27516 32320
rect 27458 32311 27516 32317
rect 27706 32308 27712 32320
rect 27764 32308 27770 32360
rect 28350 32308 28356 32360
rect 28408 32348 28414 32360
rect 28721 32351 28779 32357
rect 28721 32348 28733 32351
rect 28408 32320 28733 32348
rect 28408 32308 28414 32320
rect 28721 32317 28733 32320
rect 28767 32317 28779 32351
rect 29196 32348 29224 32379
rect 29270 32376 29276 32428
rect 29328 32376 29334 32428
rect 29638 32376 29644 32428
rect 29696 32376 29702 32428
rect 29822 32425 29828 32428
rect 29789 32419 29828 32425
rect 29789 32385 29801 32419
rect 29789 32379 29828 32385
rect 29822 32376 29828 32379
rect 29880 32376 29886 32428
rect 30190 32425 30196 32428
rect 30147 32419 30196 32425
rect 30147 32385 30159 32419
rect 30193 32385 30196 32419
rect 30147 32379 30196 32385
rect 30190 32376 30196 32379
rect 30248 32376 30254 32428
rect 29454 32348 29460 32360
rect 29196 32320 29460 32348
rect 28721 32311 28779 32317
rect 29454 32308 29460 32320
rect 29512 32308 29518 32360
rect 30392 32348 30420 32456
rect 31018 32444 31024 32456
rect 31076 32484 31082 32496
rect 31389 32487 31447 32493
rect 31389 32484 31401 32487
rect 31076 32456 31401 32484
rect 31076 32444 31082 32456
rect 31389 32453 31401 32456
rect 31435 32453 31447 32487
rect 31389 32447 31447 32453
rect 30466 32376 30472 32428
rect 30524 32416 30530 32428
rect 31113 32419 31171 32425
rect 30524 32388 31064 32416
rect 30524 32376 30530 32388
rect 29748 32320 30420 32348
rect 30561 32351 30619 32357
rect 29748 32292 29776 32320
rect 30561 32317 30573 32351
rect 30607 32317 30619 32351
rect 30561 32311 30619 32317
rect 28261 32283 28319 32289
rect 28261 32280 28273 32283
rect 26436 32252 28273 32280
rect 26436 32224 26464 32252
rect 28261 32249 28273 32252
rect 28307 32249 28319 32283
rect 28261 32243 28319 32249
rect 28997 32283 29055 32289
rect 28997 32249 29009 32283
rect 29043 32280 29055 32283
rect 29730 32280 29736 32292
rect 29043 32252 29736 32280
rect 29043 32249 29055 32252
rect 28997 32243 29055 32249
rect 29730 32240 29736 32252
rect 29788 32240 29794 32292
rect 30285 32283 30343 32289
rect 30285 32249 30297 32283
rect 30331 32280 30343 32283
rect 30576 32280 30604 32311
rect 30650 32308 30656 32360
rect 30708 32308 30714 32360
rect 30926 32308 30932 32360
rect 30984 32308 30990 32360
rect 31036 32357 31064 32388
rect 31113 32385 31125 32419
rect 31159 32385 31171 32419
rect 31113 32379 31171 32385
rect 31021 32351 31079 32357
rect 31021 32317 31033 32351
rect 31067 32317 31079 32351
rect 31128 32348 31156 32379
rect 31294 32376 31300 32428
rect 31352 32376 31358 32428
rect 31496 32416 31524 32524
rect 31573 32521 31585 32524
rect 31619 32521 31631 32555
rect 31573 32515 31631 32521
rect 31757 32555 31815 32561
rect 31757 32521 31769 32555
rect 31803 32552 31815 32555
rect 32214 32552 32220 32564
rect 31803 32524 32220 32552
rect 31803 32521 31815 32524
rect 31757 32515 31815 32521
rect 32214 32512 32220 32524
rect 32272 32512 32278 32564
rect 33410 32512 33416 32564
rect 33468 32512 33474 32564
rect 31846 32444 31852 32496
rect 31904 32484 31910 32496
rect 32447 32487 32505 32493
rect 32447 32484 32459 32487
rect 31904 32456 32459 32484
rect 31904 32444 31910 32456
rect 32447 32453 32459 32456
rect 32493 32453 32505 32487
rect 32447 32447 32505 32453
rect 32674 32444 32680 32496
rect 32732 32444 32738 32496
rect 31570 32416 31576 32428
rect 31496 32388 31576 32416
rect 31570 32376 31576 32388
rect 31628 32376 31634 32428
rect 31665 32419 31723 32425
rect 31665 32385 31677 32419
rect 31711 32385 31723 32419
rect 31665 32379 31723 32385
rect 31478 32348 31484 32360
rect 31128 32320 31484 32348
rect 31021 32311 31079 32317
rect 31478 32308 31484 32320
rect 31536 32308 31542 32360
rect 30331 32252 30604 32280
rect 30331 32249 30343 32252
rect 30285 32243 30343 32249
rect 31570 32240 31576 32292
rect 31628 32280 31634 32292
rect 31680 32280 31708 32379
rect 32582 32376 32588 32428
rect 32640 32376 32646 32428
rect 32766 32376 32772 32428
rect 32824 32376 32830 32428
rect 32953 32419 33011 32425
rect 32953 32385 32965 32419
rect 32999 32416 33011 32419
rect 33045 32419 33103 32425
rect 33045 32416 33057 32419
rect 32999 32388 33057 32416
rect 32999 32385 33011 32388
rect 32953 32379 33011 32385
rect 33045 32385 33057 32388
rect 33091 32385 33103 32419
rect 33045 32379 33103 32385
rect 33229 32419 33287 32425
rect 33229 32385 33241 32419
rect 33275 32385 33287 32419
rect 33229 32379 33287 32385
rect 32306 32308 32312 32360
rect 32364 32308 32370 32360
rect 32122 32280 32128 32292
rect 31628 32252 31708 32280
rect 31772 32252 32128 32280
rect 31628 32240 31634 32252
rect 26200 32184 26372 32212
rect 26200 32172 26206 32184
rect 26418 32172 26424 32224
rect 26476 32172 26482 32224
rect 26786 32172 26792 32224
rect 26844 32172 26850 32224
rect 27798 32172 27804 32224
rect 27856 32172 27862 32224
rect 27985 32215 28043 32221
rect 27985 32181 27997 32215
rect 28031 32212 28043 32215
rect 28166 32212 28172 32224
rect 28031 32184 28172 32212
rect 28031 32181 28043 32184
rect 27985 32175 28043 32181
rect 28166 32172 28172 32184
rect 28224 32172 28230 32224
rect 28626 32172 28632 32224
rect 28684 32172 28690 32224
rect 29454 32172 29460 32224
rect 29512 32212 29518 32224
rect 29549 32215 29607 32221
rect 29549 32212 29561 32215
rect 29512 32184 29561 32212
rect 29512 32172 29518 32184
rect 29549 32181 29561 32184
rect 29595 32212 29607 32215
rect 29638 32212 29644 32224
rect 29595 32184 29644 32212
rect 29595 32181 29607 32184
rect 29549 32175 29607 32181
rect 29638 32172 29644 32184
rect 29696 32172 29702 32224
rect 29914 32172 29920 32224
rect 29972 32212 29978 32224
rect 31772 32212 31800 32252
rect 32122 32240 32128 32252
rect 32180 32240 32186 32292
rect 29972 32184 31800 32212
rect 31941 32215 31999 32221
rect 29972 32172 29978 32184
rect 31941 32181 31953 32215
rect 31987 32212 31999 32215
rect 32858 32212 32864 32224
rect 31987 32184 32864 32212
rect 31987 32181 31999 32184
rect 31941 32175 31999 32181
rect 32858 32172 32864 32184
rect 32916 32212 32922 32224
rect 33244 32212 33272 32379
rect 32916 32184 33272 32212
rect 32916 32172 32922 32184
rect 1104 32122 36432 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 36432 32122
rect 1104 32048 36432 32070
rect 2317 32011 2375 32017
rect 2317 31977 2329 32011
rect 2363 32008 2375 32011
rect 2498 32008 2504 32020
rect 2363 31980 2504 32008
rect 2363 31977 2375 31980
rect 2317 31971 2375 31977
rect 2498 31968 2504 31980
rect 2556 31968 2562 32020
rect 3145 32011 3203 32017
rect 3145 31977 3157 32011
rect 3191 32008 3203 32011
rect 4154 32008 4160 32020
rect 3191 31980 4160 32008
rect 3191 31977 3203 31980
rect 3145 31971 3203 31977
rect 4154 31968 4160 31980
rect 4212 31968 4218 32020
rect 4430 31968 4436 32020
rect 4488 32008 4494 32020
rect 6365 32011 6423 32017
rect 6365 32008 6377 32011
rect 4488 31980 6377 32008
rect 4488 31968 4494 31980
rect 6365 31977 6377 31980
rect 6411 31977 6423 32011
rect 6365 31971 6423 31977
rect 7006 31968 7012 32020
rect 7064 32008 7070 32020
rect 7101 32011 7159 32017
rect 7101 32008 7113 32011
rect 7064 31980 7113 32008
rect 7064 31968 7070 31980
rect 7101 31977 7113 31980
rect 7147 32008 7159 32011
rect 7558 32008 7564 32020
rect 7147 31980 7564 32008
rect 7147 31977 7159 31980
rect 7101 31971 7159 31977
rect 7558 31968 7564 31980
rect 7616 31968 7622 32020
rect 8018 31968 8024 32020
rect 8076 31968 8082 32020
rect 9401 32011 9459 32017
rect 9401 31977 9413 32011
rect 9447 32008 9459 32011
rect 10226 32008 10232 32020
rect 9447 31980 10232 32008
rect 9447 31977 9459 31980
rect 9401 31971 9459 31977
rect 10226 31968 10232 31980
rect 10284 31968 10290 32020
rect 10594 31968 10600 32020
rect 10652 32008 10658 32020
rect 10652 31980 13676 32008
rect 10652 31968 10658 31980
rect 2406 31900 2412 31952
rect 2464 31940 2470 31952
rect 5537 31943 5595 31949
rect 2464 31912 3556 31940
rect 2464 31900 2470 31912
rect 1302 31832 1308 31884
rect 1360 31872 1366 31884
rect 1360 31844 2728 31872
rect 1360 31832 1366 31844
rect 2501 31807 2559 31813
rect 2501 31773 2513 31807
rect 2547 31804 2559 31807
rect 2590 31804 2596 31816
rect 2547 31776 2596 31804
rect 2547 31773 2559 31776
rect 2501 31767 2559 31773
rect 2590 31764 2596 31776
rect 2648 31764 2654 31816
rect 2700 31813 2728 31844
rect 2685 31807 2743 31813
rect 2685 31773 2697 31807
rect 2731 31773 2743 31807
rect 2685 31767 2743 31773
rect 2774 31764 2780 31816
rect 2832 31764 2838 31816
rect 3326 31764 3332 31816
rect 3384 31764 3390 31816
rect 3528 31813 3556 31912
rect 5537 31909 5549 31943
rect 5583 31940 5595 31943
rect 6546 31940 6552 31952
rect 5583 31912 6552 31940
rect 5583 31909 5595 31912
rect 5537 31903 5595 31909
rect 6546 31900 6552 31912
rect 6604 31900 6610 31952
rect 6641 31943 6699 31949
rect 6641 31909 6653 31943
rect 6687 31940 6699 31943
rect 6914 31940 6920 31952
rect 6687 31912 6920 31940
rect 6687 31909 6699 31912
rect 6641 31903 6699 31909
rect 6914 31900 6920 31912
rect 6972 31900 6978 31952
rect 7024 31912 7788 31940
rect 3789 31875 3847 31881
rect 3789 31841 3801 31875
rect 3835 31872 3847 31875
rect 4706 31872 4712 31884
rect 3835 31844 4712 31872
rect 3835 31841 3847 31844
rect 3789 31835 3847 31841
rect 3513 31807 3571 31813
rect 3513 31773 3525 31807
rect 3559 31773 3571 31807
rect 3513 31767 3571 31773
rect 3605 31807 3663 31813
rect 3605 31773 3617 31807
rect 3651 31773 3663 31807
rect 3605 31767 3663 31773
rect 2792 31736 2820 31764
rect 3620 31736 3648 31767
rect 2792 31708 3648 31736
rect 3694 31628 3700 31680
rect 3752 31668 3758 31680
rect 3804 31668 3832 31835
rect 4706 31832 4712 31844
rect 4764 31832 4770 31884
rect 5074 31832 5080 31884
rect 5132 31872 5138 31884
rect 5626 31872 5632 31884
rect 5132 31844 5632 31872
rect 5132 31832 5138 31844
rect 5626 31832 5632 31844
rect 5684 31872 5690 31884
rect 6273 31875 6331 31881
rect 6273 31872 6285 31875
rect 5684 31844 6285 31872
rect 5684 31832 5690 31844
rect 6273 31841 6285 31844
rect 6319 31841 6331 31875
rect 7024 31872 7052 31912
rect 6273 31835 6331 31841
rect 6564 31844 7052 31872
rect 5442 31764 5448 31816
rect 5500 31804 5506 31816
rect 5810 31804 5816 31816
rect 5500 31776 5816 31804
rect 5500 31764 5506 31776
rect 5810 31764 5816 31776
rect 5868 31764 5874 31816
rect 5905 31807 5963 31813
rect 5905 31773 5917 31807
rect 5951 31804 5963 31807
rect 6086 31804 6092 31816
rect 5951 31776 6092 31804
rect 5951 31773 5963 31776
rect 5905 31767 5963 31773
rect 6086 31764 6092 31776
rect 6144 31764 6150 31816
rect 6564 31813 6592 31844
rect 7466 31832 7472 31884
rect 7524 31872 7530 31884
rect 7653 31875 7711 31881
rect 7653 31872 7665 31875
rect 7524 31844 7665 31872
rect 7524 31832 7530 31844
rect 7653 31841 7665 31844
rect 7699 31841 7711 31875
rect 7760 31872 7788 31912
rect 8110 31900 8116 31952
rect 8168 31940 8174 31952
rect 8168 31912 9076 31940
rect 8168 31900 8174 31912
rect 8128 31872 8156 31900
rect 7760 31844 8156 31872
rect 7653 31835 7711 31841
rect 8386 31832 8392 31884
rect 8444 31872 8450 31884
rect 8665 31875 8723 31881
rect 8444 31844 8616 31872
rect 8444 31832 8450 31844
rect 6549 31807 6607 31813
rect 6549 31773 6561 31807
rect 6595 31773 6607 31807
rect 6549 31767 6607 31773
rect 6733 31807 6791 31813
rect 6733 31773 6745 31807
rect 6779 31773 6791 31807
rect 6733 31767 6791 31773
rect 4065 31739 4123 31745
rect 4065 31705 4077 31739
rect 4111 31736 4123 31739
rect 4338 31736 4344 31748
rect 4111 31708 4344 31736
rect 4111 31705 4123 31708
rect 4065 31699 4123 31705
rect 4338 31696 4344 31708
rect 4396 31696 4402 31748
rect 5074 31696 5080 31748
rect 5132 31696 5138 31748
rect 6748 31736 6776 31767
rect 6822 31764 6828 31816
rect 6880 31764 6886 31816
rect 7345 31807 7403 31813
rect 7345 31773 7357 31807
rect 7391 31804 7403 31807
rect 7391 31773 7420 31804
rect 7345 31767 7420 31773
rect 5828 31708 6776 31736
rect 7392 31736 7420 31767
rect 7558 31764 7564 31816
rect 7616 31764 7622 31816
rect 7834 31764 7840 31816
rect 7892 31764 7898 31816
rect 8113 31807 8171 31813
rect 8113 31773 8125 31807
rect 8159 31804 8171 31807
rect 8481 31807 8539 31813
rect 8159 31776 8340 31804
rect 8159 31773 8171 31776
rect 8113 31767 8171 31773
rect 7650 31736 7656 31748
rect 7392 31708 7656 31736
rect 3752 31640 3832 31668
rect 3752 31628 3758 31640
rect 4246 31628 4252 31680
rect 4304 31668 4310 31680
rect 4890 31668 4896 31680
rect 4304 31640 4896 31668
rect 4304 31628 4310 31640
rect 4890 31628 4896 31640
rect 4948 31628 4954 31680
rect 5534 31628 5540 31680
rect 5592 31668 5598 31680
rect 5629 31671 5687 31677
rect 5629 31668 5641 31671
rect 5592 31640 5641 31668
rect 5592 31628 5598 31640
rect 5629 31637 5641 31640
rect 5675 31637 5687 31671
rect 5629 31631 5687 31637
rect 5718 31628 5724 31680
rect 5776 31668 5782 31680
rect 5828 31668 5856 31708
rect 7650 31696 7656 31708
rect 7708 31696 7714 31748
rect 5776 31640 5856 31668
rect 5776 31628 5782 31640
rect 6086 31628 6092 31680
rect 6144 31668 6150 31680
rect 6454 31668 6460 31680
rect 6144 31640 6460 31668
rect 6144 31628 6150 31640
rect 6454 31628 6460 31640
rect 6512 31628 6518 31680
rect 8312 31677 8340 31776
rect 8481 31773 8493 31807
rect 8527 31773 8539 31807
rect 8588 31804 8616 31844
rect 8665 31841 8677 31875
rect 8711 31872 8723 31875
rect 8938 31872 8944 31884
rect 8711 31844 8944 31872
rect 8711 31841 8723 31844
rect 8665 31835 8723 31841
rect 8938 31832 8944 31844
rect 8996 31832 9002 31884
rect 9048 31872 9076 31912
rect 9582 31900 9588 31952
rect 9640 31900 9646 31952
rect 9953 31943 10011 31949
rect 9953 31909 9965 31943
rect 9999 31940 10011 31943
rect 10134 31940 10140 31952
rect 9999 31912 10140 31940
rect 9999 31909 10011 31912
rect 9953 31903 10011 31909
rect 10134 31900 10140 31912
rect 10192 31900 10198 31952
rect 10781 31943 10839 31949
rect 10781 31909 10793 31943
rect 10827 31940 10839 31943
rect 13648 31940 13676 31980
rect 13722 31968 13728 32020
rect 13780 31968 13786 32020
rect 15930 32008 15936 32020
rect 15396 31980 15936 32008
rect 13998 31940 14004 31952
rect 10827 31912 11928 31940
rect 13648 31912 14004 31940
rect 10827 31909 10839 31912
rect 10781 31903 10839 31909
rect 9674 31872 9680 31884
rect 9048 31844 9680 31872
rect 9674 31832 9680 31844
rect 9732 31832 9738 31884
rect 10042 31832 10048 31884
rect 10100 31832 10106 31884
rect 11900 31872 11928 31912
rect 13998 31900 14004 31912
rect 14056 31900 14062 31952
rect 15396 31949 15424 31980
rect 15930 31968 15936 31980
rect 15988 31968 15994 32020
rect 17589 32011 17647 32017
rect 17589 31977 17601 32011
rect 17635 32008 17647 32011
rect 17678 32008 17684 32020
rect 17635 31980 17684 32008
rect 17635 31977 17647 31980
rect 17589 31971 17647 31977
rect 17678 31968 17684 31980
rect 17736 31968 17742 32020
rect 19978 32008 19984 32020
rect 17788 31980 19984 32008
rect 15381 31943 15439 31949
rect 15381 31909 15393 31943
rect 15427 31909 15439 31943
rect 15381 31903 15439 31909
rect 15470 31900 15476 31952
rect 15528 31900 15534 31952
rect 17402 31900 17408 31952
rect 17460 31940 17466 31952
rect 17788 31940 17816 31980
rect 19978 31968 19984 31980
rect 20036 31968 20042 32020
rect 20898 31968 20904 32020
rect 20956 32008 20962 32020
rect 21266 32008 21272 32020
rect 20956 31980 21272 32008
rect 20956 31968 20962 31980
rect 21266 31968 21272 31980
rect 21324 32008 21330 32020
rect 21545 32011 21603 32017
rect 21545 32008 21557 32011
rect 21324 31980 21557 32008
rect 21324 31968 21330 31980
rect 21545 31977 21557 31980
rect 21591 31977 21603 32011
rect 21545 31971 21603 31977
rect 22094 31968 22100 32020
rect 22152 32008 22158 32020
rect 22741 32011 22799 32017
rect 22741 32008 22753 32011
rect 22152 31980 22753 32008
rect 22152 31968 22158 31980
rect 22741 31977 22753 31980
rect 22787 31977 22799 32011
rect 22741 31971 22799 31977
rect 23842 31968 23848 32020
rect 23900 32008 23906 32020
rect 24397 32011 24455 32017
rect 23900 31980 24256 32008
rect 23900 31968 23906 31980
rect 17460 31912 17816 31940
rect 17460 31900 17466 31912
rect 17862 31900 17868 31952
rect 17920 31940 17926 31952
rect 19426 31940 19432 31952
rect 17920 31912 19432 31940
rect 17920 31900 17926 31912
rect 19426 31900 19432 31912
rect 19484 31900 19490 31952
rect 21358 31940 21364 31952
rect 19536 31912 21364 31940
rect 13081 31875 13139 31881
rect 13081 31872 13093 31875
rect 11075 31844 11652 31872
rect 11900 31844 13093 31872
rect 8588 31776 9168 31804
rect 8481 31767 8539 31773
rect 8496 31736 8524 31767
rect 8496 31708 8800 31736
rect 8297 31671 8355 31677
rect 8297 31637 8309 31671
rect 8343 31668 8355 31671
rect 8662 31668 8668 31680
rect 8343 31640 8668 31668
rect 8343 31637 8355 31640
rect 8297 31631 8355 31637
rect 8662 31628 8668 31640
rect 8720 31628 8726 31680
rect 8772 31668 8800 31708
rect 9030 31696 9036 31748
rect 9088 31696 9094 31748
rect 9140 31736 9168 31776
rect 9214 31764 9220 31816
rect 9272 31764 9278 31816
rect 9493 31807 9551 31813
rect 9493 31806 9505 31807
rect 9416 31778 9505 31806
rect 9416 31736 9444 31778
rect 9493 31773 9505 31778
rect 9539 31773 9551 31807
rect 9493 31767 9551 31773
rect 9582 31764 9588 31816
rect 9640 31798 9646 31816
rect 9640 31764 9653 31798
rect 9766 31764 9772 31816
rect 9824 31764 9830 31816
rect 10594 31764 10600 31816
rect 10652 31764 10658 31816
rect 10962 31813 10968 31816
rect 10960 31804 10968 31813
rect 10923 31776 10968 31804
rect 10960 31767 10968 31776
rect 10962 31764 10968 31767
rect 11020 31764 11026 31816
rect 11075 31813 11103 31844
rect 11057 31807 11115 31813
rect 11057 31773 11069 31807
rect 11103 31773 11115 31807
rect 11057 31767 11115 31773
rect 11238 31764 11244 31816
rect 11296 31813 11302 31816
rect 11296 31807 11335 31813
rect 11323 31773 11335 31807
rect 11296 31767 11335 31773
rect 11296 31764 11302 31767
rect 11422 31764 11428 31816
rect 11480 31764 11486 31816
rect 9140 31708 9444 31736
rect 9625 31736 9653 31764
rect 9625 31708 11103 31736
rect 9122 31668 9128 31680
rect 8772 31640 9128 31668
rect 9122 31628 9128 31640
rect 9180 31668 9186 31680
rect 9950 31668 9956 31680
rect 9180 31640 9956 31668
rect 9180 31628 9186 31640
rect 9950 31628 9956 31640
rect 10008 31628 10014 31680
rect 10134 31628 10140 31680
rect 10192 31668 10198 31680
rect 10321 31671 10379 31677
rect 10321 31668 10333 31671
rect 10192 31640 10333 31668
rect 10192 31628 10198 31640
rect 10321 31637 10333 31640
rect 10367 31637 10379 31671
rect 11075 31668 11103 31708
rect 11146 31696 11152 31748
rect 11204 31696 11210 31748
rect 11256 31668 11284 31764
rect 11624 31677 11652 31844
rect 13081 31841 13093 31844
rect 13127 31841 13139 31875
rect 13081 31835 13139 31841
rect 13357 31875 13415 31881
rect 13357 31841 13369 31875
rect 13403 31872 13415 31875
rect 14090 31872 14096 31884
rect 13403 31844 14096 31872
rect 13403 31841 13415 31844
rect 13357 31835 13415 31841
rect 14090 31832 14096 31844
rect 14148 31872 14154 31884
rect 14918 31872 14924 31884
rect 14148 31844 14924 31872
rect 14148 31832 14154 31844
rect 14918 31832 14924 31844
rect 14976 31872 14982 31884
rect 18690 31872 18696 31884
rect 14976 31844 18696 31872
rect 14976 31832 14982 31844
rect 18690 31832 18696 31844
rect 18748 31832 18754 31884
rect 19242 31832 19248 31884
rect 19300 31872 19306 31884
rect 19300 31844 19472 31872
rect 19300 31832 19306 31844
rect 12066 31804 12072 31816
rect 12006 31776 12072 31804
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 13446 31764 13452 31816
rect 13504 31804 13510 31816
rect 13633 31807 13691 31813
rect 13633 31804 13645 31807
rect 13504 31776 13645 31804
rect 13504 31764 13510 31776
rect 13633 31773 13645 31776
rect 13679 31773 13691 31807
rect 13633 31767 13691 31773
rect 15102 31764 15108 31816
rect 15160 31764 15166 31816
rect 15289 31807 15347 31813
rect 15289 31773 15301 31807
rect 15335 31773 15347 31807
rect 15289 31767 15347 31773
rect 12986 31696 12992 31748
rect 13044 31736 13050 31748
rect 14366 31736 14372 31748
rect 13044 31708 14372 31736
rect 13044 31696 13050 31708
rect 14366 31696 14372 31708
rect 14424 31696 14430 31748
rect 11075 31640 11284 31668
rect 11609 31671 11667 31677
rect 10321 31631 10379 31637
rect 11609 31637 11621 31671
rect 11655 31668 11667 31671
rect 11698 31668 11704 31680
rect 11655 31640 11704 31668
rect 11655 31637 11667 31640
rect 11609 31631 11667 31637
rect 11698 31628 11704 31640
rect 11756 31628 11762 31680
rect 15304 31668 15332 31767
rect 15470 31764 15476 31816
rect 15528 31804 15534 31816
rect 15565 31807 15623 31813
rect 15565 31804 15577 31807
rect 15528 31776 15577 31804
rect 15528 31764 15534 31776
rect 15565 31773 15577 31776
rect 15611 31773 15623 31807
rect 15565 31767 15623 31773
rect 15749 31807 15807 31813
rect 15749 31773 15761 31807
rect 15795 31804 15807 31807
rect 17494 31804 17500 31816
rect 15795 31776 17500 31804
rect 15795 31773 15807 31776
rect 15749 31767 15807 31773
rect 17494 31764 17500 31776
rect 17552 31764 17558 31816
rect 17862 31764 17868 31816
rect 17920 31764 17926 31816
rect 19444 31813 19472 31844
rect 19536 31813 19564 31912
rect 21358 31900 21364 31912
rect 21416 31940 21422 31952
rect 21637 31943 21695 31949
rect 21637 31940 21649 31943
rect 21416 31912 21649 31940
rect 21416 31900 21422 31912
rect 21637 31909 21649 31912
rect 21683 31909 21695 31943
rect 21637 31903 21695 31909
rect 22554 31900 22560 31952
rect 22612 31900 22618 31952
rect 24118 31940 24124 31952
rect 22756 31912 24124 31940
rect 20530 31872 20536 31884
rect 19904 31844 20536 31872
rect 19343 31807 19401 31813
rect 19343 31773 19355 31807
rect 19389 31773 19401 31807
rect 19343 31767 19401 31773
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31773 19487 31807
rect 19429 31767 19487 31773
rect 19521 31807 19579 31813
rect 19521 31773 19533 31807
rect 19567 31773 19579 31807
rect 19521 31767 19579 31773
rect 19613 31807 19671 31813
rect 19613 31773 19625 31807
rect 19659 31804 19671 31807
rect 19702 31804 19708 31816
rect 19659 31776 19708 31804
rect 19659 31773 19671 31776
rect 19613 31767 19671 31773
rect 17310 31696 17316 31748
rect 17368 31736 17374 31748
rect 17589 31739 17647 31745
rect 17589 31736 17601 31739
rect 17368 31708 17601 31736
rect 17368 31696 17374 31708
rect 17589 31705 17601 31708
rect 17635 31705 17647 31739
rect 18414 31736 18420 31748
rect 17589 31699 17647 31705
rect 17696 31708 18420 31736
rect 15930 31668 15936 31680
rect 15304 31640 15936 31668
rect 15930 31628 15936 31640
rect 15988 31668 15994 31680
rect 17696 31668 17724 31708
rect 18414 31696 18420 31708
rect 18472 31696 18478 31748
rect 19358 31736 19386 31767
rect 19702 31764 19708 31776
rect 19760 31764 19766 31816
rect 19794 31764 19800 31816
rect 19852 31764 19858 31816
rect 19904 31813 19932 31844
rect 20530 31832 20536 31844
rect 20588 31832 20594 31884
rect 21910 31832 21916 31884
rect 21968 31832 21974 31884
rect 22756 31872 22784 31912
rect 24118 31900 24124 31912
rect 24176 31900 24182 31952
rect 24228 31940 24256 31980
rect 24397 31977 24409 32011
rect 24443 32008 24455 32011
rect 25498 32008 25504 32020
rect 24443 31980 25504 32008
rect 24443 31977 24455 31980
rect 24397 31971 24455 31977
rect 25498 31968 25504 31980
rect 25556 31968 25562 32020
rect 25590 31968 25596 32020
rect 25648 32008 25654 32020
rect 27338 32008 27344 32020
rect 25648 31980 27344 32008
rect 25648 31968 25654 31980
rect 27338 31968 27344 31980
rect 27396 31968 27402 32020
rect 27893 32011 27951 32017
rect 27893 31977 27905 32011
rect 27939 32008 27951 32011
rect 28626 32008 28632 32020
rect 27939 31980 28632 32008
rect 27939 31977 27951 31980
rect 27893 31971 27951 31977
rect 28626 31968 28632 31980
rect 28684 31968 28690 32020
rect 29270 31968 29276 32020
rect 29328 32008 29334 32020
rect 29733 32011 29791 32017
rect 29733 32008 29745 32011
rect 29328 31980 29745 32008
rect 29328 31968 29334 31980
rect 29733 31977 29745 31980
rect 29779 31977 29791 32011
rect 29733 31971 29791 31977
rect 24578 31940 24584 31952
rect 24228 31912 24584 31940
rect 24578 31900 24584 31912
rect 24636 31940 24642 31952
rect 24673 31943 24731 31949
rect 24673 31940 24685 31943
rect 24636 31912 24685 31940
rect 24636 31900 24642 31912
rect 24673 31909 24685 31912
rect 24719 31909 24731 31943
rect 24673 31903 24731 31909
rect 25130 31900 25136 31952
rect 25188 31940 25194 31952
rect 27614 31940 27620 31952
rect 25188 31912 27620 31940
rect 25188 31900 25194 31912
rect 24026 31872 24032 31884
rect 22296 31844 22784 31872
rect 22848 31844 24032 31872
rect 19889 31807 19947 31813
rect 19889 31773 19901 31807
rect 19935 31773 19947 31807
rect 19889 31767 19947 31773
rect 19978 31764 19984 31816
rect 20036 31804 20042 31816
rect 21634 31804 21640 31816
rect 20036 31776 21640 31804
rect 20036 31764 20042 31776
rect 21634 31764 21640 31776
rect 21692 31764 21698 31816
rect 21928 31804 21956 31832
rect 22296 31813 22324 31844
rect 22005 31807 22063 31813
rect 22005 31804 22017 31807
rect 21928 31776 22017 31804
rect 22005 31773 22017 31776
rect 22051 31773 22063 31807
rect 22005 31767 22063 31773
rect 22281 31807 22339 31813
rect 22281 31773 22293 31807
rect 22327 31773 22339 31807
rect 22281 31767 22339 31773
rect 22462 31764 22468 31816
rect 22520 31804 22526 31816
rect 22848 31813 22876 31844
rect 24026 31832 24032 31844
rect 24084 31872 24090 31884
rect 24762 31872 24768 31884
rect 24084 31844 24624 31872
rect 24084 31832 24090 31844
rect 22833 31807 22891 31813
rect 22520 31776 22692 31804
rect 22520 31764 22526 31776
rect 21266 31736 21272 31748
rect 19358 31708 21272 31736
rect 21266 31696 21272 31708
rect 21324 31696 21330 31748
rect 22370 31696 22376 31748
rect 22428 31696 22434 31748
rect 22557 31739 22615 31745
rect 22557 31705 22569 31739
rect 22603 31705 22615 31739
rect 22664 31736 22692 31776
rect 22833 31773 22845 31807
rect 22879 31773 22891 31807
rect 22833 31767 22891 31773
rect 23014 31764 23020 31816
rect 23072 31764 23078 31816
rect 23477 31807 23535 31813
rect 23477 31773 23489 31807
rect 23523 31804 23535 31807
rect 24121 31807 24179 31813
rect 23523 31776 24072 31804
rect 23523 31773 23535 31776
rect 23477 31767 23535 31773
rect 23109 31739 23167 31745
rect 23109 31736 23121 31739
rect 22664 31708 23121 31736
rect 22557 31699 22615 31705
rect 23109 31705 23121 31708
rect 23155 31705 23167 31739
rect 23109 31699 23167 31705
rect 15988 31640 17724 31668
rect 15988 31628 15994 31640
rect 17770 31628 17776 31680
rect 17828 31628 17834 31680
rect 20162 31628 20168 31680
rect 20220 31668 20226 31680
rect 20257 31671 20315 31677
rect 20257 31668 20269 31671
rect 20220 31640 20269 31668
rect 20220 31628 20226 31640
rect 20257 31637 20269 31640
rect 20303 31637 20315 31671
rect 22572 31668 22600 31699
rect 23658 31696 23664 31748
rect 23716 31696 23722 31748
rect 24044 31736 24072 31776
rect 24121 31773 24133 31807
rect 24167 31804 24179 31807
rect 24302 31804 24308 31816
rect 24167 31776 24308 31804
rect 24167 31773 24179 31776
rect 24121 31767 24179 31773
rect 24302 31764 24308 31776
rect 24360 31764 24366 31816
rect 24596 31813 24624 31844
rect 24688 31844 24768 31872
rect 24581 31807 24639 31813
rect 24581 31773 24593 31807
rect 24627 31773 24639 31807
rect 24581 31767 24639 31773
rect 24688 31736 24716 31844
rect 24762 31832 24768 31844
rect 24820 31832 24826 31884
rect 26142 31832 26148 31884
rect 26200 31832 26206 31884
rect 26329 31875 26387 31881
rect 26329 31841 26341 31875
rect 26375 31872 26387 31875
rect 26528 31872 26556 31912
rect 27614 31900 27620 31912
rect 27672 31900 27678 31952
rect 27706 31900 27712 31952
rect 27764 31940 27770 31952
rect 27764 31912 28304 31940
rect 27764 31900 27770 31912
rect 26375 31844 26556 31872
rect 26375 31841 26387 31844
rect 26329 31835 26387 31841
rect 27338 31832 27344 31884
rect 27396 31832 27402 31884
rect 28276 31872 28304 31912
rect 28350 31900 28356 31952
rect 28408 31940 28414 31952
rect 29549 31943 29607 31949
rect 29549 31940 29561 31943
rect 28408 31912 29561 31940
rect 28408 31900 28414 31912
rect 29549 31909 29561 31912
rect 29595 31909 29607 31943
rect 29748 31940 29776 31971
rect 29822 31968 29828 32020
rect 29880 32008 29886 32020
rect 30101 32011 30159 32017
rect 30101 32008 30113 32011
rect 29880 31980 30113 32008
rect 29880 31968 29886 31980
rect 30101 31977 30113 31980
rect 30147 31977 30159 32011
rect 30101 31971 30159 31977
rect 30374 31968 30380 32020
rect 30432 31968 30438 32020
rect 31294 31968 31300 32020
rect 31352 32008 31358 32020
rect 31481 32011 31539 32017
rect 31481 32008 31493 32011
rect 31352 31980 31493 32008
rect 31352 31968 31358 31980
rect 31481 31977 31493 31980
rect 31527 31977 31539 32011
rect 31481 31971 31539 31977
rect 32217 32011 32275 32017
rect 32217 31977 32229 32011
rect 32263 32008 32275 32011
rect 32306 32008 32312 32020
rect 32263 31980 32312 32008
rect 32263 31977 32275 31980
rect 32217 31971 32275 31977
rect 32306 31968 32312 31980
rect 32364 31968 32370 32020
rect 32582 31968 32588 32020
rect 32640 31968 32646 32020
rect 30745 31943 30803 31949
rect 30745 31940 30757 31943
rect 29748 31912 30757 31940
rect 29549 31903 29607 31909
rect 30745 31909 30757 31912
rect 30791 31940 30803 31943
rect 30834 31940 30840 31952
rect 30791 31912 30840 31940
rect 30791 31909 30803 31912
rect 30745 31903 30803 31909
rect 30834 31900 30840 31912
rect 30892 31900 30898 31952
rect 32766 31900 32772 31952
rect 32824 31900 32830 31952
rect 27632 31844 28212 31872
rect 28276 31844 28396 31872
rect 24857 31807 24915 31813
rect 24857 31804 24869 31807
rect 24835 31776 24869 31804
rect 24857 31773 24869 31776
rect 24903 31773 24915 31807
rect 24857 31767 24915 31773
rect 25041 31807 25099 31813
rect 25041 31773 25053 31807
rect 25087 31773 25099 31807
rect 25041 31767 25099 31773
rect 24044 31708 24716 31736
rect 24762 31696 24768 31748
rect 24820 31736 24826 31748
rect 24872 31736 24900 31767
rect 24820 31708 24900 31736
rect 24820 31696 24826 31708
rect 24946 31696 24952 31748
rect 25004 31736 25010 31748
rect 25056 31736 25084 31767
rect 25314 31764 25320 31816
rect 25372 31804 25378 31816
rect 25593 31807 25651 31813
rect 25593 31804 25605 31807
rect 25372 31776 25605 31804
rect 25372 31764 25378 31776
rect 25593 31773 25605 31776
rect 25639 31773 25651 31807
rect 25593 31767 25651 31773
rect 25682 31764 25688 31816
rect 25740 31764 25746 31816
rect 25866 31764 25872 31816
rect 25924 31764 25930 31816
rect 25961 31807 26019 31813
rect 25961 31773 25973 31807
rect 26007 31804 26019 31807
rect 26160 31804 26188 31832
rect 27632 31816 27660 31844
rect 26007 31776 26188 31804
rect 26237 31807 26295 31813
rect 26007 31773 26019 31776
rect 25961 31767 26019 31773
rect 26237 31773 26249 31807
rect 26283 31773 26295 31807
rect 26237 31767 26295 31773
rect 26142 31736 26148 31748
rect 25004 31708 26148 31736
rect 25004 31696 25010 31708
rect 26142 31696 26148 31708
rect 26200 31696 26206 31748
rect 26252 31736 26280 31767
rect 26418 31764 26424 31816
rect 26476 31764 26482 31816
rect 26513 31807 26571 31813
rect 26513 31773 26525 31807
rect 26559 31804 26571 31807
rect 26789 31807 26847 31813
rect 26789 31804 26801 31807
rect 26559 31776 26801 31804
rect 26559 31773 26571 31776
rect 26513 31767 26571 31773
rect 26789 31773 26801 31776
rect 26835 31773 26847 31807
rect 26789 31767 26847 31773
rect 26973 31807 27031 31813
rect 26973 31773 26985 31807
rect 27019 31804 27031 31807
rect 27062 31804 27068 31816
rect 27019 31776 27068 31804
rect 27019 31773 27031 31776
rect 26973 31767 27031 31773
rect 27062 31764 27068 31776
rect 27120 31764 27126 31816
rect 27154 31764 27160 31816
rect 27212 31764 27218 31816
rect 27246 31764 27252 31816
rect 27304 31764 27310 31816
rect 27430 31764 27436 31816
rect 27488 31764 27494 31816
rect 27614 31764 27620 31816
rect 27672 31764 27678 31816
rect 28074 31804 28080 31816
rect 27724 31776 28080 31804
rect 27724 31736 27752 31776
rect 28074 31764 28080 31776
rect 28132 31764 28138 31816
rect 28184 31813 28212 31844
rect 28169 31807 28227 31813
rect 28169 31773 28181 31807
rect 28215 31773 28227 31807
rect 28169 31767 28227 31773
rect 28258 31764 28264 31816
rect 28316 31764 28322 31816
rect 28368 31804 28396 31844
rect 28534 31832 28540 31884
rect 28592 31872 28598 31884
rect 28902 31872 28908 31884
rect 28592 31844 28908 31872
rect 28592 31832 28598 31844
rect 28902 31832 28908 31844
rect 28960 31832 28966 31884
rect 30392 31844 31064 31872
rect 30392 31816 30420 31844
rect 31036 31816 31064 31844
rect 31110 31832 31116 31884
rect 31168 31832 31174 31884
rect 31386 31832 31392 31884
rect 31444 31872 31450 31884
rect 31570 31872 31576 31884
rect 31444 31844 31576 31872
rect 31444 31832 31450 31844
rect 31570 31832 31576 31844
rect 31628 31832 31634 31884
rect 28718 31804 28724 31816
rect 28368 31776 28724 31804
rect 28718 31764 28724 31776
rect 28776 31764 28782 31816
rect 28810 31764 28816 31816
rect 28868 31804 28874 31816
rect 28868 31776 29500 31804
rect 28868 31764 28874 31776
rect 29472 31770 29500 31776
rect 29687 31773 29745 31779
rect 29687 31770 29699 31773
rect 28442 31745 28448 31748
rect 26252 31708 27752 31736
rect 28399 31739 28448 31745
rect 28399 31705 28411 31739
rect 28445 31705 28448 31739
rect 28399 31699 28448 31705
rect 28442 31696 28448 31699
rect 28500 31696 28506 31748
rect 29089 31739 29147 31745
rect 28552 31708 28948 31736
rect 23750 31668 23756 31680
rect 22572 31640 23756 31668
rect 20257 31631 20315 31637
rect 23750 31628 23756 31640
rect 23808 31628 23814 31680
rect 24029 31671 24087 31677
rect 24029 31637 24041 31671
rect 24075 31668 24087 31671
rect 24578 31668 24584 31680
rect 24075 31640 24584 31668
rect 24075 31637 24087 31640
rect 24029 31631 24087 31637
rect 24578 31628 24584 31640
rect 24636 31628 24642 31680
rect 25222 31628 25228 31680
rect 25280 31628 25286 31680
rect 25409 31671 25467 31677
rect 25409 31637 25421 31671
rect 25455 31668 25467 31671
rect 25682 31668 25688 31680
rect 25455 31640 25688 31668
rect 25455 31637 25467 31640
rect 25409 31631 25467 31637
rect 25682 31628 25688 31640
rect 25740 31628 25746 31680
rect 25774 31628 25780 31680
rect 25832 31668 25838 31680
rect 26053 31671 26111 31677
rect 26053 31668 26065 31671
rect 25832 31640 26065 31668
rect 25832 31628 25838 31640
rect 26053 31637 26065 31640
rect 26099 31637 26111 31671
rect 26053 31631 26111 31637
rect 26510 31628 26516 31680
rect 26568 31668 26574 31680
rect 27522 31668 27528 31680
rect 26568 31640 27528 31668
rect 26568 31628 26574 31640
rect 27522 31628 27528 31640
rect 27580 31668 27586 31680
rect 28552 31668 28580 31708
rect 27580 31640 28580 31668
rect 27580 31628 27586 31640
rect 28810 31628 28816 31680
rect 28868 31628 28874 31680
rect 28920 31668 28948 31708
rect 29089 31705 29101 31739
rect 29135 31736 29147 31739
rect 29362 31736 29368 31748
rect 29135 31708 29368 31736
rect 29135 31705 29147 31708
rect 29089 31699 29147 31705
rect 29362 31696 29368 31708
rect 29420 31696 29426 31748
rect 29472 31742 29699 31770
rect 29687 31739 29699 31742
rect 29733 31739 29745 31773
rect 30006 31764 30012 31816
rect 30064 31764 30070 31816
rect 30098 31764 30104 31816
rect 30156 31804 30162 31816
rect 30374 31804 30380 31816
rect 30156 31776 30380 31804
rect 30156 31764 30162 31776
rect 30374 31764 30380 31776
rect 30432 31764 30438 31816
rect 30466 31764 30472 31816
rect 30524 31764 30530 31816
rect 30926 31804 30932 31816
rect 30887 31776 30932 31804
rect 30926 31764 30932 31776
rect 30984 31764 30990 31816
rect 31018 31764 31024 31816
rect 31076 31804 31082 31816
rect 31205 31807 31263 31813
rect 31205 31804 31217 31807
rect 31076 31776 31217 31804
rect 31076 31764 31082 31776
rect 31205 31773 31217 31776
rect 31251 31773 31263 31807
rect 31205 31767 31263 31773
rect 31294 31764 31300 31816
rect 31352 31804 31358 31816
rect 31352 31776 31708 31804
rect 31352 31764 31358 31776
rect 29687 31733 29745 31739
rect 29822 31696 29828 31748
rect 29880 31736 29886 31748
rect 29917 31739 29975 31745
rect 29917 31736 29929 31739
rect 29880 31708 29929 31736
rect 29880 31696 29886 31708
rect 29917 31705 29929 31708
rect 29963 31705 29975 31739
rect 31478 31736 31484 31748
rect 29917 31699 29975 31705
rect 30392 31708 31484 31736
rect 30392 31668 30420 31708
rect 31478 31696 31484 31708
rect 31536 31696 31542 31748
rect 31680 31736 31708 31776
rect 31846 31764 31852 31816
rect 31904 31804 31910 31816
rect 32033 31807 32091 31813
rect 32033 31804 32045 31807
rect 31904 31776 32045 31804
rect 31904 31764 31910 31776
rect 32033 31773 32045 31776
rect 32079 31773 32091 31807
rect 32033 31767 32091 31773
rect 32217 31807 32275 31813
rect 32217 31773 32229 31807
rect 32263 31773 32275 31807
rect 32217 31767 32275 31773
rect 31864 31736 31892 31764
rect 31680 31708 31892 31736
rect 28920 31640 30420 31668
rect 30466 31628 30472 31680
rect 30524 31668 30530 31680
rect 31297 31671 31355 31677
rect 31297 31668 31309 31671
rect 30524 31640 31309 31668
rect 30524 31628 30530 31640
rect 31297 31637 31309 31640
rect 31343 31637 31355 31671
rect 31297 31631 31355 31637
rect 31386 31628 31392 31680
rect 31444 31668 31450 31680
rect 32232 31668 32260 31767
rect 32306 31764 32312 31816
rect 32364 31804 32370 31816
rect 32674 31804 32680 31816
rect 32364 31776 32680 31804
rect 32364 31764 32370 31776
rect 32674 31764 32680 31776
rect 32732 31764 32738 31816
rect 32398 31696 32404 31748
rect 32456 31696 32462 31748
rect 31444 31640 32260 31668
rect 31444 31628 31450 31640
rect 32582 31628 32588 31680
rect 32640 31677 32646 31680
rect 32640 31671 32659 31677
rect 32647 31637 32659 31671
rect 32640 31631 32659 31637
rect 32640 31628 32646 31631
rect 1104 31578 36432 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 36432 31578
rect 1104 31504 36432 31526
rect 4246 31464 4252 31476
rect 3804 31436 4252 31464
rect 1302 31356 1308 31408
rect 1360 31396 1366 31408
rect 2225 31399 2283 31405
rect 2225 31396 2237 31399
rect 1360 31368 2237 31396
rect 1360 31356 1366 31368
rect 2225 31365 2237 31368
rect 2271 31365 2283 31399
rect 2225 31359 2283 31365
rect 2406 31356 2412 31408
rect 2464 31356 2470 31408
rect 3804 31396 3832 31436
rect 4246 31424 4252 31436
rect 4304 31424 4310 31476
rect 4525 31467 4583 31473
rect 4525 31433 4537 31467
rect 4571 31464 4583 31467
rect 5718 31464 5724 31476
rect 4571 31436 5724 31464
rect 4571 31433 4583 31436
rect 4525 31427 4583 31433
rect 5718 31424 5724 31436
rect 5776 31424 5782 31476
rect 6733 31467 6791 31473
rect 6733 31433 6745 31467
rect 6779 31464 6791 31467
rect 6822 31464 6828 31476
rect 6779 31436 6828 31464
rect 6779 31433 6791 31436
rect 6733 31427 6791 31433
rect 6822 31424 6828 31436
rect 6880 31424 6886 31476
rect 6914 31424 6920 31476
rect 6972 31424 6978 31476
rect 7650 31464 7656 31476
rect 7116 31436 7656 31464
rect 3726 31368 3832 31396
rect 4154 31356 4160 31408
rect 4212 31356 4218 31408
rect 4614 31356 4620 31408
rect 4672 31396 4678 31408
rect 5534 31396 5540 31408
rect 4672 31368 4844 31396
rect 4672 31356 4678 31368
rect 2041 31331 2099 31337
rect 2041 31297 2053 31331
rect 2087 31297 2099 31331
rect 2041 31291 2099 31297
rect 2317 31331 2375 31337
rect 2317 31297 2329 31331
rect 2363 31297 2375 31331
rect 2317 31291 2375 31297
rect 4433 31331 4491 31337
rect 4433 31297 4445 31331
rect 4479 31328 4491 31331
rect 4706 31328 4712 31340
rect 4479 31300 4712 31328
rect 4479 31297 4491 31300
rect 4433 31291 4491 31297
rect 2056 31192 2084 31291
rect 2332 31260 2360 31291
rect 4706 31288 4712 31300
rect 4764 31288 4770 31340
rect 4816 31337 4844 31368
rect 5000 31368 5540 31396
rect 5000 31337 5028 31368
rect 5534 31356 5540 31368
rect 5592 31356 5598 31408
rect 4801 31331 4859 31337
rect 4801 31297 4813 31331
rect 4847 31297 4859 31331
rect 4801 31291 4859 31297
rect 4893 31331 4951 31337
rect 4893 31297 4905 31331
rect 4939 31297 4951 31331
rect 4893 31291 4951 31297
rect 4985 31331 5043 31337
rect 4985 31297 4997 31331
rect 5031 31297 5043 31331
rect 4985 31291 5043 31297
rect 2774 31260 2780 31272
rect 2332 31232 2780 31260
rect 2774 31220 2780 31232
rect 2832 31260 2838 31272
rect 4062 31260 4068 31272
rect 2832 31232 4068 31260
rect 2832 31220 2838 31232
rect 4062 31220 4068 31232
rect 4120 31220 4126 31272
rect 4614 31220 4620 31272
rect 4672 31260 4678 31272
rect 4908 31260 4936 31291
rect 5166 31288 5172 31340
rect 5224 31288 5230 31340
rect 5629 31331 5687 31337
rect 5629 31297 5641 31331
rect 5675 31297 5687 31331
rect 5629 31291 5687 31297
rect 4672 31232 4936 31260
rect 5445 31263 5503 31269
rect 4672 31220 4678 31232
rect 5445 31229 5457 31263
rect 5491 31229 5503 31263
rect 5445 31223 5503 31229
rect 2958 31192 2964 31204
rect 2056 31164 2964 31192
rect 2958 31152 2964 31164
rect 3016 31152 3022 31204
rect 5460 31192 5488 31223
rect 5534 31220 5540 31272
rect 5592 31220 5598 31272
rect 5644 31260 5672 31291
rect 6270 31288 6276 31340
rect 6328 31328 6334 31340
rect 6365 31331 6423 31337
rect 6365 31328 6377 31331
rect 6328 31300 6377 31328
rect 6328 31288 6334 31300
rect 6365 31297 6377 31300
rect 6411 31297 6423 31331
rect 6365 31291 6423 31297
rect 6546 31288 6552 31340
rect 6604 31328 6610 31340
rect 6822 31328 6828 31340
rect 6604 31300 6828 31328
rect 6604 31288 6610 31300
rect 6822 31288 6828 31300
rect 6880 31288 6886 31340
rect 7116 31337 7144 31436
rect 7650 31424 7656 31436
rect 7708 31424 7714 31476
rect 7926 31424 7932 31476
rect 7984 31464 7990 31476
rect 7984 31436 8708 31464
rect 7984 31424 7990 31436
rect 7466 31356 7472 31408
rect 7524 31396 7530 31408
rect 7561 31399 7619 31405
rect 7561 31396 7573 31399
rect 7524 31368 7573 31396
rect 7524 31356 7530 31368
rect 7561 31365 7573 31368
rect 7607 31365 7619 31399
rect 8680 31396 8708 31436
rect 9214 31424 9220 31476
rect 9272 31464 9278 31476
rect 9585 31467 9643 31473
rect 9585 31464 9597 31467
rect 9272 31436 9597 31464
rect 9272 31424 9278 31436
rect 9585 31433 9597 31436
rect 9631 31433 9643 31467
rect 9585 31427 9643 31433
rect 9674 31424 9680 31476
rect 9732 31464 9738 31476
rect 9769 31467 9827 31473
rect 9769 31464 9781 31467
rect 9732 31436 9781 31464
rect 9732 31424 9738 31436
rect 9769 31433 9781 31436
rect 9815 31433 9827 31467
rect 9769 31427 9827 31433
rect 10042 31424 10048 31476
rect 10100 31464 10106 31476
rect 10597 31467 10655 31473
rect 10597 31464 10609 31467
rect 10100 31436 10609 31464
rect 10100 31424 10106 31436
rect 10597 31433 10609 31436
rect 10643 31433 10655 31467
rect 10597 31427 10655 31433
rect 11241 31467 11299 31473
rect 11241 31433 11253 31467
rect 11287 31464 11299 31467
rect 11790 31464 11796 31476
rect 11287 31436 11796 31464
rect 11287 31433 11299 31436
rect 11241 31427 11299 31433
rect 11790 31424 11796 31436
rect 11848 31424 11854 31476
rect 13906 31424 13912 31476
rect 13964 31464 13970 31476
rect 13964 31436 14320 31464
rect 13964 31424 13970 31436
rect 10870 31396 10876 31408
rect 8680 31368 10876 31396
rect 7561 31359 7619 31365
rect 10870 31356 10876 31368
rect 10928 31356 10934 31408
rect 14292 31396 14320 31436
rect 14366 31424 14372 31476
rect 14424 31464 14430 31476
rect 19334 31464 19340 31476
rect 14424 31436 19340 31464
rect 14424 31424 14430 31436
rect 19334 31424 19340 31436
rect 19392 31424 19398 31476
rect 19889 31467 19947 31473
rect 19889 31433 19901 31467
rect 19935 31464 19947 31467
rect 21082 31464 21088 31476
rect 19935 31436 21088 31464
rect 19935 31433 19947 31436
rect 19889 31427 19947 31433
rect 21082 31424 21088 31436
rect 21140 31424 21146 31476
rect 21174 31424 21180 31476
rect 21232 31464 21238 31476
rect 24302 31464 24308 31476
rect 21232 31436 24308 31464
rect 21232 31424 21238 31436
rect 24302 31424 24308 31436
rect 24360 31424 24366 31476
rect 25685 31467 25743 31473
rect 25685 31464 25697 31467
rect 24688 31436 25697 31464
rect 15013 31399 15071 31405
rect 15013 31396 15025 31399
rect 10980 31368 11744 31396
rect 14214 31368 15025 31396
rect 7101 31331 7159 31337
rect 7101 31297 7113 31331
rect 7147 31297 7159 31331
rect 7101 31291 7159 31297
rect 7374 31288 7380 31340
rect 7432 31288 7438 31340
rect 7834 31288 7840 31340
rect 7892 31328 7898 31340
rect 8297 31331 8355 31337
rect 8297 31328 8309 31331
rect 7892 31300 8309 31328
rect 7892 31288 7898 31300
rect 8297 31297 8309 31300
rect 8343 31297 8355 31331
rect 8297 31291 8355 31297
rect 8478 31288 8484 31340
rect 8536 31288 8542 31340
rect 8573 31331 8631 31337
rect 8573 31297 8585 31331
rect 8619 31328 8631 31331
rect 8619 31300 8892 31328
rect 8619 31297 8631 31300
rect 8573 31291 8631 31297
rect 6914 31260 6920 31272
rect 5644 31232 6920 31260
rect 6914 31220 6920 31232
rect 6972 31220 6978 31272
rect 7193 31263 7251 31269
rect 7193 31229 7205 31263
rect 7239 31260 7251 31263
rect 7558 31260 7564 31272
rect 7239 31232 7564 31260
rect 7239 31229 7251 31232
rect 7193 31223 7251 31229
rect 7558 31220 7564 31232
rect 7616 31220 7622 31272
rect 5718 31192 5724 31204
rect 5460 31164 5724 31192
rect 5718 31152 5724 31164
rect 5776 31152 5782 31204
rect 7285 31195 7343 31201
rect 7285 31161 7297 31195
rect 7331 31192 7343 31195
rect 7466 31192 7472 31204
rect 7331 31164 7472 31192
rect 7331 31161 7343 31164
rect 7285 31155 7343 31161
rect 7466 31152 7472 31164
rect 7524 31152 7530 31204
rect 7929 31195 7987 31201
rect 7929 31161 7941 31195
rect 7975 31192 7987 31195
rect 8113 31195 8171 31201
rect 8113 31192 8125 31195
rect 7975 31164 8125 31192
rect 7975 31161 7987 31164
rect 7929 31155 7987 31161
rect 8113 31161 8125 31164
rect 8159 31161 8171 31195
rect 8113 31155 8171 31161
rect 8570 31152 8576 31204
rect 8628 31192 8634 31204
rect 8665 31195 8723 31201
rect 8665 31192 8677 31195
rect 8628 31164 8677 31192
rect 8628 31152 8634 31164
rect 8665 31161 8677 31164
rect 8711 31161 8723 31195
rect 8864 31192 8892 31300
rect 8938 31288 8944 31340
rect 8996 31288 9002 31340
rect 9122 31288 9128 31340
rect 9180 31288 9186 31340
rect 9214 31288 9220 31340
rect 9272 31288 9278 31340
rect 9401 31331 9459 31337
rect 9401 31297 9413 31331
rect 9447 31297 9459 31331
rect 9401 31291 9459 31297
rect 9033 31263 9091 31269
rect 9033 31229 9045 31263
rect 9079 31260 9091 31263
rect 9416 31260 9444 31291
rect 9490 31288 9496 31340
rect 9548 31328 9554 31340
rect 9710 31331 9768 31337
rect 9710 31328 9722 31331
rect 9548 31300 9722 31328
rect 9548 31288 9554 31300
rect 9710 31297 9722 31300
rect 9756 31297 9768 31331
rect 9710 31291 9768 31297
rect 9950 31288 9956 31340
rect 10008 31328 10014 31340
rect 10686 31328 10692 31340
rect 10008 31300 10692 31328
rect 10008 31288 10014 31300
rect 10686 31288 10692 31300
rect 10744 31328 10750 31340
rect 10980 31337 11008 31368
rect 11716 31340 11744 31368
rect 15013 31365 15025 31368
rect 15059 31365 15071 31399
rect 17586 31396 17592 31408
rect 15013 31359 15071 31365
rect 16960 31368 17592 31396
rect 10781 31331 10839 31337
rect 10781 31328 10793 31331
rect 10744 31300 10793 31328
rect 10744 31288 10750 31300
rect 10781 31297 10793 31300
rect 10827 31297 10839 31331
rect 10781 31291 10839 31297
rect 10965 31331 11023 31337
rect 10965 31297 10977 31331
rect 11011 31297 11023 31331
rect 10965 31291 11023 31297
rect 11149 31331 11207 31337
rect 11149 31297 11161 31331
rect 11195 31297 11207 31331
rect 11149 31291 11207 31297
rect 9079 31232 9444 31260
rect 9079 31229 9091 31232
rect 9033 31223 9091 31229
rect 10134 31220 10140 31272
rect 10192 31260 10198 31272
rect 10229 31263 10287 31269
rect 10229 31260 10241 31263
rect 10192 31232 10241 31260
rect 10192 31220 10198 31232
rect 10229 31229 10241 31232
rect 10275 31260 10287 31263
rect 10502 31260 10508 31272
rect 10275 31232 10508 31260
rect 10275 31229 10287 31232
rect 10229 31223 10287 31229
rect 10502 31220 10508 31232
rect 10560 31220 10566 31272
rect 9122 31192 9128 31204
rect 8864 31164 9128 31192
rect 8665 31155 8723 31161
rect 9122 31152 9128 31164
rect 9180 31152 9186 31204
rect 9401 31195 9459 31201
rect 9401 31161 9413 31195
rect 9447 31192 9459 31195
rect 9766 31192 9772 31204
rect 9447 31164 9772 31192
rect 9447 31161 9459 31164
rect 9401 31155 9459 31161
rect 9766 31152 9772 31164
rect 9824 31152 9830 31204
rect 11164 31192 11192 31291
rect 11330 31288 11336 31340
rect 11388 31288 11394 31340
rect 11698 31288 11704 31340
rect 11756 31288 11762 31340
rect 11974 31328 11980 31340
rect 11808 31300 11980 31328
rect 11808 31269 11836 31300
rect 11974 31288 11980 31300
rect 12032 31288 12038 31340
rect 12345 31331 12403 31337
rect 12345 31297 12357 31331
rect 12391 31297 12403 31331
rect 12345 31291 12403 31297
rect 11793 31263 11851 31269
rect 11793 31229 11805 31263
rect 11839 31229 11851 31263
rect 11793 31223 11851 31229
rect 11882 31220 11888 31272
rect 11940 31260 11946 31272
rect 12069 31263 12127 31269
rect 12069 31260 12081 31263
rect 11940 31232 12081 31260
rect 11940 31220 11946 31232
rect 12069 31229 12081 31232
rect 12115 31260 12127 31263
rect 12360 31260 12388 31291
rect 14918 31288 14924 31340
rect 14976 31288 14982 31340
rect 15378 31288 15384 31340
rect 15436 31288 15442 31340
rect 12115 31232 12388 31260
rect 12529 31263 12587 31269
rect 12115 31229 12127 31232
rect 12069 31223 12127 31229
rect 12529 31229 12541 31263
rect 12575 31260 12587 31263
rect 13173 31263 13231 31269
rect 13173 31260 13185 31263
rect 12575 31232 13185 31260
rect 12575 31229 12587 31232
rect 12529 31223 12587 31229
rect 13173 31229 13185 31232
rect 13219 31229 13231 31263
rect 13173 31223 13231 31229
rect 11164 31164 12296 31192
rect 1762 31084 1768 31136
rect 1820 31124 1826 31136
rect 1857 31127 1915 31133
rect 1857 31124 1869 31127
rect 1820 31096 1869 31124
rect 1820 31084 1826 31096
rect 1857 31093 1869 31096
rect 1903 31093 1915 31127
rect 1857 31087 1915 31093
rect 4890 31084 4896 31136
rect 4948 31124 4954 31136
rect 5626 31124 5632 31136
rect 4948 31096 5632 31124
rect 4948 31084 4954 31096
rect 5626 31084 5632 31096
rect 5684 31084 5690 31136
rect 5810 31084 5816 31136
rect 5868 31124 5874 31136
rect 5997 31127 6055 31133
rect 5997 31124 6009 31127
rect 5868 31096 6009 31124
rect 5868 31084 5874 31096
rect 5997 31093 6009 31096
rect 6043 31093 6055 31127
rect 5997 31087 6055 31093
rect 6086 31084 6092 31136
rect 6144 31124 6150 31136
rect 8021 31127 8079 31133
rect 8021 31124 8033 31127
rect 6144 31096 8033 31124
rect 6144 31084 6150 31096
rect 8021 31093 8033 31096
rect 8067 31093 8079 31127
rect 8021 31087 8079 31093
rect 8478 31084 8484 31136
rect 8536 31084 8542 31136
rect 9030 31084 9036 31136
rect 9088 31124 9094 31136
rect 10137 31127 10195 31133
rect 10137 31124 10149 31127
rect 9088 31096 10149 31124
rect 9088 31084 9094 31096
rect 10137 31093 10149 31096
rect 10183 31093 10195 31127
rect 10137 31087 10195 31093
rect 11330 31084 11336 31136
rect 11388 31124 11394 31136
rect 12161 31127 12219 31133
rect 12161 31124 12173 31127
rect 11388 31096 12173 31124
rect 11388 31084 11394 31096
rect 12161 31093 12173 31096
rect 12207 31093 12219 31127
rect 12268 31124 12296 31164
rect 12342 31152 12348 31204
rect 12400 31192 12406 31204
rect 12544 31192 12572 31223
rect 13906 31220 13912 31272
rect 13964 31260 13970 31272
rect 14645 31263 14703 31269
rect 14645 31260 14657 31263
rect 13964 31232 14657 31260
rect 13964 31220 13970 31232
rect 14645 31229 14657 31232
rect 14691 31229 14703 31263
rect 14645 31223 14703 31229
rect 15654 31220 15660 31272
rect 15712 31260 15718 31272
rect 16206 31260 16212 31272
rect 15712 31232 16212 31260
rect 15712 31220 15718 31232
rect 16206 31220 16212 31232
rect 16264 31260 16270 31272
rect 16960 31269 16988 31368
rect 17586 31356 17592 31368
rect 17644 31356 17650 31408
rect 17770 31356 17776 31408
rect 17828 31396 17834 31408
rect 20993 31399 21051 31405
rect 20993 31396 21005 31399
rect 17828 31368 21005 31396
rect 17828 31356 17834 31368
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31297 17187 31331
rect 17129 31291 17187 31297
rect 16945 31263 17003 31269
rect 16945 31260 16957 31263
rect 16264 31232 16957 31260
rect 16264 31220 16270 31232
rect 16945 31229 16957 31232
rect 16991 31229 17003 31263
rect 17144 31260 17172 31291
rect 17862 31288 17868 31340
rect 17920 31328 17926 31340
rect 18601 31331 18659 31337
rect 18601 31328 18613 31331
rect 17920 31300 18613 31328
rect 17920 31288 17926 31300
rect 18601 31297 18613 31300
rect 18647 31297 18659 31331
rect 18601 31291 18659 31297
rect 18782 31288 18788 31340
rect 18840 31288 18846 31340
rect 18874 31288 18880 31340
rect 18932 31288 18938 31340
rect 18989 31331 19047 31337
rect 18989 31297 19001 31331
rect 19035 31328 19047 31331
rect 19076 31328 19104 31368
rect 20993 31365 21005 31368
rect 21039 31365 21051 31399
rect 22094 31396 22100 31408
rect 20993 31359 21051 31365
rect 21284 31368 22100 31396
rect 21284 31340 21312 31368
rect 22094 31356 22100 31368
rect 22152 31356 22158 31408
rect 24688 31405 24716 31436
rect 25685 31433 25697 31436
rect 25731 31433 25743 31467
rect 25685 31427 25743 31433
rect 25866 31424 25872 31476
rect 25924 31464 25930 31476
rect 26973 31467 27031 31473
rect 26973 31464 26985 31467
rect 25924 31436 26985 31464
rect 25924 31424 25930 31436
rect 26973 31433 26985 31436
rect 27019 31433 27031 31467
rect 26973 31427 27031 31433
rect 27890 31424 27896 31476
rect 27948 31464 27954 31476
rect 30742 31464 30748 31476
rect 27948 31436 28121 31464
rect 27948 31424 27954 31436
rect 24673 31399 24731 31405
rect 24673 31365 24685 31399
rect 24719 31365 24731 31399
rect 24673 31359 24731 31365
rect 25314 31356 25320 31408
rect 25372 31356 25378 31408
rect 25409 31399 25467 31405
rect 25409 31365 25421 31399
rect 25455 31396 25467 31399
rect 25777 31399 25835 31405
rect 25777 31396 25789 31399
rect 25455 31368 25789 31396
rect 25455 31365 25467 31368
rect 25409 31359 25467 31365
rect 25777 31365 25789 31368
rect 25823 31365 25835 31399
rect 25777 31359 25835 31365
rect 25961 31399 26019 31405
rect 25961 31365 25973 31399
rect 26007 31396 26019 31399
rect 26602 31396 26608 31408
rect 26007 31368 26608 31396
rect 26007 31365 26019 31368
rect 25961 31359 26019 31365
rect 26602 31356 26608 31368
rect 26660 31356 26666 31408
rect 26694 31356 26700 31408
rect 26752 31396 26758 31408
rect 27125 31399 27183 31405
rect 27125 31396 27137 31399
rect 26752 31368 27137 31396
rect 26752 31356 26758 31368
rect 27125 31365 27137 31368
rect 27171 31365 27183 31399
rect 27125 31359 27183 31365
rect 27341 31399 27399 31405
rect 27341 31365 27353 31399
rect 27387 31365 27399 31399
rect 27341 31359 27399 31365
rect 19035 31300 19104 31328
rect 20073 31331 20131 31337
rect 19035 31297 19047 31300
rect 18989 31291 19047 31297
rect 20073 31297 20085 31331
rect 20119 31297 20131 31331
rect 20073 31291 20131 31297
rect 18046 31260 18052 31272
rect 17144 31232 18052 31260
rect 16945 31223 17003 31229
rect 18046 31220 18052 31232
rect 18104 31220 18110 31272
rect 18693 31263 18751 31269
rect 18693 31229 18705 31263
rect 18739 31260 18751 31263
rect 20088 31260 20116 31291
rect 20162 31288 20168 31340
rect 20220 31288 20226 31340
rect 20254 31288 20260 31340
rect 20312 31328 20318 31340
rect 20349 31331 20407 31337
rect 20349 31328 20361 31331
rect 20312 31300 20361 31328
rect 20312 31288 20318 31300
rect 20349 31297 20361 31300
rect 20395 31297 20407 31331
rect 20349 31291 20407 31297
rect 20438 31288 20444 31340
rect 20496 31288 20502 31340
rect 20533 31331 20591 31337
rect 20533 31297 20545 31331
rect 20579 31297 20591 31331
rect 20533 31291 20591 31297
rect 18739 31232 20116 31260
rect 18739 31229 18751 31232
rect 18693 31223 18751 31229
rect 12400 31164 12572 31192
rect 12400 31152 12406 31164
rect 15746 31152 15752 31204
rect 15804 31192 15810 31204
rect 18064 31192 18092 31220
rect 19150 31192 19156 31204
rect 15804 31164 17356 31192
rect 18064 31164 19156 31192
rect 15804 31152 15810 31164
rect 17328 31136 17356 31164
rect 19150 31152 19156 31164
rect 19208 31192 19214 31204
rect 20548 31192 20576 31291
rect 20714 31288 20720 31340
rect 20772 31288 20778 31340
rect 20809 31331 20867 31337
rect 20809 31297 20821 31331
rect 20855 31297 20867 31331
rect 20809 31291 20867 31297
rect 20622 31220 20628 31272
rect 20680 31260 20686 31272
rect 20824 31260 20852 31291
rect 20898 31288 20904 31340
rect 20956 31288 20962 31340
rect 21085 31331 21143 31337
rect 21085 31297 21097 31331
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 21177 31331 21235 31337
rect 21177 31297 21189 31331
rect 21223 31328 21235 31331
rect 21266 31328 21272 31340
rect 21223 31300 21272 31328
rect 21223 31297 21235 31300
rect 21177 31291 21235 31297
rect 20680 31232 20852 31260
rect 20680 31220 20686 31232
rect 19208 31164 20576 31192
rect 19208 31152 19214 31164
rect 20806 31152 20812 31204
rect 20864 31192 20870 31204
rect 21100 31192 21128 31291
rect 21266 31288 21272 31300
rect 21324 31288 21330 31340
rect 21361 31331 21419 31337
rect 21361 31297 21373 31331
rect 21407 31297 21419 31331
rect 21361 31291 21419 31297
rect 22925 31331 22983 31337
rect 22925 31297 22937 31331
rect 22971 31328 22983 31331
rect 23198 31328 23204 31340
rect 22971 31300 23204 31328
rect 22971 31297 22983 31300
rect 22925 31291 22983 31297
rect 21177 31195 21235 31201
rect 21177 31192 21189 31195
rect 20864 31164 21189 31192
rect 20864 31152 20870 31164
rect 21177 31161 21189 31164
rect 21223 31161 21235 31195
rect 21177 31155 21235 31161
rect 13262 31124 13268 31136
rect 12268 31096 13268 31124
rect 12161 31087 12219 31093
rect 13262 31084 13268 31096
rect 13320 31084 13326 31136
rect 14274 31084 14280 31136
rect 14332 31124 14338 31136
rect 16850 31124 16856 31136
rect 14332 31096 16856 31124
rect 14332 31084 14338 31096
rect 16850 31084 16856 31096
rect 16908 31084 16914 31136
rect 17310 31084 17316 31136
rect 17368 31084 17374 31136
rect 17586 31084 17592 31136
rect 17644 31124 17650 31136
rect 18782 31124 18788 31136
rect 17644 31096 18788 31124
rect 17644 31084 17650 31096
rect 18782 31084 18788 31096
rect 18840 31084 18846 31136
rect 20530 31084 20536 31136
rect 20588 31084 20594 31136
rect 20714 31084 20720 31136
rect 20772 31124 20778 31136
rect 21376 31124 21404 31291
rect 23198 31288 23204 31300
rect 23256 31288 23262 31340
rect 23566 31288 23572 31340
rect 23624 31288 23630 31340
rect 25199 31331 25257 31337
rect 25199 31297 25211 31331
rect 25245 31328 25257 31331
rect 25501 31331 25559 31337
rect 25245 31300 25452 31328
rect 25245 31297 25257 31300
rect 25199 31291 25257 31297
rect 23014 31220 23020 31272
rect 23072 31220 23078 31272
rect 23584 31260 23612 31288
rect 25424 31272 25452 31300
rect 25501 31297 25513 31331
rect 25547 31328 25559 31331
rect 25866 31328 25872 31340
rect 25547 31300 25872 31328
rect 25547 31297 25559 31300
rect 25501 31291 25559 31297
rect 25866 31288 25872 31300
rect 25924 31288 25930 31340
rect 26145 31331 26203 31337
rect 26145 31297 26157 31331
rect 26191 31297 26203 31331
rect 26145 31291 26203 31297
rect 24302 31260 24308 31272
rect 23584 31232 24308 31260
rect 24302 31220 24308 31232
rect 24360 31220 24366 31272
rect 24946 31220 24952 31272
rect 25004 31220 25010 31272
rect 25041 31263 25099 31269
rect 25041 31229 25053 31263
rect 25087 31229 25099 31263
rect 25041 31223 25099 31229
rect 20772 31096 21404 31124
rect 20772 31084 20778 31096
rect 22554 31084 22560 31136
rect 22612 31124 22618 31136
rect 23014 31124 23020 31136
rect 22612 31096 23020 31124
rect 22612 31084 22618 31096
rect 23014 31084 23020 31096
rect 23072 31084 23078 31136
rect 23198 31084 23204 31136
rect 23256 31124 23262 31136
rect 25056 31124 25084 31223
rect 25406 31220 25412 31272
rect 25464 31220 25470 31272
rect 25590 31220 25596 31272
rect 25648 31260 25654 31272
rect 26160 31260 26188 31291
rect 26234 31288 26240 31340
rect 26292 31288 26298 31340
rect 26878 31288 26884 31340
rect 26936 31328 26942 31340
rect 27356 31328 27384 31359
rect 28093 31350 28121 31436
rect 28828 31436 30748 31464
rect 28718 31396 28724 31408
rect 28552 31368 28724 31396
rect 28169 31353 28227 31359
rect 28169 31350 28181 31353
rect 26936 31300 27384 31328
rect 27433 31331 27491 31337
rect 26936 31288 26942 31300
rect 27433 31297 27445 31331
rect 27479 31328 27491 31331
rect 27522 31328 27528 31340
rect 27479 31300 27528 31328
rect 27479 31297 27491 31300
rect 27433 31291 27491 31297
rect 27522 31288 27528 31300
rect 27580 31288 27586 31340
rect 27617 31331 27675 31337
rect 27617 31297 27629 31331
rect 27663 31328 27675 31331
rect 27706 31328 27712 31340
rect 27663 31300 27712 31328
rect 27663 31297 27675 31300
rect 27617 31291 27675 31297
rect 27706 31288 27712 31300
rect 27764 31288 27770 31340
rect 27893 31331 27951 31337
rect 27893 31297 27905 31331
rect 27939 31297 27951 31331
rect 28093 31322 28181 31350
rect 28169 31319 28181 31322
rect 28215 31319 28227 31353
rect 28552 31337 28580 31368
rect 28718 31356 28724 31368
rect 28776 31356 28782 31408
rect 28169 31313 28227 31319
rect 28537 31331 28595 31337
rect 27893 31291 27951 31297
rect 28537 31297 28549 31331
rect 28583 31297 28595 31331
rect 28537 31291 28595 31297
rect 26418 31260 26424 31272
rect 25648 31232 26424 31260
rect 25648 31220 25654 31232
rect 26418 31220 26424 31232
rect 26476 31220 26482 31272
rect 26510 31220 26516 31272
rect 26568 31220 26574 31272
rect 26896 31260 26924 31288
rect 27908 31260 27936 31291
rect 28626 31288 28632 31340
rect 28684 31328 28690 31340
rect 28828 31337 28856 31436
rect 30742 31424 30748 31436
rect 30800 31464 30806 31476
rect 30837 31467 30895 31473
rect 30837 31464 30849 31467
rect 30800 31436 30849 31464
rect 30800 31424 30806 31436
rect 30837 31433 30849 31436
rect 30883 31433 30895 31467
rect 30837 31427 30895 31433
rect 31018 31424 31024 31476
rect 31076 31424 31082 31476
rect 32493 31467 32551 31473
rect 31128 31436 31984 31464
rect 29178 31356 29184 31408
rect 29236 31396 29242 31408
rect 31128 31396 31156 31436
rect 29236 31368 31156 31396
rect 31741 31399 31799 31405
rect 29236 31356 29242 31368
rect 31741 31365 31753 31399
rect 31787 31396 31799 31399
rect 31846 31396 31852 31408
rect 31787 31368 31852 31396
rect 31787 31365 31799 31368
rect 31741 31359 31799 31365
rect 31846 31356 31852 31368
rect 31904 31356 31910 31408
rect 31956 31405 31984 31436
rect 32493 31433 32505 31467
rect 32539 31464 32551 31467
rect 32674 31464 32680 31476
rect 32539 31436 32680 31464
rect 32539 31433 32551 31436
rect 32493 31427 32551 31433
rect 32674 31424 32680 31436
rect 32732 31464 32738 31476
rect 33045 31467 33103 31473
rect 33045 31464 33057 31467
rect 32732 31436 33057 31464
rect 32732 31424 32738 31436
rect 33045 31433 33057 31436
rect 33091 31433 33103 31467
rect 33045 31427 33103 31433
rect 31941 31399 31999 31405
rect 31941 31365 31953 31399
rect 31987 31396 31999 31399
rect 32398 31396 32404 31408
rect 31987 31368 32404 31396
rect 31987 31365 31999 31368
rect 31941 31359 31999 31365
rect 32398 31356 32404 31368
rect 32456 31356 32462 31408
rect 32766 31356 32772 31408
rect 32824 31396 32830 31408
rect 32953 31399 33011 31405
rect 32953 31396 32965 31399
rect 32824 31368 32965 31396
rect 32824 31356 32830 31368
rect 32953 31365 32965 31368
rect 32999 31365 33011 31399
rect 32953 31359 33011 31365
rect 28813 31331 28871 31337
rect 28813 31328 28825 31331
rect 28684 31300 28825 31328
rect 28684 31288 28690 31300
rect 28813 31297 28825 31300
rect 28859 31297 28871 31331
rect 28813 31291 28871 31297
rect 28902 31288 28908 31340
rect 28960 31328 28966 31340
rect 29089 31331 29147 31337
rect 29089 31328 29101 31331
rect 28960 31300 29101 31328
rect 28960 31288 28966 31300
rect 29089 31297 29101 31300
rect 29135 31297 29147 31331
rect 29089 31291 29147 31297
rect 29641 31331 29699 31337
rect 29641 31297 29653 31331
rect 29687 31297 29699 31331
rect 29641 31291 29699 31297
rect 26712 31232 26924 31260
rect 27724 31232 27936 31260
rect 29656 31260 29684 31291
rect 29822 31288 29828 31340
rect 29880 31288 29886 31340
rect 30190 31288 30196 31340
rect 30248 31288 30254 31340
rect 30374 31288 30380 31340
rect 30432 31288 30438 31340
rect 30466 31288 30472 31340
rect 30524 31288 30530 31340
rect 32582 31328 32588 31340
rect 30668 31300 32588 31328
rect 30558 31260 30564 31272
rect 29656 31232 30564 31260
rect 25222 31152 25228 31204
rect 25280 31192 25286 31204
rect 26712 31192 26740 31232
rect 25280 31164 26740 31192
rect 26789 31195 26847 31201
rect 25280 31152 25286 31164
rect 26789 31161 26801 31195
rect 26835 31161 26847 31195
rect 26789 31155 26847 31161
rect 23256 31096 25084 31124
rect 23256 31084 23262 31096
rect 25590 31084 25596 31136
rect 25648 31124 25654 31136
rect 26326 31124 26332 31136
rect 25648 31096 26332 31124
rect 25648 31084 25654 31096
rect 26326 31084 26332 31096
rect 26384 31084 26390 31136
rect 26510 31084 26516 31136
rect 26568 31124 26574 31136
rect 26804 31124 26832 31155
rect 27614 31152 27620 31204
rect 27672 31192 27678 31204
rect 27724 31192 27752 31232
rect 30558 31220 30564 31232
rect 30616 31260 30622 31272
rect 30668 31269 30696 31300
rect 32582 31288 32588 31300
rect 32640 31288 32646 31340
rect 32674 31288 32680 31340
rect 32732 31288 32738 31340
rect 33229 31331 33287 31337
rect 33229 31297 33241 31331
rect 33275 31328 33287 31331
rect 33318 31328 33324 31340
rect 33275 31300 33324 31328
rect 33275 31297 33287 31300
rect 33229 31291 33287 31297
rect 30653 31263 30711 31269
rect 30653 31260 30665 31263
rect 30616 31232 30665 31260
rect 30616 31220 30622 31232
rect 30653 31229 30665 31232
rect 30699 31229 30711 31263
rect 30653 31223 30711 31229
rect 30742 31220 30748 31272
rect 30800 31260 30806 31272
rect 31294 31260 31300 31272
rect 30800 31232 31300 31260
rect 30800 31220 30806 31232
rect 31294 31220 31300 31232
rect 31352 31220 31358 31272
rect 31588 31232 32444 31260
rect 27672 31164 27752 31192
rect 27801 31195 27859 31201
rect 27672 31152 27678 31164
rect 27801 31161 27813 31195
rect 27847 31192 27859 31195
rect 27890 31192 27896 31204
rect 27847 31164 27896 31192
rect 27847 31161 27859 31164
rect 27801 31155 27859 31161
rect 27890 31152 27896 31164
rect 27948 31152 27954 31204
rect 28074 31152 28080 31204
rect 28132 31152 28138 31204
rect 28169 31195 28227 31201
rect 28169 31161 28181 31195
rect 28215 31192 28227 31195
rect 28258 31192 28264 31204
rect 28215 31164 28264 31192
rect 28215 31161 28227 31164
rect 28169 31155 28227 31161
rect 28258 31152 28264 31164
rect 28316 31152 28322 31204
rect 30098 31192 30104 31204
rect 28460 31164 30104 31192
rect 26568 31096 26832 31124
rect 27197 31127 27255 31133
rect 26568 31084 26574 31096
rect 27197 31093 27209 31127
rect 27243 31124 27255 31127
rect 27338 31124 27344 31136
rect 27243 31096 27344 31124
rect 27243 31093 27255 31096
rect 27197 31087 27255 31093
rect 27338 31084 27344 31096
rect 27396 31084 27402 31136
rect 27430 31084 27436 31136
rect 27488 31124 27494 31136
rect 27525 31127 27583 31133
rect 27525 31124 27537 31127
rect 27488 31096 27537 31124
rect 27488 31084 27494 31096
rect 27525 31093 27537 31096
rect 27571 31124 27583 31127
rect 28460 31124 28488 31164
rect 30098 31152 30104 31164
rect 30156 31152 30162 31204
rect 30282 31152 30288 31204
rect 30340 31192 30346 31204
rect 31588 31201 31616 31232
rect 31389 31195 31447 31201
rect 31389 31192 31401 31195
rect 30340 31164 31401 31192
rect 30340 31152 30346 31164
rect 31389 31161 31401 31164
rect 31435 31161 31447 31195
rect 31389 31155 31447 31161
rect 31573 31195 31631 31201
rect 31573 31161 31585 31195
rect 31619 31161 31631 31195
rect 31573 31155 31631 31161
rect 32214 31152 32220 31204
rect 32272 31192 32278 31204
rect 32309 31195 32367 31201
rect 32309 31192 32321 31195
rect 32272 31164 32321 31192
rect 32272 31152 32278 31164
rect 32309 31161 32321 31164
rect 32355 31161 32367 31195
rect 32416 31192 32444 31232
rect 33244 31192 33272 31291
rect 33318 31288 33324 31300
rect 33376 31288 33382 31340
rect 32416 31164 33272 31192
rect 32309 31155 32367 31161
rect 27571 31096 28488 31124
rect 28905 31127 28963 31133
rect 27571 31093 27583 31096
rect 27525 31087 27583 31093
rect 28905 31093 28917 31127
rect 28951 31124 28963 31127
rect 28994 31124 29000 31136
rect 28951 31096 29000 31124
rect 28951 31093 28963 31096
rect 28905 31087 28963 31093
rect 28994 31084 29000 31096
rect 29052 31124 29058 31136
rect 30006 31124 30012 31136
rect 29052 31096 30012 31124
rect 29052 31084 29058 31096
rect 30006 31084 30012 31096
rect 30064 31084 30070 31136
rect 30190 31084 30196 31136
rect 30248 31124 30254 31136
rect 31021 31127 31079 31133
rect 31021 31124 31033 31127
rect 30248 31096 31033 31124
rect 30248 31084 30254 31096
rect 31021 31093 31033 31096
rect 31067 31093 31079 31127
rect 31021 31087 31079 31093
rect 31797 31127 31855 31133
rect 31797 31093 31809 31127
rect 31843 31124 31855 31127
rect 32232 31124 32260 31152
rect 31843 31096 32260 31124
rect 32861 31127 32919 31133
rect 31843 31093 31855 31096
rect 31797 31087 31855 31093
rect 32861 31093 32873 31127
rect 32907 31124 32919 31127
rect 33042 31124 33048 31136
rect 32907 31096 33048 31124
rect 32907 31093 32919 31096
rect 32861 31087 32919 31093
rect 33042 31084 33048 31096
rect 33100 31084 33106 31136
rect 33134 31084 33140 31136
rect 33192 31124 33198 31136
rect 33413 31127 33471 31133
rect 33413 31124 33425 31127
rect 33192 31096 33425 31124
rect 33192 31084 33198 31096
rect 33413 31093 33425 31096
rect 33459 31093 33471 31127
rect 33413 31087 33471 31093
rect 1104 31034 36432 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 36432 31034
rect 1104 30960 36432 30982
rect 4062 30880 4068 30932
rect 4120 30920 4126 30932
rect 4525 30923 4583 30929
rect 4120 30892 4292 30920
rect 4120 30880 4126 30892
rect 3142 30812 3148 30864
rect 3200 30852 3206 30864
rect 3200 30824 4200 30852
rect 3200 30812 3206 30824
rect 1489 30787 1547 30793
rect 1489 30753 1501 30787
rect 1535 30784 1547 30787
rect 3694 30784 3700 30796
rect 1535 30756 3700 30784
rect 1535 30753 1547 30756
rect 1489 30747 1547 30753
rect 3694 30744 3700 30756
rect 3752 30744 3758 30796
rect 3234 30676 3240 30728
rect 3292 30716 3298 30728
rect 4172 30725 4200 30824
rect 4264 30784 4292 30892
rect 4525 30889 4537 30923
rect 4571 30920 4583 30923
rect 4614 30920 4620 30932
rect 4571 30892 4620 30920
rect 4571 30889 4583 30892
rect 4525 30883 4583 30889
rect 4614 30880 4620 30892
rect 4672 30880 4678 30932
rect 4801 30923 4859 30929
rect 4801 30889 4813 30923
rect 4847 30920 4859 30923
rect 4890 30920 4896 30932
rect 4847 30892 4896 30920
rect 4847 30889 4859 30892
rect 4801 30883 4859 30889
rect 4890 30880 4896 30892
rect 4948 30880 4954 30932
rect 4982 30880 4988 30932
rect 5040 30920 5046 30932
rect 5261 30923 5319 30929
rect 5261 30920 5273 30923
rect 5040 30892 5273 30920
rect 5040 30880 5046 30892
rect 5261 30889 5273 30892
rect 5307 30920 5319 30923
rect 5718 30920 5724 30932
rect 5307 30892 5724 30920
rect 5307 30889 5319 30892
rect 5261 30883 5319 30889
rect 5718 30880 5724 30892
rect 5776 30880 5782 30932
rect 5902 30880 5908 30932
rect 5960 30920 5966 30932
rect 6825 30923 6883 30929
rect 6825 30920 6837 30923
rect 5960 30892 6837 30920
rect 5960 30880 5966 30892
rect 6825 30889 6837 30892
rect 6871 30889 6883 30923
rect 6825 30883 6883 30889
rect 7469 30923 7527 30929
rect 7469 30889 7481 30923
rect 7515 30920 7527 30923
rect 7558 30920 7564 30932
rect 7515 30892 7564 30920
rect 7515 30889 7527 30892
rect 7469 30883 7527 30889
rect 7558 30880 7564 30892
rect 7616 30880 7622 30932
rect 7834 30880 7840 30932
rect 7892 30920 7898 30932
rect 8389 30923 8447 30929
rect 8389 30920 8401 30923
rect 7892 30892 8401 30920
rect 7892 30880 7898 30892
rect 8389 30889 8401 30892
rect 8435 30889 8447 30923
rect 8389 30883 8447 30889
rect 8478 30880 8484 30932
rect 8536 30920 8542 30932
rect 8662 30920 8668 30932
rect 8536 30892 8668 30920
rect 8536 30880 8542 30892
rect 8662 30880 8668 30892
rect 8720 30920 8726 30932
rect 9214 30920 9220 30932
rect 8720 30892 9220 30920
rect 8720 30880 8726 30892
rect 9214 30880 9220 30892
rect 9272 30880 9278 30932
rect 11238 30920 11244 30932
rect 9416 30892 11244 30920
rect 6365 30855 6423 30861
rect 6365 30852 6377 30855
rect 4540 30824 6377 30852
rect 4430 30784 4436 30796
rect 4264 30756 4436 30784
rect 4264 30725 4292 30756
rect 4430 30744 4436 30756
rect 4488 30744 4494 30796
rect 4540 30725 4568 30824
rect 6365 30821 6377 30824
rect 6411 30821 6423 30855
rect 6365 30815 6423 30821
rect 7282 30812 7288 30864
rect 7340 30812 7346 30864
rect 5166 30744 5172 30796
rect 5224 30784 5230 30796
rect 6181 30787 6239 30793
rect 6181 30784 6193 30787
rect 5224 30756 6193 30784
rect 5224 30744 5230 30756
rect 6181 30753 6193 30756
rect 6227 30784 6239 30787
rect 7300 30784 7328 30812
rect 6227 30756 7328 30784
rect 7576 30784 7604 30880
rect 7742 30812 7748 30864
rect 7800 30852 7806 30864
rect 9416 30852 9444 30892
rect 11238 30880 11244 30892
rect 11296 30920 11302 30932
rect 11701 30923 11759 30929
rect 11701 30920 11713 30923
rect 11296 30892 11713 30920
rect 11296 30880 11302 30892
rect 11701 30889 11713 30892
rect 11747 30889 11759 30923
rect 14274 30920 14280 30932
rect 11701 30883 11759 30889
rect 11808 30892 14280 30920
rect 7800 30824 9444 30852
rect 7800 30812 7806 30824
rect 9674 30812 9680 30864
rect 9732 30852 9738 30864
rect 9769 30855 9827 30861
rect 9769 30852 9781 30855
rect 9732 30824 9781 30852
rect 9732 30812 9738 30824
rect 9769 30821 9781 30824
rect 9815 30821 9827 30855
rect 9769 30815 9827 30821
rect 10137 30855 10195 30861
rect 10137 30821 10149 30855
rect 10183 30821 10195 30855
rect 10137 30815 10195 30821
rect 10965 30855 11023 30861
rect 10965 30821 10977 30855
rect 11011 30852 11023 30855
rect 11146 30852 11152 30864
rect 11011 30824 11152 30852
rect 11011 30821 11023 30824
rect 10965 30815 11023 30821
rect 8021 30787 8079 30793
rect 7576 30756 7696 30784
rect 6227 30753 6239 30756
rect 6181 30747 6239 30753
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 3292 30688 3801 30716
rect 3292 30676 3298 30688
rect 3789 30685 3801 30688
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 3973 30719 4031 30725
rect 3973 30685 3985 30719
rect 4019 30716 4031 30719
rect 4157 30719 4215 30725
rect 4019 30688 4108 30716
rect 4019 30685 4031 30688
rect 3973 30679 4031 30685
rect 1762 30608 1768 30660
rect 1820 30608 1826 30660
rect 3050 30648 3056 30660
rect 2990 30620 3056 30648
rect 3050 30608 3056 30620
rect 3108 30608 3114 30660
rect 3513 30651 3571 30657
rect 3513 30617 3525 30651
rect 3559 30617 3571 30651
rect 3513 30611 3571 30617
rect 1302 30540 1308 30592
rect 1360 30580 1366 30592
rect 3528 30580 3556 30611
rect 1360 30552 3556 30580
rect 4080 30580 4108 30688
rect 4157 30685 4169 30719
rect 4203 30685 4215 30719
rect 4157 30679 4215 30685
rect 4249 30719 4307 30725
rect 4249 30685 4261 30719
rect 4295 30685 4307 30719
rect 4249 30679 4307 30685
rect 4341 30719 4399 30725
rect 4341 30685 4353 30719
rect 4387 30685 4399 30719
rect 4341 30679 4399 30685
rect 4525 30719 4583 30725
rect 4525 30685 4537 30719
rect 4571 30685 4583 30719
rect 4525 30679 4583 30685
rect 4356 30648 4384 30679
rect 4798 30676 4804 30728
rect 4856 30676 4862 30728
rect 5534 30716 5540 30728
rect 5092 30688 5540 30716
rect 4816 30648 4844 30676
rect 4356 30620 4844 30648
rect 4522 30580 4528 30592
rect 4080 30552 4528 30580
rect 1360 30540 1366 30552
rect 4522 30540 4528 30552
rect 4580 30540 4586 30592
rect 4632 30589 4660 30620
rect 4982 30608 4988 30660
rect 5040 30608 5046 30660
rect 5092 30589 5120 30688
rect 5534 30676 5540 30688
rect 5592 30716 5598 30728
rect 6641 30719 6699 30725
rect 6641 30716 6653 30719
rect 5592 30688 6653 30716
rect 5592 30676 5598 30688
rect 6641 30685 6653 30688
rect 6687 30685 6699 30719
rect 6641 30679 6699 30685
rect 6730 30676 6736 30728
rect 6788 30676 6794 30728
rect 6914 30676 6920 30728
rect 6972 30676 6978 30728
rect 7098 30676 7104 30728
rect 7156 30676 7162 30728
rect 7190 30676 7196 30728
rect 7248 30716 7254 30728
rect 7285 30719 7343 30725
rect 7285 30716 7297 30719
rect 7248 30688 7297 30716
rect 7248 30676 7254 30688
rect 7285 30685 7297 30688
rect 7331 30685 7343 30719
rect 7285 30679 7343 30685
rect 5445 30651 5503 30657
rect 5445 30617 5457 30651
rect 5491 30648 5503 30651
rect 5718 30648 5724 30660
rect 5491 30620 5724 30648
rect 5491 30617 5503 30620
rect 5445 30611 5503 30617
rect 5718 30608 5724 30620
rect 5776 30608 5782 30660
rect 5905 30651 5963 30657
rect 5905 30617 5917 30651
rect 5951 30648 5963 30651
rect 6086 30648 6092 30660
rect 5951 30620 6092 30648
rect 5951 30617 5963 30620
rect 5905 30611 5963 30617
rect 6086 30608 6092 30620
rect 6144 30608 6150 30660
rect 6365 30651 6423 30657
rect 6365 30617 6377 30651
rect 6411 30648 6423 30651
rect 6454 30648 6460 30660
rect 6411 30620 6460 30648
rect 6411 30617 6423 30620
rect 6365 30611 6423 30617
rect 6454 30608 6460 30620
rect 6512 30608 6518 30660
rect 4617 30583 4675 30589
rect 4617 30549 4629 30583
rect 4663 30549 4675 30583
rect 4617 30543 4675 30549
rect 4785 30583 4843 30589
rect 4785 30549 4797 30583
rect 4831 30580 4843 30583
rect 5077 30583 5135 30589
rect 5077 30580 5089 30583
rect 4831 30552 5089 30580
rect 4831 30549 4843 30552
rect 4785 30543 4843 30549
rect 5077 30549 5089 30552
rect 5123 30549 5135 30583
rect 5077 30543 5135 30549
rect 5245 30583 5303 30589
rect 5245 30549 5257 30583
rect 5291 30580 5303 30583
rect 5350 30580 5356 30592
rect 5291 30552 5356 30580
rect 5291 30549 5303 30552
rect 5245 30543 5303 30549
rect 5350 30540 5356 30552
rect 5408 30540 5414 30592
rect 5534 30540 5540 30592
rect 5592 30540 5598 30592
rect 5994 30540 6000 30592
rect 6052 30540 6058 30592
rect 6546 30540 6552 30592
rect 6604 30540 6610 30592
rect 7300 30580 7328 30679
rect 7558 30676 7564 30728
rect 7616 30676 7622 30728
rect 7668 30648 7696 30756
rect 8021 30753 8033 30787
rect 8067 30784 8079 30787
rect 8067 30756 8432 30784
rect 8067 30753 8079 30756
rect 8021 30747 8079 30753
rect 7926 30676 7932 30728
rect 7984 30676 7990 30728
rect 8110 30676 8116 30728
rect 8168 30676 8174 30728
rect 8404 30725 8432 30756
rect 8662 30744 8668 30796
rect 8720 30784 8726 30796
rect 9306 30784 9312 30796
rect 8720 30756 9312 30784
rect 8720 30744 8726 30756
rect 9306 30744 9312 30756
rect 9364 30744 9370 30796
rect 9493 30787 9551 30793
rect 9493 30753 9505 30787
rect 9539 30784 9551 30787
rect 10152 30784 10180 30815
rect 11146 30812 11152 30824
rect 11204 30812 11210 30864
rect 9539 30756 10180 30784
rect 9539 30753 9551 30756
rect 9493 30747 9551 30753
rect 10226 30744 10232 30796
rect 10284 30784 10290 30796
rect 10689 30787 10747 30793
rect 10689 30784 10701 30787
rect 10284 30756 10701 30784
rect 10284 30744 10290 30756
rect 10689 30753 10701 30756
rect 10735 30753 10747 30787
rect 10689 30747 10747 30753
rect 11422 30744 11428 30796
rect 11480 30744 11486 30796
rect 8205 30719 8263 30725
rect 8205 30685 8217 30719
rect 8251 30685 8263 30719
rect 8205 30679 8263 30685
rect 8389 30719 8447 30725
rect 8389 30685 8401 30719
rect 8435 30685 8447 30719
rect 8389 30679 8447 30685
rect 9401 30719 9459 30725
rect 9401 30685 9413 30719
rect 9447 30716 9459 30719
rect 9582 30716 9588 30728
rect 9447 30688 9588 30716
rect 9447 30685 9459 30688
rect 9401 30679 9459 30685
rect 8220 30648 8248 30679
rect 9582 30676 9588 30688
rect 9640 30676 9646 30728
rect 10410 30676 10416 30728
rect 10468 30716 10474 30728
rect 11808 30725 11836 30892
rect 14274 30880 14280 30892
rect 14332 30880 14338 30932
rect 14384 30892 17540 30920
rect 14384 30852 14412 30892
rect 13740 30824 14412 30852
rect 14829 30855 14887 30861
rect 11333 30719 11391 30725
rect 11333 30716 11345 30719
rect 10468 30688 11345 30716
rect 10468 30676 10474 30688
rect 11333 30685 11345 30688
rect 11379 30685 11391 30719
rect 11333 30679 11391 30685
rect 11793 30719 11851 30725
rect 11793 30685 11805 30719
rect 11839 30685 11851 30719
rect 11793 30679 11851 30685
rect 11974 30676 11980 30728
rect 12032 30716 12038 30728
rect 12342 30716 12348 30728
rect 12032 30688 12348 30716
rect 12032 30676 12038 30688
rect 12342 30676 12348 30688
rect 12400 30716 12406 30728
rect 13541 30719 13599 30725
rect 13541 30716 13553 30719
rect 12400 30688 13553 30716
rect 12400 30676 12406 30688
rect 13541 30685 13553 30688
rect 13587 30685 13599 30719
rect 13541 30679 13599 30685
rect 7668 30620 8248 30648
rect 9490 30608 9496 30660
rect 9548 30648 9554 30660
rect 13740 30648 13768 30824
rect 14829 30821 14841 30855
rect 14875 30852 14887 30855
rect 15010 30852 15016 30864
rect 14875 30824 15016 30852
rect 14875 30821 14887 30824
rect 14829 30815 14887 30821
rect 13817 30787 13875 30793
rect 13817 30753 13829 30787
rect 13863 30753 13875 30787
rect 13817 30747 13875 30753
rect 13832 30716 13860 30747
rect 14844 30728 14872 30815
rect 15010 30812 15016 30824
rect 15068 30812 15074 30864
rect 15286 30812 15292 30864
rect 15344 30852 15350 30864
rect 15930 30852 15936 30864
rect 15344 30824 15936 30852
rect 15344 30812 15350 30824
rect 15930 30812 15936 30824
rect 15988 30852 15994 30864
rect 16485 30855 16543 30861
rect 15988 30824 16436 30852
rect 15988 30812 15994 30824
rect 16206 30744 16212 30796
rect 16264 30744 16270 30796
rect 16408 30784 16436 30824
rect 16485 30821 16497 30855
rect 16531 30852 16543 30855
rect 17512 30852 17540 30892
rect 17862 30880 17868 30932
rect 17920 30920 17926 30932
rect 18049 30923 18107 30929
rect 18049 30920 18061 30923
rect 17920 30892 18061 30920
rect 17920 30880 17926 30892
rect 18049 30889 18061 30892
rect 18095 30889 18107 30923
rect 18049 30883 18107 30889
rect 21358 30880 21364 30932
rect 21416 30880 21422 30932
rect 21726 30880 21732 30932
rect 21784 30920 21790 30932
rect 21784 30892 22784 30920
rect 21784 30880 21790 30892
rect 19337 30855 19395 30861
rect 19337 30852 19349 30855
rect 16531 30824 16712 30852
rect 17512 30824 19349 30852
rect 16531 30821 16543 30824
rect 16485 30815 16543 30821
rect 16408 30756 16620 30784
rect 14277 30719 14335 30725
rect 14277 30716 14289 30719
rect 13832 30688 14289 30716
rect 14277 30685 14289 30688
rect 14323 30716 14335 30719
rect 14826 30716 14832 30728
rect 14323 30688 14832 30716
rect 14323 30685 14335 30688
rect 14277 30679 14335 30685
rect 14826 30676 14832 30688
rect 14884 30676 14890 30728
rect 15746 30676 15752 30728
rect 15804 30716 15810 30728
rect 15841 30719 15899 30725
rect 15841 30716 15853 30719
rect 15804 30688 15853 30716
rect 15804 30676 15810 30688
rect 15841 30685 15853 30688
rect 15887 30685 15899 30719
rect 15841 30679 15899 30685
rect 15934 30719 15992 30725
rect 15934 30685 15946 30719
rect 15980 30685 15992 30719
rect 15934 30679 15992 30685
rect 9548 30620 13768 30648
rect 9548 30608 9554 30620
rect 14090 30608 14096 30660
rect 14148 30608 14154 30660
rect 14642 30608 14648 30660
rect 14700 30608 14706 30660
rect 15654 30608 15660 30660
rect 15712 30648 15718 30660
rect 15948 30648 15976 30679
rect 16114 30676 16120 30728
rect 16172 30676 16178 30728
rect 16224 30716 16252 30744
rect 16592 30725 16620 30756
rect 16684 30725 16712 30824
rect 19337 30821 19349 30824
rect 19383 30821 19395 30855
rect 20990 30852 20996 30864
rect 19337 30815 19395 30821
rect 19444 30824 20996 30852
rect 19444 30784 19472 30824
rect 20990 30812 20996 30824
rect 21048 30812 21054 30864
rect 21177 30855 21235 30861
rect 21177 30821 21189 30855
rect 21223 30852 21235 30855
rect 21910 30852 21916 30864
rect 21223 30824 21916 30852
rect 21223 30821 21235 30824
rect 21177 30815 21235 30821
rect 21910 30812 21916 30824
rect 21968 30852 21974 30864
rect 21968 30824 22508 30852
rect 21968 30812 21974 30824
rect 20162 30784 20168 30796
rect 18984 30756 19472 30784
rect 19628 30756 20168 30784
rect 16306 30719 16364 30725
rect 16306 30716 16318 30719
rect 16224 30688 16318 30716
rect 16306 30685 16318 30688
rect 16352 30685 16364 30719
rect 16306 30679 16364 30685
rect 16577 30719 16635 30725
rect 16577 30685 16589 30719
rect 16623 30685 16635 30719
rect 16577 30679 16635 30685
rect 16669 30719 16727 30725
rect 16669 30685 16681 30719
rect 16715 30685 16727 30719
rect 16669 30679 16727 30685
rect 16853 30719 16911 30725
rect 16853 30685 16865 30719
rect 16899 30685 16911 30719
rect 16853 30679 16911 30685
rect 16945 30719 17003 30725
rect 16945 30685 16957 30719
rect 16991 30716 17003 30719
rect 17954 30716 17960 30728
rect 16991 30688 17960 30716
rect 16991 30685 17003 30688
rect 16945 30679 17003 30685
rect 15712 30620 15976 30648
rect 15712 30608 15718 30620
rect 16206 30608 16212 30660
rect 16264 30608 16270 30660
rect 16868 30648 16896 30679
rect 17954 30676 17960 30688
rect 18012 30716 18018 30728
rect 18874 30716 18880 30728
rect 18012 30688 18880 30716
rect 18012 30676 18018 30688
rect 18874 30676 18880 30688
rect 18932 30676 18938 30728
rect 18984 30725 19012 30756
rect 18969 30719 19027 30725
rect 18969 30685 18981 30719
rect 19015 30685 19027 30719
rect 18969 30679 19027 30685
rect 16868 30620 17264 30648
rect 17236 30592 17264 30620
rect 17678 30608 17684 30660
rect 17736 30608 17742 30660
rect 17862 30608 17868 30660
rect 17920 30608 17926 30660
rect 18984 30648 19012 30679
rect 19334 30676 19340 30728
rect 19392 30716 19398 30728
rect 19628 30725 19656 30756
rect 20162 30744 20168 30756
rect 20220 30744 20226 30796
rect 20898 30744 20904 30796
rect 20956 30784 20962 30796
rect 20956 30756 22232 30784
rect 20956 30744 20962 30756
rect 19521 30719 19579 30725
rect 19521 30716 19533 30719
rect 19392 30688 19533 30716
rect 19392 30676 19398 30688
rect 19521 30685 19533 30688
rect 19567 30685 19579 30719
rect 19521 30679 19579 30685
rect 19613 30719 19671 30725
rect 19613 30685 19625 30719
rect 19659 30685 19671 30719
rect 19613 30679 19671 30685
rect 19794 30676 19800 30728
rect 19852 30676 19858 30728
rect 19889 30719 19947 30725
rect 19889 30685 19901 30719
rect 19935 30716 19947 30719
rect 20254 30716 20260 30728
rect 19935 30688 20260 30716
rect 19935 30685 19947 30688
rect 19889 30679 19947 30685
rect 17972 30620 19012 30648
rect 7745 30583 7803 30589
rect 7745 30580 7757 30583
rect 7300 30552 7757 30580
rect 7745 30549 7757 30552
rect 7791 30580 7803 30583
rect 8110 30580 8116 30592
rect 7791 30552 8116 30580
rect 7791 30549 7803 30552
rect 7745 30543 7803 30549
rect 8110 30540 8116 30552
rect 8168 30540 8174 30592
rect 10502 30540 10508 30592
rect 10560 30540 10566 30592
rect 10597 30583 10655 30589
rect 10597 30549 10609 30583
rect 10643 30580 10655 30583
rect 10870 30580 10876 30592
rect 10643 30552 10876 30580
rect 10643 30549 10655 30552
rect 10597 30543 10655 30549
rect 10870 30540 10876 30552
rect 10928 30540 10934 30592
rect 13170 30540 13176 30592
rect 13228 30540 13234 30592
rect 13262 30540 13268 30592
rect 13320 30580 13326 30592
rect 13633 30583 13691 30589
rect 13633 30580 13645 30583
rect 13320 30552 13645 30580
rect 13320 30540 13326 30552
rect 13633 30549 13645 30552
rect 13679 30549 13691 30583
rect 13633 30543 13691 30549
rect 14461 30583 14519 30589
rect 14461 30549 14473 30583
rect 14507 30580 14519 30583
rect 15194 30580 15200 30592
rect 14507 30552 15200 30580
rect 14507 30549 14519 30552
rect 14461 30543 14519 30549
rect 15194 30540 15200 30552
rect 15252 30540 15258 30592
rect 17126 30540 17132 30592
rect 17184 30540 17190 30592
rect 17218 30540 17224 30592
rect 17276 30580 17282 30592
rect 17972 30580 18000 30620
rect 19242 30608 19248 30660
rect 19300 30648 19306 30660
rect 19904 30648 19932 30679
rect 20254 30676 20260 30688
rect 20312 30676 20318 30728
rect 20714 30676 20720 30728
rect 20772 30716 20778 30728
rect 21726 30716 21732 30728
rect 20772 30688 21732 30716
rect 20772 30676 20778 30688
rect 21726 30676 21732 30688
rect 21784 30676 21790 30728
rect 22002 30676 22008 30728
rect 22060 30676 22066 30728
rect 22204 30725 22232 30756
rect 22480 30725 22508 30824
rect 22756 30784 22784 30892
rect 22830 30880 22836 30932
rect 22888 30920 22894 30932
rect 24581 30923 24639 30929
rect 24581 30920 24593 30923
rect 22888 30892 24593 30920
rect 22888 30880 22894 30892
rect 24581 30889 24593 30892
rect 24627 30889 24639 30923
rect 24581 30883 24639 30889
rect 25866 30880 25872 30932
rect 25924 30920 25930 30932
rect 27433 30923 27491 30929
rect 25924 30892 27016 30920
rect 25924 30880 25930 30892
rect 23014 30812 23020 30864
rect 23072 30852 23078 30864
rect 23201 30855 23259 30861
rect 23201 30852 23213 30855
rect 23072 30824 23213 30852
rect 23072 30812 23078 30824
rect 23201 30821 23213 30824
rect 23247 30821 23259 30855
rect 23201 30815 23259 30821
rect 23382 30812 23388 30864
rect 23440 30852 23446 30864
rect 26881 30855 26939 30861
rect 23440 30824 23888 30852
rect 23440 30812 23446 30824
rect 22756 30756 23428 30784
rect 22756 30725 22784 30756
rect 22189 30719 22247 30725
rect 22189 30685 22201 30719
rect 22235 30685 22247 30719
rect 22189 30679 22247 30685
rect 22465 30719 22523 30725
rect 22465 30685 22477 30719
rect 22511 30685 22523 30719
rect 22465 30679 22523 30685
rect 22741 30719 22799 30725
rect 22741 30685 22753 30719
rect 22787 30685 22799 30719
rect 22741 30679 22799 30685
rect 22833 30719 22891 30725
rect 22833 30685 22845 30719
rect 22879 30716 22891 30719
rect 23198 30716 23204 30728
rect 22879 30688 23204 30716
rect 22879 30685 22891 30688
rect 22833 30679 22891 30685
rect 19300 30620 19932 30648
rect 19300 30608 19306 30620
rect 20622 30608 20628 30660
rect 20680 30648 20686 30660
rect 20680 30620 22094 30648
rect 20680 30608 20686 30620
rect 17276 30552 18000 30580
rect 17276 30540 17282 30552
rect 18874 30540 18880 30592
rect 18932 30540 18938 30592
rect 19150 30540 19156 30592
rect 19208 30580 19214 30592
rect 21358 30580 21364 30592
rect 19208 30552 21364 30580
rect 19208 30540 19214 30552
rect 21358 30540 21364 30552
rect 21416 30540 21422 30592
rect 22066 30580 22094 30620
rect 23032 30580 23060 30688
rect 23198 30676 23204 30688
rect 23256 30676 23262 30728
rect 23400 30725 23428 30756
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30685 23443 30719
rect 23385 30679 23443 30685
rect 23474 30676 23480 30728
rect 23532 30716 23538 30728
rect 23860 30725 23888 30824
rect 26881 30821 26893 30855
rect 26927 30821 26939 30855
rect 26988 30852 27016 30892
rect 27433 30889 27445 30923
rect 27479 30920 27491 30923
rect 27614 30920 27620 30932
rect 27479 30892 27620 30920
rect 27479 30889 27491 30892
rect 27433 30883 27491 30889
rect 27614 30880 27620 30892
rect 27672 30880 27678 30932
rect 27709 30923 27767 30929
rect 27709 30889 27721 30923
rect 27755 30920 27767 30923
rect 28074 30920 28080 30932
rect 27755 30892 28080 30920
rect 27755 30889 27767 30892
rect 27709 30883 27767 30889
rect 28074 30880 28080 30892
rect 28132 30920 28138 30932
rect 30745 30923 30803 30929
rect 28132 30892 28856 30920
rect 28132 30880 28138 30892
rect 28169 30855 28227 30861
rect 28169 30852 28181 30855
rect 26988 30824 28181 30852
rect 26881 30815 26939 30821
rect 28169 30821 28181 30824
rect 28215 30821 28227 30855
rect 28169 30815 28227 30821
rect 26896 30784 26924 30815
rect 27522 30784 27528 30796
rect 24596 30756 27528 30784
rect 23569 30719 23627 30725
rect 23569 30716 23581 30719
rect 23532 30688 23581 30716
rect 23532 30676 23538 30688
rect 23569 30685 23581 30688
rect 23615 30685 23627 30719
rect 23569 30679 23627 30685
rect 23845 30719 23903 30725
rect 23845 30685 23857 30719
rect 23891 30685 23903 30719
rect 23845 30679 23903 30685
rect 23934 30676 23940 30728
rect 23992 30716 23998 30728
rect 24596 30725 24624 30756
rect 27522 30744 27528 30756
rect 27580 30744 27586 30796
rect 28534 30784 28540 30796
rect 27816 30756 28540 30784
rect 24397 30719 24455 30725
rect 24397 30716 24409 30719
rect 23992 30688 24409 30716
rect 23992 30676 23998 30688
rect 24397 30685 24409 30688
rect 24443 30685 24455 30719
rect 24397 30679 24455 30685
rect 24581 30719 24639 30725
rect 24581 30685 24593 30719
rect 24627 30685 24639 30719
rect 24581 30679 24639 30685
rect 24854 30676 24860 30728
rect 24912 30716 24918 30728
rect 25038 30716 25044 30728
rect 24912 30688 25044 30716
rect 24912 30676 24918 30688
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 26602 30676 26608 30728
rect 26660 30676 26666 30728
rect 27062 30676 27068 30728
rect 27120 30676 27126 30728
rect 27249 30719 27307 30725
rect 27249 30685 27261 30719
rect 27295 30716 27307 30719
rect 27430 30716 27436 30728
rect 27295 30688 27436 30716
rect 27295 30685 27307 30688
rect 27249 30679 27307 30685
rect 27430 30676 27436 30688
rect 27488 30676 27494 30728
rect 27614 30676 27620 30728
rect 27672 30676 27678 30728
rect 27816 30725 27844 30756
rect 28534 30744 28540 30756
rect 28592 30744 28598 30796
rect 27801 30719 27859 30725
rect 27801 30685 27813 30719
rect 27847 30685 27859 30719
rect 27801 30679 27859 30685
rect 27890 30676 27896 30728
rect 27948 30676 27954 30728
rect 28074 30676 28080 30728
rect 28132 30676 28138 30728
rect 28169 30719 28227 30725
rect 28169 30685 28181 30719
rect 28215 30685 28227 30719
rect 28169 30679 28227 30685
rect 28353 30719 28411 30725
rect 28353 30685 28365 30719
rect 28399 30716 28411 30719
rect 28718 30716 28724 30728
rect 28399 30688 28724 30716
rect 28399 30685 28411 30688
rect 28353 30679 28411 30685
rect 24029 30651 24087 30657
rect 24029 30617 24041 30651
rect 24075 30617 24087 30651
rect 24029 30611 24087 30617
rect 22066 30552 23060 30580
rect 23198 30540 23204 30592
rect 23256 30580 23262 30592
rect 23477 30583 23535 30589
rect 23477 30580 23489 30583
rect 23256 30552 23489 30580
rect 23256 30540 23262 30552
rect 23477 30549 23489 30552
rect 23523 30549 23535 30583
rect 23477 30543 23535 30549
rect 23566 30540 23572 30592
rect 23624 30580 23630 30592
rect 24044 30580 24072 30611
rect 24210 30608 24216 30660
rect 24268 30608 24274 30660
rect 24302 30608 24308 30660
rect 24360 30648 24366 30660
rect 24360 30620 25162 30648
rect 24360 30608 24366 30620
rect 26326 30608 26332 30660
rect 26384 30608 26390 30660
rect 26418 30608 26424 30660
rect 26476 30648 26482 30660
rect 27525 30651 27583 30657
rect 27525 30648 27537 30651
rect 26476 30620 27537 30648
rect 26476 30608 26482 30620
rect 27525 30617 27537 30620
rect 27571 30648 27583 30651
rect 27706 30648 27712 30660
rect 27571 30620 27712 30648
rect 27571 30617 27583 30620
rect 27525 30611 27583 30617
rect 27706 30608 27712 30620
rect 27764 30608 27770 30660
rect 27908 30648 27936 30676
rect 28184 30648 28212 30679
rect 28718 30676 28724 30688
rect 28776 30676 28782 30728
rect 27908 30620 28212 30648
rect 28626 30608 28632 30660
rect 28684 30608 28690 30660
rect 28828 30648 28856 30892
rect 30745 30889 30757 30923
rect 30791 30889 30803 30923
rect 30745 30883 30803 30889
rect 31205 30923 31263 30929
rect 31205 30889 31217 30923
rect 31251 30920 31263 30923
rect 31478 30920 31484 30932
rect 31251 30892 31484 30920
rect 31251 30889 31263 30892
rect 31205 30883 31263 30889
rect 28902 30812 28908 30864
rect 28960 30852 28966 30864
rect 28960 30824 29132 30852
rect 28960 30812 28966 30824
rect 28994 30744 29000 30796
rect 29052 30744 29058 30796
rect 28905 30719 28963 30725
rect 28905 30685 28917 30719
rect 28951 30716 28963 30719
rect 29012 30716 29040 30744
rect 29104 30725 29132 30824
rect 30466 30812 30472 30864
rect 30524 30852 30530 30864
rect 30760 30852 30788 30883
rect 31478 30880 31484 30892
rect 31536 30880 31542 30932
rect 31662 30852 31668 30864
rect 30524 30824 31668 30852
rect 30524 30812 30530 30824
rect 31662 30812 31668 30824
rect 31720 30812 31726 30864
rect 30282 30744 30288 30796
rect 30340 30784 30346 30796
rect 30340 30756 31340 30784
rect 30340 30744 30346 30756
rect 28951 30688 29040 30716
rect 29089 30719 29147 30725
rect 28951 30685 28963 30688
rect 28905 30679 28963 30685
rect 29089 30685 29101 30719
rect 29135 30685 29147 30719
rect 29089 30679 29147 30685
rect 29362 30676 29368 30728
rect 29420 30716 29426 30728
rect 29917 30719 29975 30725
rect 29420 30688 29868 30716
rect 29420 30676 29426 30688
rect 29733 30651 29791 30657
rect 29733 30648 29745 30651
rect 28828 30620 29745 30648
rect 29733 30617 29745 30620
rect 29779 30617 29791 30651
rect 29840 30648 29868 30688
rect 29917 30685 29929 30719
rect 29963 30716 29975 30719
rect 30006 30716 30012 30728
rect 29963 30688 30012 30716
rect 29963 30685 29975 30688
rect 29917 30679 29975 30685
rect 30006 30676 30012 30688
rect 30064 30676 30070 30728
rect 30190 30676 30196 30728
rect 30248 30716 30254 30728
rect 31312 30725 31340 30756
rect 31113 30719 31171 30725
rect 31113 30716 31125 30719
rect 30248 30688 31125 30716
rect 30248 30676 30254 30688
rect 31113 30685 31125 30688
rect 31159 30685 31171 30719
rect 31113 30679 31171 30685
rect 31297 30719 31355 30725
rect 31297 30685 31309 30719
rect 31343 30716 31355 30719
rect 36262 30716 36268 30728
rect 31343 30688 36268 30716
rect 31343 30685 31355 30688
rect 31297 30679 31355 30685
rect 36262 30676 36268 30688
rect 36320 30676 36326 30728
rect 30561 30651 30619 30657
rect 30561 30648 30573 30651
rect 29840 30620 30573 30648
rect 29733 30611 29791 30617
rect 30561 30617 30573 30620
rect 30607 30617 30619 30651
rect 30561 30611 30619 30617
rect 30742 30608 30748 30660
rect 30800 30608 30806 30660
rect 24762 30580 24768 30592
rect 23624 30552 24768 30580
rect 23624 30540 23630 30552
rect 24762 30540 24768 30552
rect 24820 30540 24826 30592
rect 24854 30540 24860 30592
rect 24912 30540 24918 30592
rect 25406 30540 25412 30592
rect 25464 30580 25470 30592
rect 26142 30580 26148 30592
rect 25464 30552 26148 30580
rect 25464 30540 25470 30552
rect 26142 30540 26148 30552
rect 26200 30540 26206 30592
rect 27614 30540 27620 30592
rect 27672 30580 27678 30592
rect 27985 30583 28043 30589
rect 27985 30580 27997 30583
rect 27672 30552 27997 30580
rect 27672 30540 27678 30552
rect 27985 30549 27997 30552
rect 28031 30549 28043 30583
rect 27985 30543 28043 30549
rect 28166 30540 28172 30592
rect 28224 30580 28230 30592
rect 28810 30580 28816 30592
rect 28224 30552 28816 30580
rect 28224 30540 28230 30552
rect 28810 30540 28816 30552
rect 28868 30540 28874 30592
rect 29546 30540 29552 30592
rect 29604 30540 29610 30592
rect 30929 30583 30987 30589
rect 30929 30549 30941 30583
rect 30975 30580 30987 30583
rect 31294 30580 31300 30592
rect 30975 30552 31300 30580
rect 30975 30549 30987 30552
rect 30929 30543 30987 30549
rect 31294 30540 31300 30552
rect 31352 30540 31358 30592
rect 1104 30490 36432 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 36432 30490
rect 1104 30416 36432 30438
rect 3050 30336 3056 30388
rect 3108 30376 3114 30388
rect 5718 30376 5724 30388
rect 3108 30348 5304 30376
rect 3108 30336 3114 30348
rect 3068 30308 3096 30336
rect 5276 30320 5304 30348
rect 5368 30348 5724 30376
rect 5258 30308 5264 30320
rect 2898 30280 3096 30308
rect 5198 30280 5264 30308
rect 5258 30268 5264 30280
rect 5316 30268 5322 30320
rect 3605 30243 3663 30249
rect 3605 30209 3617 30243
rect 3651 30240 3663 30243
rect 3694 30240 3700 30252
rect 3651 30212 3700 30240
rect 3651 30209 3663 30212
rect 3605 30203 3663 30209
rect 3694 30200 3700 30212
rect 3752 30200 3758 30252
rect 1302 30132 1308 30184
rect 1360 30172 1366 30184
rect 1581 30175 1639 30181
rect 1581 30172 1593 30175
rect 1360 30144 1593 30172
rect 1360 30132 1366 30144
rect 1581 30141 1593 30144
rect 1627 30141 1639 30175
rect 1581 30135 1639 30141
rect 3329 30175 3387 30181
rect 3329 30141 3341 30175
rect 3375 30172 3387 30175
rect 3375 30144 3648 30172
rect 3375 30141 3387 30144
rect 3329 30135 3387 30141
rect 3620 30116 3648 30144
rect 3970 30132 3976 30184
rect 4028 30132 4034 30184
rect 5258 30132 5264 30184
rect 5316 30172 5322 30184
rect 5368 30172 5396 30348
rect 5718 30336 5724 30348
rect 5776 30376 5782 30388
rect 5776 30348 5948 30376
rect 5776 30336 5782 30348
rect 5920 30308 5948 30348
rect 5994 30336 6000 30388
rect 6052 30376 6058 30388
rect 6089 30379 6147 30385
rect 6089 30376 6101 30379
rect 6052 30348 6101 30376
rect 6052 30336 6058 30348
rect 6089 30345 6101 30348
rect 6135 30345 6147 30379
rect 6089 30339 6147 30345
rect 6270 30336 6276 30388
rect 6328 30376 6334 30388
rect 10134 30376 10140 30388
rect 6328 30348 10140 30376
rect 6328 30336 6334 30348
rect 10134 30336 10140 30348
rect 10192 30336 10198 30388
rect 10686 30336 10692 30388
rect 10744 30385 10750 30388
rect 10744 30379 10763 30385
rect 10751 30345 10763 30379
rect 10744 30339 10763 30345
rect 10744 30336 10750 30339
rect 10870 30336 10876 30388
rect 10928 30336 10934 30388
rect 11422 30336 11428 30388
rect 11480 30376 11486 30388
rect 11609 30379 11667 30385
rect 11609 30376 11621 30379
rect 11480 30348 11621 30376
rect 11480 30336 11486 30348
rect 11609 30345 11621 30348
rect 11655 30345 11667 30379
rect 11609 30339 11667 30345
rect 14090 30336 14096 30388
rect 14148 30336 14154 30388
rect 14642 30336 14648 30388
rect 14700 30376 14706 30388
rect 19058 30376 19064 30388
rect 14700 30348 19064 30376
rect 14700 30336 14706 30348
rect 19058 30336 19064 30348
rect 19116 30336 19122 30388
rect 19610 30376 19616 30388
rect 19358 30348 19616 30376
rect 5920 30280 8800 30308
rect 5718 30200 5724 30252
rect 5776 30240 5782 30252
rect 6730 30240 6736 30252
rect 5776 30212 6736 30240
rect 5776 30200 5782 30212
rect 6730 30200 6736 30212
rect 6788 30200 6794 30252
rect 7282 30200 7288 30252
rect 7340 30240 7346 30252
rect 7745 30243 7803 30249
rect 7745 30240 7757 30243
rect 7340 30212 7757 30240
rect 7340 30200 7346 30212
rect 7745 30209 7757 30212
rect 7791 30209 7803 30243
rect 7745 30203 7803 30209
rect 5316 30144 5396 30172
rect 5316 30132 5322 30144
rect 5810 30132 5816 30184
rect 5868 30132 5874 30184
rect 7006 30132 7012 30184
rect 7064 30172 7070 30184
rect 7469 30175 7527 30181
rect 7469 30172 7481 30175
rect 7064 30144 7481 30172
rect 7064 30132 7070 30144
rect 7469 30141 7481 30144
rect 7515 30141 7527 30175
rect 7469 30135 7527 30141
rect 7650 30132 7656 30184
rect 7708 30132 7714 30184
rect 8570 30132 8576 30184
rect 8628 30172 8634 30184
rect 8665 30175 8723 30181
rect 8665 30172 8677 30175
rect 8628 30144 8677 30172
rect 8628 30132 8634 30144
rect 8665 30141 8677 30144
rect 8711 30141 8723 30175
rect 8772 30172 8800 30280
rect 9122 30268 9128 30320
rect 9180 30268 9186 30320
rect 10045 30311 10103 30317
rect 10045 30277 10057 30311
rect 10091 30308 10103 30311
rect 10226 30308 10232 30320
rect 10091 30280 10232 30308
rect 10091 30277 10103 30280
rect 10045 30271 10103 30277
rect 10226 30268 10232 30280
rect 10284 30268 10290 30320
rect 10505 30311 10563 30317
rect 10505 30308 10517 30311
rect 10336 30280 10517 30308
rect 8846 30200 8852 30252
rect 8904 30200 8910 30252
rect 8938 30200 8944 30252
rect 8996 30240 9002 30252
rect 9217 30243 9275 30249
rect 9217 30240 9229 30243
rect 8996 30212 9229 30240
rect 8996 30200 9002 30212
rect 9217 30209 9229 30212
rect 9263 30209 9275 30243
rect 9217 30203 9275 30209
rect 10137 30243 10195 30249
rect 10137 30209 10149 30243
rect 10183 30240 10195 30243
rect 10336 30240 10364 30280
rect 10505 30277 10517 30280
rect 10551 30308 10563 30311
rect 10594 30308 10600 30320
rect 10551 30280 10600 30308
rect 10551 30277 10563 30280
rect 10505 30271 10563 30277
rect 10594 30268 10600 30280
rect 10652 30308 10658 30320
rect 10888 30308 10916 30336
rect 14108 30308 14136 30336
rect 10652 30280 10824 30308
rect 10888 30280 11560 30308
rect 10652 30268 10658 30280
rect 10183 30212 10364 30240
rect 10183 30209 10195 30212
rect 10137 30203 10195 30209
rect 9582 30172 9588 30184
rect 8772 30144 9588 30172
rect 8665 30135 8723 30141
rect 9582 30132 9588 30144
rect 9640 30172 9646 30184
rect 9769 30175 9827 30181
rect 9769 30172 9781 30175
rect 9640 30144 9781 30172
rect 9640 30132 9646 30144
rect 9769 30141 9781 30144
rect 9815 30141 9827 30175
rect 9769 30135 9827 30141
rect 10254 30175 10312 30181
rect 10254 30141 10266 30175
rect 10300 30172 10312 30175
rect 10796 30172 10824 30280
rect 10962 30200 10968 30252
rect 11020 30240 11026 30252
rect 11020 30212 11192 30240
rect 11020 30200 11026 30212
rect 11054 30172 11060 30184
rect 10300 30144 10732 30172
rect 10796 30144 11060 30172
rect 10300 30141 10312 30144
rect 10254 30135 10312 30141
rect 3602 30064 3608 30116
rect 3660 30064 3666 30116
rect 6914 30064 6920 30116
rect 6972 30104 6978 30116
rect 10413 30107 10471 30113
rect 10413 30104 10425 30107
rect 6972 30076 10425 30104
rect 6972 30064 6978 30076
rect 10413 30073 10425 30076
rect 10459 30073 10471 30107
rect 10413 30067 10471 30073
rect 10704 30104 10732 30144
rect 11054 30132 11060 30144
rect 11112 30132 11118 30184
rect 11164 30172 11192 30212
rect 11238 30200 11244 30252
rect 11296 30200 11302 30252
rect 11532 30249 11560 30280
rect 13280 30280 14136 30308
rect 11517 30243 11575 30249
rect 11517 30209 11529 30243
rect 11563 30209 11575 30243
rect 11517 30203 11575 30209
rect 11701 30243 11759 30249
rect 11701 30209 11713 30243
rect 11747 30209 11759 30243
rect 11701 30203 11759 30209
rect 11716 30172 11744 30203
rect 11790 30200 11796 30252
rect 11848 30200 11854 30252
rect 13280 30249 13308 30280
rect 14274 30268 14280 30320
rect 14332 30308 14338 30320
rect 18049 30311 18107 30317
rect 14332 30280 14964 30308
rect 14332 30268 14338 30280
rect 13265 30243 13323 30249
rect 13265 30209 13277 30243
rect 13311 30209 13323 30243
rect 13265 30203 13323 30209
rect 14001 30243 14059 30249
rect 14001 30209 14013 30243
rect 14047 30209 14059 30243
rect 14001 30203 14059 30209
rect 14185 30243 14243 30249
rect 14185 30209 14197 30243
rect 14231 30240 14243 30243
rect 14231 30212 14780 30240
rect 14231 30209 14243 30212
rect 14185 30203 14243 30209
rect 11164 30144 11744 30172
rect 13170 30132 13176 30184
rect 13228 30132 13234 30184
rect 14016 30172 14044 30203
rect 14274 30172 14280 30184
rect 13556 30144 14280 30172
rect 13556 30104 13584 30144
rect 14274 30132 14280 30144
rect 14332 30132 14338 30184
rect 10704 30076 13584 30104
rect 13633 30107 13691 30113
rect 5166 29996 5172 30048
rect 5224 30036 5230 30048
rect 5445 30039 5503 30045
rect 5445 30036 5457 30039
rect 5224 30008 5457 30036
rect 5224 29996 5230 30008
rect 5445 30005 5457 30008
rect 5491 30036 5503 30039
rect 7098 30036 7104 30048
rect 5491 30008 7104 30036
rect 5491 30005 5503 30008
rect 5445 29999 5503 30005
rect 7098 29996 7104 30008
rect 7156 30036 7162 30048
rect 7926 30036 7932 30048
rect 7156 30008 7932 30036
rect 7156 29996 7162 30008
rect 7926 29996 7932 30008
rect 7984 29996 7990 30048
rect 8110 29996 8116 30048
rect 8168 29996 8174 30048
rect 8386 29996 8392 30048
rect 8444 30036 8450 30048
rect 8846 30036 8852 30048
rect 8444 30008 8852 30036
rect 8444 29996 8450 30008
rect 8846 29996 8852 30008
rect 8904 30036 8910 30048
rect 9582 30036 9588 30048
rect 8904 30008 9588 30036
rect 8904 29996 8910 30008
rect 9582 29996 9588 30008
rect 9640 29996 9646 30048
rect 10704 30045 10732 30076
rect 13633 30073 13645 30107
rect 13679 30104 13691 30107
rect 13906 30104 13912 30116
rect 13679 30076 13912 30104
rect 13679 30073 13691 30076
rect 13633 30067 13691 30073
rect 13906 30064 13912 30076
rect 13964 30064 13970 30116
rect 13998 30064 14004 30116
rect 14056 30104 14062 30116
rect 14553 30107 14611 30113
rect 14553 30104 14565 30107
rect 14056 30076 14565 30104
rect 14056 30064 14062 30076
rect 14553 30073 14565 30076
rect 14599 30073 14611 30107
rect 14752 30104 14780 30212
rect 14826 30200 14832 30252
rect 14884 30200 14890 30252
rect 14936 30249 14964 30280
rect 18049 30277 18061 30311
rect 18095 30308 18107 30311
rect 18598 30308 18604 30320
rect 18095 30280 18604 30308
rect 18095 30277 18107 30280
rect 18049 30271 18107 30277
rect 18598 30268 18604 30280
rect 18656 30308 18662 30320
rect 18656 30280 18828 30308
rect 18656 30268 18662 30280
rect 14921 30243 14979 30249
rect 14921 30209 14933 30243
rect 14967 30240 14979 30243
rect 15102 30240 15108 30252
rect 14967 30212 15108 30240
rect 14967 30209 14979 30212
rect 14921 30203 14979 30209
rect 15102 30200 15108 30212
rect 15160 30200 15166 30252
rect 17586 30200 17592 30252
rect 17644 30240 17650 30252
rect 17865 30243 17923 30249
rect 17865 30240 17877 30243
rect 17644 30212 17877 30240
rect 17644 30200 17650 30212
rect 17865 30209 17877 30212
rect 17911 30209 17923 30243
rect 17865 30203 17923 30209
rect 18141 30243 18199 30249
rect 18141 30209 18153 30243
rect 18187 30240 18199 30243
rect 18187 30212 18460 30240
rect 18187 30209 18199 30212
rect 18141 30203 18199 30209
rect 17678 30132 17684 30184
rect 17736 30132 17742 30184
rect 18322 30132 18328 30184
rect 18380 30132 18386 30184
rect 18432 30172 18460 30212
rect 18506 30200 18512 30252
rect 18564 30200 18570 30252
rect 18800 30249 18828 30280
rect 18966 30268 18972 30320
rect 19024 30308 19030 30320
rect 19153 30311 19211 30317
rect 19024 30280 19104 30308
rect 19024 30268 19030 30280
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 18874 30200 18880 30252
rect 18932 30200 18938 30252
rect 19076 30249 19104 30280
rect 19153 30277 19165 30311
rect 19199 30308 19211 30311
rect 19358 30308 19386 30348
rect 19610 30336 19616 30348
rect 19668 30336 19674 30388
rect 20714 30336 20720 30388
rect 20772 30376 20778 30388
rect 21818 30376 21824 30388
rect 20772 30348 21824 30376
rect 20772 30336 20778 30348
rect 21818 30336 21824 30348
rect 21876 30376 21882 30388
rect 22189 30379 22247 30385
rect 22189 30376 22201 30379
rect 21876 30348 22201 30376
rect 21876 30336 21882 30348
rect 22189 30345 22201 30348
rect 22235 30345 22247 30379
rect 22189 30339 22247 30345
rect 24854 30336 24860 30388
rect 24912 30376 24918 30388
rect 24912 30348 25452 30376
rect 24912 30336 24918 30348
rect 20732 30308 20760 30336
rect 19199 30280 19386 30308
rect 19444 30280 20760 30308
rect 19199 30277 19211 30280
rect 19153 30271 19211 30277
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30240 19119 30243
rect 19107 30212 19196 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 18966 30172 18972 30184
rect 18432 30144 18972 30172
rect 14752 30076 14964 30104
rect 14553 30067 14611 30073
rect 10689 30039 10747 30045
rect 10689 30005 10701 30039
rect 10735 30005 10747 30039
rect 10689 29999 10747 30005
rect 10778 29996 10784 30048
rect 10836 30036 10842 30048
rect 11057 30039 11115 30045
rect 11057 30036 11069 30039
rect 10836 30008 11069 30036
rect 10836 29996 10842 30008
rect 11057 30005 11069 30008
rect 11103 30005 11115 30039
rect 11057 29999 11115 30005
rect 11606 29996 11612 30048
rect 11664 30036 11670 30048
rect 11885 30039 11943 30045
rect 11885 30036 11897 30039
rect 11664 30008 11897 30036
rect 11664 29996 11670 30008
rect 11885 30005 11897 30008
rect 11931 30036 11943 30039
rect 13262 30036 13268 30048
rect 11931 30008 13268 30036
rect 11931 30005 11943 30008
rect 11885 29999 11943 30005
rect 13262 29996 13268 30008
rect 13320 29996 13326 30048
rect 14936 30045 14964 30076
rect 16850 30064 16856 30116
rect 16908 30104 16914 30116
rect 18233 30107 18291 30113
rect 18233 30104 18245 30107
rect 16908 30076 18245 30104
rect 16908 30064 16914 30076
rect 18233 30073 18245 30076
rect 18279 30073 18291 30107
rect 18233 30067 18291 30073
rect 14921 30039 14979 30045
rect 14921 30005 14933 30039
rect 14967 30036 14979 30039
rect 18432 30036 18460 30144
rect 18966 30132 18972 30144
rect 19024 30132 19030 30184
rect 19168 30104 19196 30212
rect 19242 30200 19248 30252
rect 19300 30200 19306 30252
rect 19334 30132 19340 30184
rect 19392 30132 19398 30184
rect 19444 30181 19472 30280
rect 21634 30268 21640 30320
rect 21692 30308 21698 30320
rect 23198 30308 23204 30320
rect 21692 30280 23204 30308
rect 21692 30268 21698 30280
rect 19705 30243 19763 30249
rect 19705 30209 19717 30243
rect 19751 30240 19763 30243
rect 20622 30240 20628 30252
rect 19751 30212 20628 30240
rect 19751 30209 19763 30212
rect 19705 30203 19763 30209
rect 20622 30200 20628 30212
rect 20680 30200 20686 30252
rect 20714 30200 20720 30252
rect 20772 30240 20778 30252
rect 22002 30240 22008 30252
rect 20772 30212 22008 30240
rect 20772 30200 20778 30212
rect 22002 30200 22008 30212
rect 22060 30200 22066 30252
rect 22462 30240 22468 30252
rect 22301 30212 22468 30240
rect 19429 30175 19487 30181
rect 19429 30141 19441 30175
rect 19475 30141 19487 30175
rect 19429 30135 19487 30141
rect 22301 30116 22329 30212
rect 22462 30200 22468 30212
rect 22520 30241 22526 30252
rect 22664 30249 22692 30280
rect 23198 30268 23204 30280
rect 23256 30268 23262 30320
rect 23842 30308 23848 30320
rect 23492 30280 23848 30308
rect 22557 30243 22615 30249
rect 22557 30241 22569 30243
rect 22520 30213 22569 30241
rect 22520 30200 22526 30213
rect 22557 30209 22569 30213
rect 22603 30209 22615 30243
rect 22557 30203 22615 30209
rect 22649 30243 22707 30249
rect 22649 30209 22661 30243
rect 22695 30209 22707 30243
rect 22649 30203 22707 30209
rect 22738 30200 22744 30252
rect 22796 30200 22802 30252
rect 22830 30200 22836 30252
rect 22888 30249 22894 30252
rect 23492 30249 23520 30280
rect 23842 30268 23848 30280
rect 23900 30268 23906 30320
rect 24302 30268 24308 30320
rect 24360 30308 24366 30320
rect 24486 30308 24492 30320
rect 24360 30280 24492 30308
rect 24360 30268 24366 30280
rect 24486 30268 24492 30280
rect 24544 30308 24550 30320
rect 25424 30308 25452 30348
rect 26878 30336 26884 30388
rect 26936 30376 26942 30388
rect 27062 30376 27068 30388
rect 26936 30348 27068 30376
rect 26936 30336 26942 30348
rect 27062 30336 27068 30348
rect 27120 30376 27126 30388
rect 27430 30376 27436 30388
rect 27120 30348 27436 30376
rect 27120 30336 27126 30348
rect 27430 30336 27436 30348
rect 27488 30336 27494 30388
rect 27706 30376 27712 30388
rect 27632 30348 27712 30376
rect 27448 30308 27476 30336
rect 27632 30317 27660 30348
rect 27706 30336 27712 30348
rect 27764 30336 27770 30388
rect 27982 30336 27988 30388
rect 28040 30376 28046 30388
rect 28040 30348 29960 30376
rect 28040 30336 28046 30348
rect 24544 30280 24610 30308
rect 25424 30280 27200 30308
rect 24544 30268 24550 30280
rect 22888 30243 22917 30249
rect 22905 30240 22917 30243
rect 23293 30243 23351 30249
rect 23293 30240 23305 30243
rect 22905 30212 23305 30240
rect 22905 30209 22917 30212
rect 22888 30203 22917 30209
rect 23293 30209 23305 30212
rect 23339 30209 23351 30243
rect 23293 30203 23351 30209
rect 23477 30243 23535 30249
rect 23477 30209 23489 30243
rect 23523 30209 23535 30243
rect 23477 30203 23535 30209
rect 23569 30243 23627 30249
rect 23569 30209 23581 30243
rect 23615 30209 23627 30243
rect 23569 30203 23627 30209
rect 22888 30200 22894 30203
rect 22370 30132 22376 30184
rect 22428 30132 22434 30184
rect 23017 30175 23075 30181
rect 23017 30172 23029 30175
rect 22664 30144 23029 30172
rect 22278 30104 22284 30116
rect 19168 30076 22284 30104
rect 22278 30064 22284 30076
rect 22336 30064 22342 30116
rect 22388 30104 22416 30132
rect 22664 30116 22692 30144
rect 23017 30141 23029 30144
rect 23063 30141 23075 30175
rect 23584 30172 23612 30203
rect 23750 30200 23756 30252
rect 23808 30200 23814 30252
rect 26142 30200 26148 30252
rect 26200 30240 26206 30252
rect 26329 30243 26387 30249
rect 26329 30240 26341 30243
rect 26200 30212 26341 30240
rect 26200 30200 26206 30212
rect 26329 30209 26341 30212
rect 26375 30209 26387 30243
rect 26329 30203 26387 30209
rect 26421 30243 26479 30249
rect 26421 30209 26433 30243
rect 26467 30209 26479 30243
rect 26421 30203 26479 30209
rect 26513 30243 26571 30249
rect 26513 30209 26525 30243
rect 26559 30240 26571 30243
rect 26602 30240 26608 30252
rect 26559 30212 26608 30240
rect 26559 30209 26571 30212
rect 26513 30203 26571 30209
rect 23017 30135 23075 30141
rect 23492 30144 23612 30172
rect 22388 30076 22600 30104
rect 14967 30008 18460 30036
rect 14967 30005 14979 30008
rect 14921 29999 14979 30005
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 19521 30039 19579 30045
rect 19521 30036 19533 30039
rect 19392 30008 19533 30036
rect 19392 29996 19398 30008
rect 19521 30005 19533 30008
rect 19567 30005 19579 30039
rect 19521 29999 19579 30005
rect 19610 29996 19616 30048
rect 19668 30036 19674 30048
rect 20070 30036 20076 30048
rect 19668 30008 20076 30036
rect 19668 29996 19674 30008
rect 20070 29996 20076 30008
rect 20128 30036 20134 30048
rect 22094 30036 22100 30048
rect 20128 30008 22100 30036
rect 20128 29996 20134 30008
rect 22094 29996 22100 30008
rect 22152 29996 22158 30048
rect 22373 30039 22431 30045
rect 22373 30005 22385 30039
rect 22419 30036 22431 30039
rect 22462 30036 22468 30048
rect 22419 30008 22468 30036
rect 22419 30005 22431 30008
rect 22373 29999 22431 30005
rect 22462 29996 22468 30008
rect 22520 29996 22526 30048
rect 22572 30036 22600 30076
rect 22646 30064 22652 30116
rect 22704 30064 22710 30116
rect 23492 30104 23520 30144
rect 23934 30132 23940 30184
rect 23992 30132 23998 30184
rect 24029 30175 24087 30181
rect 24029 30141 24041 30175
rect 24075 30172 24087 30175
rect 25777 30175 25835 30181
rect 24075 30144 24164 30172
rect 24075 30141 24087 30144
rect 24029 30135 24087 30141
rect 22848 30076 23520 30104
rect 22848 30036 22876 30076
rect 22572 30008 22876 30036
rect 22922 29996 22928 30048
rect 22980 30036 22986 30048
rect 23109 30039 23167 30045
rect 23109 30036 23121 30039
rect 22980 30008 23121 30036
rect 22980 29996 22986 30008
rect 23109 30005 23121 30008
rect 23155 30005 23167 30039
rect 23109 29999 23167 30005
rect 23198 29996 23204 30048
rect 23256 30036 23262 30048
rect 24136 30036 24164 30144
rect 25777 30141 25789 30175
rect 25823 30172 25835 30175
rect 26053 30175 26111 30181
rect 25823 30144 26004 30172
rect 25823 30141 25835 30144
rect 25777 30135 25835 30141
rect 25976 30104 26004 30144
rect 26053 30141 26065 30175
rect 26099 30172 26111 30175
rect 26234 30172 26240 30184
rect 26099 30144 26240 30172
rect 26099 30141 26111 30144
rect 26053 30135 26111 30141
rect 26234 30132 26240 30144
rect 26292 30132 26298 30184
rect 26145 30107 26203 30113
rect 26145 30104 26157 30107
rect 25976 30076 26157 30104
rect 26145 30073 26157 30076
rect 26191 30073 26203 30107
rect 26145 30067 26203 30073
rect 26436 30036 26464 30203
rect 26602 30200 26608 30212
rect 26660 30200 26666 30252
rect 27172 30249 27200 30280
rect 27264 30280 27476 30308
rect 27617 30311 27675 30317
rect 27264 30249 27292 30280
rect 27617 30277 27629 30311
rect 27663 30277 27675 30311
rect 28074 30308 28080 30320
rect 27617 30271 27675 30277
rect 27908 30280 28080 30308
rect 26697 30243 26755 30249
rect 26697 30209 26709 30243
rect 26743 30209 26755 30243
rect 26697 30203 26755 30209
rect 27157 30243 27215 30249
rect 27157 30209 27169 30243
rect 27203 30209 27215 30243
rect 27157 30203 27215 30209
rect 27249 30243 27307 30249
rect 27249 30209 27261 30243
rect 27295 30209 27307 30243
rect 27249 30203 27307 30209
rect 26712 30172 26740 30203
rect 27338 30200 27344 30252
rect 27396 30240 27402 30252
rect 27908 30249 27936 30280
rect 28074 30268 28080 30280
rect 28132 30308 28138 30320
rect 28169 30311 28227 30317
rect 28169 30308 28181 30311
rect 28132 30280 28181 30308
rect 28132 30268 28138 30280
rect 28169 30277 28181 30280
rect 28215 30308 28227 30311
rect 28258 30308 28264 30320
rect 28215 30280 28264 30308
rect 28215 30277 28227 30280
rect 28169 30271 28227 30277
rect 28258 30268 28264 30280
rect 28316 30268 28322 30320
rect 28813 30311 28871 30317
rect 28813 30308 28825 30311
rect 28552 30280 28825 30308
rect 27709 30243 27767 30249
rect 27709 30240 27721 30243
rect 27396 30212 27721 30240
rect 27396 30200 27402 30212
rect 27709 30209 27721 30212
rect 27755 30209 27767 30243
rect 27709 30203 27767 30209
rect 27893 30243 27951 30249
rect 27893 30209 27905 30243
rect 27939 30209 27951 30243
rect 27893 30203 27951 30209
rect 28442 30200 28448 30252
rect 28500 30240 28506 30252
rect 28552 30240 28580 30280
rect 28813 30277 28825 30280
rect 28859 30277 28871 30311
rect 28813 30271 28871 30277
rect 28500 30212 28580 30240
rect 28500 30200 28506 30212
rect 28629 30209 28687 30215
rect 27525 30175 27583 30181
rect 26712 30144 27476 30172
rect 27448 30048 27476 30144
rect 27525 30141 27537 30175
rect 27571 30172 27583 30175
rect 28166 30172 28172 30184
rect 27571 30144 28172 30172
rect 27571 30141 27583 30144
rect 27525 30135 27583 30141
rect 27908 30116 27936 30144
rect 28166 30132 28172 30144
rect 28224 30132 28230 30184
rect 28258 30132 28264 30184
rect 28316 30172 28322 30184
rect 28353 30175 28411 30181
rect 28353 30172 28365 30175
rect 28316 30144 28365 30172
rect 28316 30132 28322 30144
rect 28353 30141 28365 30144
rect 28399 30141 28411 30175
rect 28537 30175 28595 30181
rect 28537 30172 28549 30175
rect 28353 30135 28411 30141
rect 28460 30144 28549 30172
rect 27890 30064 27896 30116
rect 27948 30064 27954 30116
rect 28074 30064 28080 30116
rect 28132 30104 28138 30116
rect 28460 30104 28488 30144
rect 28537 30141 28549 30144
rect 28583 30141 28595 30175
rect 28629 30175 28641 30209
rect 28675 30175 28687 30209
rect 28718 30200 28724 30252
rect 28776 30200 28782 30252
rect 28902 30200 28908 30252
rect 28960 30200 28966 30252
rect 28994 30200 29000 30252
rect 29052 30200 29058 30252
rect 29362 30240 29368 30252
rect 29104 30212 29368 30240
rect 28629 30169 28687 30175
rect 29104 30172 29132 30212
rect 29362 30200 29368 30212
rect 29420 30200 29426 30252
rect 29546 30200 29552 30252
rect 29604 30240 29610 30252
rect 29825 30243 29883 30249
rect 29825 30240 29837 30243
rect 29604 30212 29837 30240
rect 29604 30200 29610 30212
rect 29825 30209 29837 30212
rect 29871 30209 29883 30243
rect 29932 30240 29960 30348
rect 30006 30268 30012 30320
rect 30064 30308 30070 30320
rect 30064 30280 34284 30308
rect 30064 30268 30070 30280
rect 30190 30240 30196 30252
rect 29932 30212 30196 30240
rect 29825 30203 29883 30209
rect 30190 30200 30196 30212
rect 30248 30240 30254 30252
rect 30285 30243 30343 30249
rect 30285 30240 30297 30243
rect 30248 30212 30297 30240
rect 30248 30200 30254 30212
rect 30285 30209 30297 30212
rect 30331 30209 30343 30243
rect 30285 30203 30343 30209
rect 30392 30212 30604 30240
rect 28537 30135 28595 30141
rect 28132 30076 28488 30104
rect 28644 30104 28672 30169
rect 28966 30164 29132 30172
rect 28828 30144 29132 30164
rect 28828 30136 28994 30144
rect 28828 30104 28856 30136
rect 29178 30132 29184 30184
rect 29236 30172 29242 30184
rect 29457 30175 29515 30181
rect 29457 30172 29469 30175
rect 29236 30144 29469 30172
rect 29236 30132 29242 30144
rect 29457 30141 29469 30144
rect 29503 30172 29515 30175
rect 30392 30172 30420 30212
rect 29503 30144 30420 30172
rect 30576 30172 30604 30212
rect 30650 30200 30656 30252
rect 30708 30200 30714 30252
rect 30837 30243 30895 30249
rect 30837 30209 30849 30243
rect 30883 30240 30895 30243
rect 31110 30240 31116 30252
rect 30883 30212 31116 30240
rect 30883 30209 30895 30212
rect 30837 30203 30895 30209
rect 31110 30200 31116 30212
rect 31168 30240 31174 30252
rect 31478 30240 31484 30252
rect 31168 30212 31484 30240
rect 31168 30200 31174 30212
rect 31478 30200 31484 30212
rect 31536 30200 31542 30252
rect 33042 30200 33048 30252
rect 33100 30200 33106 30252
rect 33152 30249 33180 30280
rect 33138 30243 33196 30249
rect 33138 30209 33150 30243
rect 33184 30209 33196 30243
rect 33138 30203 33196 30209
rect 33318 30200 33324 30252
rect 33376 30200 33382 30252
rect 33410 30200 33416 30252
rect 33468 30200 33474 30252
rect 34256 30249 34284 30280
rect 33510 30243 33568 30249
rect 33510 30209 33522 30243
rect 33556 30209 33568 30243
rect 33510 30203 33568 30209
rect 34241 30243 34299 30249
rect 34241 30209 34253 30243
rect 34287 30209 34299 30243
rect 34241 30203 34299 30209
rect 32398 30172 32404 30184
rect 30576 30144 32404 30172
rect 29503 30141 29515 30144
rect 29457 30135 29515 30141
rect 32398 30132 32404 30144
rect 32456 30132 32462 30184
rect 33520 30172 33548 30203
rect 34422 30200 34428 30252
rect 34480 30200 34486 30252
rect 34330 30172 34336 30184
rect 33152 30144 34336 30172
rect 30466 30104 30472 30116
rect 28644 30076 28856 30104
rect 28132 30064 28138 30076
rect 23256 30008 26464 30036
rect 23256 29996 23262 30008
rect 26878 29996 26884 30048
rect 26936 30036 26942 30048
rect 26973 30039 27031 30045
rect 26973 30036 26985 30039
rect 26936 30008 26985 30036
rect 26936 29996 26942 30008
rect 26973 30005 26985 30008
rect 27019 30005 27031 30039
rect 26973 29999 27031 30005
rect 27430 29996 27436 30048
rect 27488 30036 27494 30048
rect 27709 30039 27767 30045
rect 27709 30036 27721 30039
rect 27488 30008 27721 30036
rect 27488 29996 27494 30008
rect 27709 30005 27721 30008
rect 27755 30005 27767 30039
rect 27709 29999 27767 30005
rect 28534 29996 28540 30048
rect 28592 30036 28598 30048
rect 28828 30036 28856 30076
rect 28966 30076 30472 30104
rect 28966 30048 28994 30076
rect 30466 30064 30472 30076
rect 30524 30064 30530 30116
rect 28592 30008 28856 30036
rect 28592 29996 28598 30008
rect 28902 29996 28908 30048
rect 28960 30008 28994 30048
rect 28960 29996 28966 30008
rect 29638 29996 29644 30048
rect 29696 30036 29702 30048
rect 29917 30039 29975 30045
rect 29917 30036 29929 30039
rect 29696 30008 29929 30036
rect 29696 29996 29702 30008
rect 29917 30005 29929 30008
rect 29963 30005 29975 30039
rect 29917 29999 29975 30005
rect 30558 29996 30564 30048
rect 30616 30036 30622 30048
rect 31570 30036 31576 30048
rect 30616 30008 31576 30036
rect 30616 29996 30622 30008
rect 31570 29996 31576 30008
rect 31628 30036 31634 30048
rect 33152 30036 33180 30144
rect 34330 30132 34336 30144
rect 34388 30132 34394 30184
rect 33226 30064 33232 30116
rect 33284 30104 33290 30116
rect 34057 30107 34115 30113
rect 34057 30104 34069 30107
rect 33284 30076 34069 30104
rect 33284 30064 33290 30076
rect 34057 30073 34069 30076
rect 34103 30073 34115 30107
rect 34057 30067 34115 30073
rect 31628 30008 33180 30036
rect 31628 29996 31634 30008
rect 33594 29996 33600 30048
rect 33652 30036 33658 30048
rect 33689 30039 33747 30045
rect 33689 30036 33701 30039
rect 33652 30008 33701 30036
rect 33652 29996 33658 30008
rect 33689 30005 33701 30008
rect 33735 30005 33747 30039
rect 33689 29999 33747 30005
rect 1104 29946 36432 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 36432 29946
rect 1104 29872 36432 29894
rect 1302 29792 1308 29844
rect 1360 29832 1366 29844
rect 1360 29804 3556 29832
rect 1360 29792 1366 29804
rect 3528 29764 3556 29804
rect 3602 29792 3608 29844
rect 3660 29832 3666 29844
rect 3789 29835 3847 29841
rect 3789 29832 3801 29835
rect 3660 29804 3801 29832
rect 3660 29792 3666 29804
rect 3789 29801 3801 29804
rect 3835 29801 3847 29835
rect 3789 29795 3847 29801
rect 3970 29792 3976 29844
rect 4028 29832 4034 29844
rect 4801 29835 4859 29841
rect 4801 29832 4813 29835
rect 4028 29804 4813 29832
rect 4028 29792 4034 29804
rect 4801 29801 4813 29804
rect 4847 29801 4859 29835
rect 4801 29795 4859 29801
rect 8938 29792 8944 29844
rect 8996 29792 9002 29844
rect 9214 29792 9220 29844
rect 9272 29832 9278 29844
rect 10410 29832 10416 29844
rect 9272 29804 10416 29832
rect 9272 29792 9278 29804
rect 10410 29792 10416 29804
rect 10468 29792 10474 29844
rect 10502 29792 10508 29844
rect 10560 29832 10566 29844
rect 10689 29835 10747 29841
rect 10689 29832 10701 29835
rect 10560 29804 10701 29832
rect 10560 29792 10566 29804
rect 10689 29801 10701 29804
rect 10735 29832 10747 29835
rect 10962 29832 10968 29844
rect 10735 29804 10968 29832
rect 10735 29801 10747 29804
rect 10689 29795 10747 29801
rect 10962 29792 10968 29804
rect 11020 29792 11026 29844
rect 15470 29792 15476 29844
rect 15528 29832 15534 29844
rect 15528 29804 16160 29832
rect 15528 29792 15534 29804
rect 3528 29736 4292 29764
rect 1489 29699 1547 29705
rect 1489 29665 1501 29699
rect 1535 29696 1547 29699
rect 3142 29696 3148 29708
rect 1535 29668 3148 29696
rect 1535 29665 1547 29668
rect 1489 29659 1547 29665
rect 3142 29656 3148 29668
rect 3200 29656 3206 29708
rect 3234 29656 3240 29708
rect 3292 29656 3298 29708
rect 3513 29699 3571 29705
rect 3513 29665 3525 29699
rect 3559 29696 3571 29699
rect 3694 29696 3700 29708
rect 3559 29668 3700 29696
rect 3559 29665 3571 29668
rect 3513 29659 3571 29665
rect 3694 29656 3700 29668
rect 3752 29656 3758 29708
rect 4264 29705 4292 29736
rect 4249 29699 4307 29705
rect 4249 29665 4261 29699
rect 4295 29665 4307 29699
rect 4249 29659 4307 29665
rect 4341 29699 4399 29705
rect 4341 29665 4353 29699
rect 4387 29665 4399 29699
rect 4341 29659 4399 29665
rect 5445 29699 5503 29705
rect 5445 29665 5457 29699
rect 5491 29696 5503 29699
rect 6270 29696 6276 29708
rect 5491 29668 6276 29696
rect 5491 29665 5503 29668
rect 5445 29659 5503 29665
rect 4062 29588 4068 29640
rect 4120 29628 4126 29640
rect 4356 29628 4384 29659
rect 6270 29656 6276 29668
rect 6328 29656 6334 29708
rect 7098 29656 7104 29708
rect 7156 29696 7162 29708
rect 8386 29696 8392 29708
rect 7156 29668 8392 29696
rect 7156 29656 7162 29668
rect 4120 29600 4384 29628
rect 5261 29631 5319 29637
rect 4120 29588 4126 29600
rect 5261 29597 5273 29631
rect 5307 29628 5319 29631
rect 5534 29628 5540 29640
rect 5307 29600 5540 29628
rect 5307 29597 5319 29600
rect 5261 29591 5319 29597
rect 5534 29588 5540 29600
rect 5592 29588 5598 29640
rect 5626 29588 5632 29640
rect 5684 29628 5690 29640
rect 5810 29628 5816 29640
rect 5684 29600 5816 29628
rect 5684 29588 5690 29600
rect 5810 29588 5816 29600
rect 5868 29628 5874 29640
rect 6546 29628 6552 29640
rect 5868 29600 6552 29628
rect 5868 29588 5874 29600
rect 6546 29588 6552 29600
rect 6604 29588 6610 29640
rect 7377 29631 7435 29637
rect 7377 29597 7389 29631
rect 7423 29628 7435 29631
rect 7558 29628 7564 29640
rect 7423 29600 7564 29628
rect 7423 29597 7435 29600
rect 7377 29591 7435 29597
rect 7558 29588 7564 29600
rect 7616 29588 7622 29640
rect 7760 29637 7788 29668
rect 8386 29656 8392 29668
rect 8444 29656 8450 29708
rect 7745 29631 7803 29637
rect 7745 29597 7757 29631
rect 7791 29597 7803 29631
rect 7745 29591 7803 29597
rect 8110 29588 8116 29640
rect 8168 29588 8174 29640
rect 8297 29631 8355 29637
rect 8297 29597 8309 29631
rect 8343 29628 8355 29631
rect 8662 29628 8668 29640
rect 8343 29600 8668 29628
rect 8343 29597 8355 29600
rect 8297 29591 8355 29597
rect 8662 29588 8668 29600
rect 8720 29588 8726 29640
rect 4157 29563 4215 29569
rect 2806 29532 3096 29560
rect 3068 29504 3096 29532
rect 4157 29529 4169 29563
rect 4203 29560 4215 29563
rect 5350 29560 5356 29572
rect 4203 29532 5356 29560
rect 4203 29529 4215 29532
rect 4157 29523 4215 29529
rect 5350 29520 5356 29532
rect 5408 29520 5414 29572
rect 3050 29452 3056 29504
rect 3108 29452 3114 29504
rect 4706 29452 4712 29504
rect 4764 29492 4770 29504
rect 5166 29492 5172 29504
rect 4764 29464 5172 29492
rect 4764 29452 4770 29464
rect 5166 29452 5172 29464
rect 5224 29452 5230 29504
rect 5718 29452 5724 29504
rect 5776 29452 5782 29504
rect 8956 29501 8984 29792
rect 9122 29724 9128 29776
rect 9180 29764 9186 29776
rect 11885 29767 11943 29773
rect 11885 29764 11897 29767
rect 9180 29736 11897 29764
rect 9180 29724 9186 29736
rect 11885 29733 11897 29736
rect 11931 29733 11943 29767
rect 13078 29764 13084 29776
rect 11885 29727 11943 29733
rect 12176 29736 13084 29764
rect 9585 29699 9643 29705
rect 9585 29665 9597 29699
rect 9631 29696 9643 29699
rect 9766 29696 9772 29708
rect 9631 29668 9772 29696
rect 9631 29665 9643 29668
rect 9585 29659 9643 29665
rect 9766 29656 9772 29668
rect 9824 29656 9830 29708
rect 11606 29696 11612 29708
rect 10152 29668 11612 29696
rect 9306 29588 9312 29640
rect 9364 29628 9370 29640
rect 10152 29628 10180 29668
rect 11606 29656 11612 29668
rect 11664 29656 11670 29708
rect 12176 29705 12204 29736
rect 13078 29724 13084 29736
rect 13136 29724 13142 29776
rect 13354 29724 13360 29776
rect 13412 29724 13418 29776
rect 16022 29764 16028 29776
rect 13740 29736 16028 29764
rect 12161 29699 12219 29705
rect 12161 29665 12173 29699
rect 12207 29665 12219 29699
rect 13372 29696 13400 29724
rect 13449 29699 13507 29705
rect 13449 29696 13461 29699
rect 12161 29659 12219 29665
rect 12820 29668 13308 29696
rect 13372 29668 13461 29696
rect 9364 29600 10180 29628
rect 10229 29631 10287 29637
rect 9364 29588 9370 29600
rect 10229 29597 10241 29631
rect 10275 29628 10287 29631
rect 10410 29628 10416 29640
rect 10275 29600 10416 29628
rect 10275 29597 10287 29600
rect 10229 29591 10287 29597
rect 10410 29588 10416 29600
rect 10468 29588 10474 29640
rect 10505 29631 10563 29637
rect 10505 29597 10517 29631
rect 10551 29628 10563 29631
rect 10594 29628 10600 29640
rect 10551 29600 10600 29628
rect 10551 29597 10563 29600
rect 10505 29591 10563 29597
rect 10594 29588 10600 29600
rect 10652 29588 10658 29640
rect 10689 29631 10747 29637
rect 10689 29597 10701 29631
rect 10735 29628 10747 29631
rect 10778 29628 10784 29640
rect 10735 29600 10784 29628
rect 10735 29597 10747 29600
rect 10689 29591 10747 29597
rect 10778 29588 10784 29600
rect 10836 29588 10842 29640
rect 11790 29588 11796 29640
rect 11848 29588 11854 29640
rect 12250 29588 12256 29640
rect 12308 29588 12314 29640
rect 12618 29588 12624 29640
rect 12676 29588 12682 29640
rect 12820 29637 12848 29668
rect 12805 29631 12863 29637
rect 12805 29597 12817 29631
rect 12851 29597 12863 29631
rect 12805 29591 12863 29597
rect 12897 29631 12955 29637
rect 12897 29597 12909 29631
rect 12943 29628 12955 29631
rect 12943 29600 13124 29628
rect 12943 29597 12955 29600
rect 12897 29591 12955 29597
rect 12989 29563 13047 29569
rect 12989 29560 13001 29563
rect 9324 29532 13001 29560
rect 8941 29495 8999 29501
rect 8941 29461 8953 29495
rect 8987 29461 8999 29495
rect 8941 29455 8999 29461
rect 9214 29452 9220 29504
rect 9272 29492 9278 29504
rect 9324 29501 9352 29532
rect 12989 29529 13001 29532
rect 13035 29529 13047 29563
rect 13096 29560 13124 29600
rect 13096 29532 13216 29560
rect 12989 29523 13047 29529
rect 13188 29504 13216 29532
rect 13280 29504 13308 29668
rect 13449 29665 13461 29668
rect 13495 29665 13507 29699
rect 13449 29659 13507 29665
rect 13357 29631 13415 29637
rect 13357 29597 13369 29631
rect 13403 29628 13415 29631
rect 13630 29628 13636 29640
rect 13403 29600 13636 29628
rect 13403 29597 13415 29600
rect 13357 29591 13415 29597
rect 13630 29588 13636 29600
rect 13688 29588 13694 29640
rect 13740 29637 13768 29736
rect 16022 29724 16028 29736
rect 16080 29724 16086 29776
rect 16132 29764 16160 29804
rect 17310 29792 17316 29844
rect 17368 29832 17374 29844
rect 18417 29835 18475 29841
rect 18417 29832 18429 29835
rect 17368 29804 18429 29832
rect 17368 29792 17374 29804
rect 18417 29801 18429 29804
rect 18463 29801 18475 29835
rect 18417 29795 18475 29801
rect 18598 29792 18604 29844
rect 18656 29792 18662 29844
rect 18966 29792 18972 29844
rect 19024 29832 19030 29844
rect 19245 29835 19303 29841
rect 19245 29832 19257 29835
rect 19024 29804 19257 29832
rect 19024 29792 19030 29804
rect 19245 29801 19257 29804
rect 19291 29801 19303 29835
rect 23934 29832 23940 29844
rect 19245 29795 19303 29801
rect 19634 29804 23940 29832
rect 16132 29736 17540 29764
rect 14090 29656 14096 29708
rect 14148 29656 14154 29708
rect 14292 29668 14509 29696
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29597 13783 29631
rect 13725 29591 13783 29597
rect 13740 29560 13768 29591
rect 13814 29588 13820 29640
rect 13872 29628 13878 29640
rect 14292 29628 14320 29668
rect 13872 29600 14320 29628
rect 13872 29588 13878 29600
rect 14366 29588 14372 29640
rect 14424 29588 14430 29640
rect 14481 29637 14509 29668
rect 15286 29656 15292 29708
rect 15344 29656 15350 29708
rect 15841 29699 15899 29705
rect 15841 29665 15853 29699
rect 15887 29696 15899 29699
rect 16574 29696 16580 29708
rect 15887 29668 16580 29696
rect 15887 29665 15899 29668
rect 15841 29659 15899 29665
rect 16574 29656 16580 29668
rect 16632 29656 16638 29708
rect 17402 29696 17408 29708
rect 16868 29668 17408 29696
rect 14466 29631 14524 29637
rect 14466 29597 14478 29631
rect 14512 29597 14524 29631
rect 14466 29591 14524 29597
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29628 15715 29631
rect 15746 29628 15752 29640
rect 15703 29600 15752 29628
rect 15703 29597 15715 29600
rect 15657 29591 15715 29597
rect 15746 29588 15752 29600
rect 15804 29588 15810 29640
rect 16117 29631 16175 29637
rect 16117 29597 16129 29631
rect 16163 29628 16175 29631
rect 16868 29628 16896 29668
rect 17402 29656 17408 29668
rect 17460 29656 17466 29708
rect 17512 29696 17540 29736
rect 18322 29724 18328 29776
rect 18380 29764 18386 29776
rect 18782 29764 18788 29776
rect 18380 29736 18788 29764
rect 18380 29724 18386 29736
rect 18782 29724 18788 29736
rect 18840 29764 18846 29776
rect 19634 29764 19662 29804
rect 23934 29792 23940 29804
rect 23992 29832 23998 29844
rect 23992 29804 26280 29832
rect 23992 29792 23998 29804
rect 18840 29736 19662 29764
rect 18840 29724 18846 29736
rect 19702 29724 19708 29776
rect 19760 29724 19766 29776
rect 20162 29724 20168 29776
rect 20220 29764 20226 29776
rect 21266 29764 21272 29776
rect 20220 29736 21272 29764
rect 20220 29724 20226 29736
rect 21266 29724 21272 29736
rect 21324 29764 21330 29776
rect 21542 29764 21548 29776
rect 21324 29736 21548 29764
rect 21324 29724 21330 29736
rect 21542 29724 21548 29736
rect 21600 29724 21606 29776
rect 22094 29724 22100 29776
rect 22152 29724 22158 29776
rect 22186 29724 22192 29776
rect 22244 29724 22250 29776
rect 22278 29724 22284 29776
rect 22336 29764 22342 29776
rect 22336 29736 23796 29764
rect 22336 29724 22342 29736
rect 19521 29699 19579 29705
rect 19521 29696 19533 29699
rect 17512 29668 19533 29696
rect 19521 29665 19533 29668
rect 19567 29665 19579 29699
rect 19521 29659 19579 29665
rect 19613 29699 19671 29705
rect 19613 29665 19625 29699
rect 19659 29696 19671 29699
rect 19720 29696 19748 29724
rect 19659 29668 21588 29696
rect 19659 29665 19671 29668
rect 19613 29659 19671 29665
rect 16163 29600 16896 29628
rect 16945 29631 17003 29637
rect 16163 29597 16175 29600
rect 16117 29591 16175 29597
rect 16945 29597 16957 29631
rect 16991 29597 17003 29631
rect 16945 29591 17003 29597
rect 13372 29532 13768 29560
rect 13372 29504 13400 29532
rect 13998 29520 14004 29572
rect 14056 29560 14062 29572
rect 14093 29563 14151 29569
rect 14093 29560 14105 29563
rect 14056 29532 14105 29560
rect 14056 29520 14062 29532
rect 14093 29529 14105 29532
rect 14139 29529 14151 29563
rect 14093 29523 14151 29529
rect 14277 29563 14335 29569
rect 14277 29529 14289 29563
rect 14323 29529 14335 29563
rect 14277 29523 14335 29529
rect 9309 29495 9367 29501
rect 9309 29492 9321 29495
rect 9272 29464 9321 29492
rect 9272 29452 9278 29464
rect 9309 29461 9321 29464
rect 9355 29461 9367 29495
rect 9309 29455 9367 29461
rect 9401 29495 9459 29501
rect 9401 29461 9413 29495
rect 9447 29492 9459 29495
rect 9490 29492 9496 29504
rect 9447 29464 9496 29492
rect 9447 29461 9459 29464
rect 9401 29455 9459 29461
rect 9490 29452 9496 29464
rect 9548 29452 9554 29504
rect 10226 29452 10232 29504
rect 10284 29492 10290 29504
rect 10321 29495 10379 29501
rect 10321 29492 10333 29495
rect 10284 29464 10333 29492
rect 10284 29452 10290 29464
rect 10321 29461 10333 29464
rect 10367 29461 10379 29495
rect 10321 29455 10379 29461
rect 13170 29452 13176 29504
rect 13228 29452 13234 29504
rect 13262 29452 13268 29504
rect 13320 29452 13326 29504
rect 13354 29452 13360 29504
rect 13412 29452 13418 29504
rect 13630 29452 13636 29504
rect 13688 29492 13694 29504
rect 14292 29492 14320 29523
rect 15562 29520 15568 29572
rect 15620 29560 15626 29572
rect 16206 29560 16212 29572
rect 15620 29532 16212 29560
rect 15620 29520 15626 29532
rect 16206 29520 16212 29532
rect 16264 29520 16270 29572
rect 16301 29563 16359 29569
rect 16301 29529 16313 29563
rect 16347 29529 16359 29563
rect 16301 29523 16359 29529
rect 16439 29563 16497 29569
rect 16439 29529 16451 29563
rect 16485 29560 16497 29563
rect 16960 29560 16988 29591
rect 17034 29588 17040 29640
rect 17092 29628 17098 29640
rect 17129 29631 17187 29637
rect 17129 29628 17141 29631
rect 17092 29600 17141 29628
rect 17092 29588 17098 29600
rect 17129 29597 17141 29600
rect 17175 29628 17187 29631
rect 17678 29628 17684 29640
rect 17175 29600 17684 29628
rect 17175 29597 17187 29600
rect 17129 29591 17187 29597
rect 17678 29588 17684 29600
rect 17736 29588 17742 29640
rect 17954 29588 17960 29640
rect 18012 29628 18018 29640
rect 18141 29631 18199 29637
rect 18141 29628 18153 29631
rect 18012 29600 18153 29628
rect 18012 29588 18018 29600
rect 18141 29597 18153 29600
rect 18187 29597 18199 29631
rect 18141 29591 18199 29597
rect 18506 29588 18512 29640
rect 18564 29588 18570 29640
rect 18877 29631 18935 29637
rect 18877 29597 18889 29631
rect 18923 29628 18935 29631
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 18923 29600 19441 29628
rect 18923 29597 18935 29600
rect 18877 29591 18935 29597
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 19702 29588 19708 29640
rect 19760 29588 19766 29640
rect 17770 29560 17776 29572
rect 16485 29532 16896 29560
rect 16960 29532 17776 29560
rect 16485 29529 16497 29532
rect 16439 29523 16497 29529
rect 13688 29464 14320 29492
rect 15657 29495 15715 29501
rect 13688 29452 13694 29464
rect 15657 29461 15669 29495
rect 15703 29492 15715 29495
rect 15838 29492 15844 29504
rect 15703 29464 15844 29492
rect 15703 29461 15715 29464
rect 15657 29455 15715 29461
rect 15838 29452 15844 29464
rect 15896 29452 15902 29504
rect 15933 29495 15991 29501
rect 15933 29461 15945 29495
rect 15979 29492 15991 29495
rect 16114 29492 16120 29504
rect 15979 29464 16120 29492
rect 15979 29461 15991 29464
rect 15933 29455 15991 29461
rect 16114 29452 16120 29464
rect 16172 29452 16178 29504
rect 16316 29492 16344 29523
rect 16666 29492 16672 29504
rect 16316 29464 16672 29492
rect 16666 29452 16672 29464
rect 16724 29452 16730 29504
rect 16758 29452 16764 29504
rect 16816 29452 16822 29504
rect 16868 29492 16896 29532
rect 17770 29520 17776 29532
rect 17828 29520 17834 29572
rect 17862 29520 17868 29572
rect 17920 29560 17926 29572
rect 17920 29532 18368 29560
rect 17920 29520 17926 29532
rect 17034 29492 17040 29504
rect 16868 29464 17040 29492
rect 17034 29452 17040 29464
rect 17092 29492 17098 29504
rect 17954 29492 17960 29504
rect 17092 29464 17960 29492
rect 17092 29452 17098 29464
rect 17954 29452 17960 29464
rect 18012 29452 18018 29504
rect 18230 29452 18236 29504
rect 18288 29452 18294 29504
rect 18340 29492 18368 29532
rect 18414 29520 18420 29572
rect 18472 29560 18478 29572
rect 19610 29560 19616 29572
rect 18472 29532 19616 29560
rect 18472 29520 18478 29532
rect 19610 29520 19616 29532
rect 19668 29520 19674 29572
rect 19812 29492 19840 29668
rect 20625 29631 20683 29637
rect 20625 29597 20637 29631
rect 20671 29597 20683 29631
rect 20625 29591 20683 29597
rect 20640 29560 20668 29591
rect 20806 29588 20812 29640
rect 20864 29588 20870 29640
rect 20898 29588 20904 29640
rect 20956 29588 20962 29640
rect 20990 29588 20996 29640
rect 21048 29588 21054 29640
rect 21177 29631 21235 29637
rect 21177 29597 21189 29631
rect 21223 29628 21235 29631
rect 21266 29628 21272 29640
rect 21223 29600 21272 29628
rect 21223 29597 21235 29600
rect 21177 29591 21235 29597
rect 21266 29588 21272 29600
rect 21324 29588 21330 29640
rect 21450 29560 21456 29572
rect 20640 29532 21456 29560
rect 21450 29520 21456 29532
rect 21508 29520 21514 29572
rect 21560 29560 21588 29668
rect 22002 29656 22008 29708
rect 22060 29696 22066 29708
rect 22060 29668 22876 29696
rect 22060 29656 22066 29668
rect 22848 29640 22876 29668
rect 21637 29631 21695 29637
rect 21637 29597 21649 29631
rect 21683 29628 21695 29631
rect 21726 29628 21732 29640
rect 21683 29600 21732 29628
rect 21683 29597 21695 29600
rect 21637 29591 21695 29597
rect 21726 29588 21732 29600
rect 21784 29588 21790 29640
rect 22646 29588 22652 29640
rect 22704 29588 22710 29640
rect 22830 29588 22836 29640
rect 22888 29588 22894 29640
rect 23290 29588 23296 29640
rect 23348 29588 23354 29640
rect 23768 29637 23796 29736
rect 24486 29724 24492 29776
rect 24544 29764 24550 29776
rect 25409 29767 25467 29773
rect 25409 29764 25421 29767
rect 24544 29736 25421 29764
rect 24544 29724 24550 29736
rect 25409 29733 25421 29736
rect 25455 29733 25467 29767
rect 25409 29727 25467 29733
rect 25961 29767 26019 29773
rect 25961 29733 25973 29767
rect 26007 29764 26019 29767
rect 26142 29764 26148 29776
rect 26007 29736 26148 29764
rect 26007 29733 26019 29736
rect 25961 29727 26019 29733
rect 26142 29724 26148 29736
rect 26200 29724 26206 29776
rect 26252 29764 26280 29804
rect 26326 29792 26332 29844
rect 26384 29832 26390 29844
rect 26881 29835 26939 29841
rect 26881 29832 26893 29835
rect 26384 29804 26893 29832
rect 26384 29792 26390 29804
rect 26881 29801 26893 29804
rect 26927 29801 26939 29835
rect 26881 29795 26939 29801
rect 27154 29792 27160 29844
rect 27212 29832 27218 29844
rect 28169 29835 28227 29841
rect 28169 29832 28181 29835
rect 27212 29804 28181 29832
rect 27212 29792 27218 29804
rect 28169 29801 28181 29804
rect 28215 29801 28227 29835
rect 28169 29795 28227 29801
rect 28442 29792 28448 29844
rect 28500 29832 28506 29844
rect 28902 29832 28908 29844
rect 28500 29804 28908 29832
rect 28500 29792 28506 29804
rect 28902 29792 28908 29804
rect 28960 29792 28966 29844
rect 29178 29792 29184 29844
rect 29236 29832 29242 29844
rect 29822 29832 29828 29844
rect 29236 29804 29828 29832
rect 29236 29792 29242 29804
rect 29822 29792 29828 29804
rect 29880 29832 29886 29844
rect 32030 29832 32036 29844
rect 29880 29804 32036 29832
rect 29880 29792 29886 29804
rect 32030 29792 32036 29804
rect 32088 29792 32094 29844
rect 27893 29767 27951 29773
rect 26252 29736 27660 29764
rect 26970 29696 26976 29708
rect 25608 29668 26976 29696
rect 25608 29637 25636 29668
rect 26970 29656 26976 29668
rect 27028 29656 27034 29708
rect 27522 29656 27528 29708
rect 27580 29656 27586 29708
rect 27632 29696 27660 29736
rect 27893 29733 27905 29767
rect 27939 29764 27951 29767
rect 28534 29764 28540 29776
rect 27939 29736 28540 29764
rect 27939 29733 27951 29736
rect 27893 29727 27951 29733
rect 28534 29724 28540 29736
rect 28592 29724 28598 29776
rect 28994 29764 29000 29776
rect 28644 29736 29000 29764
rect 28644 29696 28672 29736
rect 28994 29724 29000 29736
rect 29052 29724 29058 29776
rect 29086 29724 29092 29776
rect 29144 29764 29150 29776
rect 29144 29736 32076 29764
rect 29144 29724 29150 29736
rect 27632 29668 28672 29696
rect 28902 29656 28908 29708
rect 28960 29696 28966 29708
rect 32048 29705 32076 29736
rect 31757 29699 31815 29705
rect 31757 29696 31769 29699
rect 28960 29668 31769 29696
rect 28960 29656 28966 29668
rect 31757 29665 31769 29668
rect 31803 29665 31815 29699
rect 31757 29659 31815 29665
rect 32033 29699 32091 29705
rect 32033 29665 32045 29699
rect 32079 29665 32091 29699
rect 32033 29659 32091 29665
rect 23753 29631 23811 29637
rect 23753 29597 23765 29631
rect 23799 29597 23811 29631
rect 23753 29591 23811 29597
rect 25593 29631 25651 29637
rect 25593 29597 25605 29631
rect 25639 29597 25651 29631
rect 25593 29591 25651 29597
rect 25774 29588 25780 29640
rect 25832 29588 25838 29640
rect 26421 29631 26479 29637
rect 26421 29597 26433 29631
rect 26467 29628 26479 29631
rect 26786 29628 26792 29640
rect 26467 29600 26792 29628
rect 26467 29597 26479 29600
rect 26421 29591 26479 29597
rect 26786 29588 26792 29600
rect 26844 29588 26850 29640
rect 26878 29588 26884 29640
rect 26936 29588 26942 29640
rect 27062 29588 27068 29640
rect 27120 29588 27126 29640
rect 27157 29631 27215 29637
rect 27157 29597 27169 29631
rect 27203 29628 27215 29631
rect 27338 29628 27344 29640
rect 27203 29600 27344 29628
rect 27203 29597 27215 29600
rect 27157 29591 27215 29597
rect 27338 29588 27344 29600
rect 27396 29588 27402 29640
rect 27706 29588 27712 29640
rect 27764 29628 27770 29640
rect 28077 29631 28135 29637
rect 28077 29628 28089 29631
rect 27764 29600 28089 29628
rect 27764 29588 27770 29600
rect 28077 29597 28089 29600
rect 28123 29597 28135 29631
rect 28077 29591 28135 29597
rect 28258 29588 28264 29640
rect 28316 29588 28322 29640
rect 28442 29588 28448 29640
rect 28500 29628 28506 29640
rect 30466 29628 30472 29640
rect 28500 29600 30472 29628
rect 28500 29588 28506 29600
rect 30466 29588 30472 29600
rect 30524 29588 30530 29640
rect 31205 29631 31263 29637
rect 31205 29628 31217 29631
rect 30760 29600 31217 29628
rect 30760 29572 30788 29600
rect 31205 29597 31217 29600
rect 31251 29597 31263 29631
rect 31205 29591 31263 29597
rect 31389 29631 31447 29637
rect 31389 29597 31401 29631
rect 31435 29597 31447 29631
rect 31389 29591 31447 29597
rect 31665 29631 31723 29637
rect 31665 29597 31677 29631
rect 31711 29597 31723 29631
rect 31665 29591 31723 29597
rect 32125 29631 32183 29637
rect 32125 29597 32137 29631
rect 32171 29628 32183 29631
rect 32950 29628 32956 29640
rect 32171 29600 32956 29628
rect 32171 29597 32183 29600
rect 32125 29591 32183 29597
rect 21560 29532 23060 29560
rect 23032 29504 23060 29532
rect 23658 29520 23664 29572
rect 23716 29560 23722 29572
rect 24581 29563 24639 29569
rect 24581 29560 24593 29563
rect 23716 29532 24593 29560
rect 23716 29520 23722 29532
rect 24581 29529 24593 29532
rect 24627 29560 24639 29563
rect 25041 29563 25099 29569
rect 25041 29560 25053 29563
rect 24627 29532 25053 29560
rect 24627 29529 24639 29532
rect 24581 29523 24639 29529
rect 25041 29529 25053 29532
rect 25087 29529 25099 29563
rect 25041 29523 25099 29529
rect 25222 29520 25228 29572
rect 25280 29560 25286 29572
rect 25280 29532 26096 29560
rect 25280 29520 25286 29532
rect 18340 29464 19840 29492
rect 20990 29452 20996 29504
rect 21048 29492 21054 29504
rect 21361 29495 21419 29501
rect 21361 29492 21373 29495
rect 21048 29464 21373 29492
rect 21048 29452 21054 29464
rect 21361 29461 21373 29464
rect 21407 29461 21419 29495
rect 21361 29455 21419 29461
rect 21634 29452 21640 29504
rect 21692 29492 21698 29504
rect 21729 29495 21787 29501
rect 21729 29492 21741 29495
rect 21692 29464 21741 29492
rect 21692 29452 21698 29464
rect 21729 29461 21741 29464
rect 21775 29461 21787 29495
rect 21729 29455 21787 29461
rect 23014 29452 23020 29504
rect 23072 29492 23078 29504
rect 24857 29495 24915 29501
rect 24857 29492 24869 29495
rect 23072 29464 24869 29492
rect 23072 29452 23078 29464
rect 24857 29461 24869 29464
rect 24903 29492 24915 29495
rect 25682 29492 25688 29504
rect 24903 29464 25688 29492
rect 24903 29461 24915 29464
rect 24857 29455 24915 29461
rect 25682 29452 25688 29464
rect 25740 29452 25746 29504
rect 26068 29492 26096 29532
rect 26142 29520 26148 29572
rect 26200 29560 26206 29572
rect 26200 29532 26556 29560
rect 26200 29520 26206 29532
rect 26237 29495 26295 29501
rect 26237 29492 26249 29495
rect 26068 29464 26249 29492
rect 26237 29461 26249 29464
rect 26283 29461 26295 29495
rect 26528 29492 26556 29532
rect 26602 29520 26608 29572
rect 26660 29520 26666 29572
rect 27522 29520 27528 29572
rect 27580 29560 27586 29572
rect 30282 29560 30288 29572
rect 27580 29532 30288 29560
rect 27580 29520 27586 29532
rect 30282 29520 30288 29532
rect 30340 29520 30346 29572
rect 30742 29520 30748 29572
rect 30800 29520 30806 29572
rect 30834 29520 30840 29572
rect 30892 29560 30898 29572
rect 31404 29560 31432 29591
rect 30892 29532 31432 29560
rect 31680 29560 31708 29591
rect 32950 29588 32956 29600
rect 33008 29588 33014 29640
rect 31938 29560 31944 29572
rect 31680 29532 31944 29560
rect 30892 29520 30898 29532
rect 31938 29520 31944 29532
rect 31996 29520 32002 29572
rect 26697 29495 26755 29501
rect 26697 29492 26709 29495
rect 26528 29464 26709 29492
rect 26237 29455 26295 29461
rect 26697 29461 26709 29464
rect 26743 29461 26755 29495
rect 26697 29455 26755 29461
rect 27982 29452 27988 29504
rect 28040 29452 28046 29504
rect 28166 29452 28172 29504
rect 28224 29492 28230 29504
rect 28810 29492 28816 29504
rect 28224 29464 28816 29492
rect 28224 29452 28230 29464
rect 28810 29452 28816 29464
rect 28868 29492 28874 29504
rect 30926 29492 30932 29504
rect 28868 29464 30932 29492
rect 28868 29452 28874 29464
rect 30926 29452 30932 29464
rect 30984 29452 30990 29504
rect 31110 29452 31116 29504
rect 31168 29492 31174 29504
rect 31478 29492 31484 29504
rect 31168 29464 31484 29492
rect 31168 29452 31174 29464
rect 31478 29452 31484 29464
rect 31536 29452 31542 29504
rect 31570 29452 31576 29504
rect 31628 29452 31634 29504
rect 31846 29452 31852 29504
rect 31904 29452 31910 29504
rect 32306 29452 32312 29504
rect 32364 29452 32370 29504
rect 1104 29402 36432 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 36432 29402
rect 1104 29328 36432 29350
rect 4341 29291 4399 29297
rect 4341 29288 4353 29291
rect 1780 29260 4353 29288
rect 1302 29180 1308 29232
rect 1360 29220 1366 29232
rect 1780 29229 1808 29260
rect 4341 29257 4353 29260
rect 4387 29257 4399 29291
rect 4341 29251 4399 29257
rect 7742 29248 7748 29300
rect 7800 29288 7806 29300
rect 13265 29291 13323 29297
rect 13265 29288 13277 29291
rect 7800 29260 13277 29288
rect 7800 29248 7806 29260
rect 13265 29257 13277 29260
rect 13311 29257 13323 29291
rect 13265 29251 13323 29257
rect 16022 29248 16028 29300
rect 16080 29288 16086 29300
rect 16080 29260 18000 29288
rect 16080 29248 16086 29260
rect 1765 29223 1823 29229
rect 1765 29220 1777 29223
rect 1360 29192 1777 29220
rect 1360 29180 1366 29192
rect 1765 29189 1777 29192
rect 1811 29189 1823 29223
rect 1765 29183 1823 29189
rect 3050 29180 3056 29232
rect 3108 29180 3114 29232
rect 3602 29180 3608 29232
rect 3660 29220 3666 29232
rect 4249 29223 4307 29229
rect 3660 29192 3832 29220
rect 3660 29180 3666 29192
rect 3804 29161 3832 29192
rect 4249 29189 4261 29223
rect 4295 29220 4307 29223
rect 4798 29220 4804 29232
rect 4295 29192 4804 29220
rect 4295 29189 4307 29192
rect 4249 29183 4307 29189
rect 4798 29180 4804 29192
rect 4856 29180 4862 29232
rect 6454 29180 6460 29232
rect 6512 29220 6518 29232
rect 6512 29192 6960 29220
rect 6512 29180 6518 29192
rect 6932 29161 6960 29192
rect 7098 29180 7104 29232
rect 7156 29220 7162 29232
rect 7929 29223 7987 29229
rect 7156 29192 7328 29220
rect 7156 29180 7162 29192
rect 3789 29155 3847 29161
rect 3789 29121 3801 29155
rect 3835 29121 3847 29155
rect 3789 29115 3847 29121
rect 6825 29155 6883 29161
rect 6825 29121 6837 29155
rect 6871 29121 6883 29155
rect 6825 29115 6883 29121
rect 6917 29155 6975 29161
rect 6917 29121 6929 29155
rect 6963 29121 6975 29155
rect 6917 29115 6975 29121
rect 3513 29087 3571 29093
rect 3513 29053 3525 29087
rect 3559 29084 3571 29087
rect 3559 29056 3924 29084
rect 3559 29053 3571 29056
rect 3513 29047 3571 29053
rect 3896 29025 3924 29056
rect 4062 29044 4068 29096
rect 4120 29084 4126 29096
rect 4433 29087 4491 29093
rect 4433 29084 4445 29087
rect 4120 29056 4445 29084
rect 4120 29044 4126 29056
rect 4433 29053 4445 29056
rect 4479 29053 4491 29087
rect 4433 29047 4491 29053
rect 3881 29019 3939 29025
rect 3881 28985 3893 29019
rect 3927 28985 3939 29019
rect 3881 28979 3939 28985
rect 6840 29016 6868 29115
rect 7190 29112 7196 29164
rect 7248 29112 7254 29164
rect 7300 29152 7328 29192
rect 7929 29189 7941 29223
rect 7975 29220 7987 29223
rect 9398 29220 9404 29232
rect 7975 29192 9404 29220
rect 7975 29189 7987 29192
rect 7929 29183 7987 29189
rect 9398 29180 9404 29192
rect 9456 29180 9462 29232
rect 10229 29223 10287 29229
rect 10229 29189 10241 29223
rect 10275 29220 10287 29223
rect 10318 29220 10324 29232
rect 10275 29192 10324 29220
rect 10275 29189 10287 29192
rect 10229 29183 10287 29189
rect 10318 29180 10324 29192
rect 10376 29180 10382 29232
rect 10686 29180 10692 29232
rect 10744 29220 10750 29232
rect 14366 29220 14372 29232
rect 10744 29192 14372 29220
rect 10744 29180 10750 29192
rect 14366 29180 14372 29192
rect 14424 29180 14430 29232
rect 15286 29180 15292 29232
rect 15344 29220 15350 29232
rect 16390 29220 16396 29232
rect 15344 29192 16396 29220
rect 15344 29180 15350 29192
rect 16390 29180 16396 29192
rect 16448 29180 16454 29232
rect 16758 29180 16764 29232
rect 16816 29220 16822 29232
rect 16816 29195 17356 29220
rect 16816 29192 17371 29195
rect 16816 29180 16822 29192
rect 17313 29189 17371 29192
rect 7358 29155 7416 29161
rect 7358 29152 7370 29155
rect 7300 29124 7370 29152
rect 7358 29121 7370 29124
rect 7404 29121 7416 29155
rect 7358 29115 7416 29121
rect 7742 29112 7748 29164
rect 7800 29112 7806 29164
rect 8662 29112 8668 29164
rect 8720 29152 8726 29164
rect 9214 29152 9220 29164
rect 8720 29124 9220 29152
rect 8720 29112 8726 29124
rect 9214 29112 9220 29124
rect 9272 29112 9278 29164
rect 9582 29112 9588 29164
rect 9640 29112 9646 29164
rect 9950 29112 9956 29164
rect 10008 29112 10014 29164
rect 11790 29112 11796 29164
rect 11848 29152 11854 29164
rect 12069 29155 12127 29161
rect 12069 29152 12081 29155
rect 11848 29124 12081 29152
rect 11848 29112 11854 29124
rect 12069 29121 12081 29124
rect 12115 29121 12127 29155
rect 12069 29115 12127 29121
rect 12250 29112 12256 29164
rect 12308 29152 12314 29164
rect 12529 29155 12587 29161
rect 12529 29152 12541 29155
rect 12308 29124 12541 29152
rect 12308 29112 12314 29124
rect 12529 29121 12541 29124
rect 12575 29152 12587 29155
rect 12710 29152 12716 29164
rect 12575 29124 12716 29152
rect 12575 29121 12587 29124
rect 12529 29115 12587 29121
rect 12710 29112 12716 29124
rect 12768 29112 12774 29164
rect 12894 29112 12900 29164
rect 12952 29112 12958 29164
rect 13081 29155 13139 29161
rect 13081 29121 13093 29155
rect 13127 29152 13139 29155
rect 13262 29152 13268 29164
rect 13127 29124 13268 29152
rect 13127 29121 13139 29124
rect 13081 29115 13139 29121
rect 13262 29112 13268 29124
rect 13320 29152 13326 29164
rect 13320 29124 13584 29152
rect 13320 29112 13326 29124
rect 7466 29044 7472 29096
rect 7524 29044 7530 29096
rect 7561 29087 7619 29093
rect 7561 29053 7573 29087
rect 7607 29053 7619 29087
rect 7561 29047 7619 29053
rect 9309 29087 9367 29093
rect 9309 29053 9321 29087
rect 9355 29084 9367 29087
rect 9398 29084 9404 29096
rect 9355 29056 9404 29084
rect 9355 29053 9367 29056
rect 9309 29047 9367 29053
rect 7006 29016 7012 29028
rect 6840 28988 7012 29016
rect 2406 28908 2412 28960
rect 2464 28948 2470 28960
rect 5258 28948 5264 28960
rect 2464 28920 5264 28948
rect 2464 28908 2470 28920
rect 5258 28908 5264 28920
rect 5316 28908 5322 28960
rect 5350 28908 5356 28960
rect 5408 28948 5414 28960
rect 6840 28948 6868 28988
rect 7006 28976 7012 28988
rect 7064 29016 7070 29028
rect 7576 29016 7604 29047
rect 9398 29044 9404 29056
rect 9456 29044 9462 29096
rect 11146 29044 11152 29096
rect 11204 29084 11210 29096
rect 12621 29087 12679 29093
rect 11204 29056 12572 29084
rect 11204 29044 11210 29056
rect 8110 29016 8116 29028
rect 7064 28988 8116 29016
rect 7064 28976 7070 28988
rect 8110 28976 8116 28988
rect 8168 28976 8174 29028
rect 10042 28976 10048 29028
rect 10100 29016 10106 29028
rect 12161 29019 12219 29025
rect 10100 28988 12112 29016
rect 10100 28976 10106 28988
rect 5408 28920 6868 28948
rect 5408 28908 5414 28920
rect 9582 28908 9588 28960
rect 9640 28948 9646 28960
rect 11698 28948 11704 28960
rect 9640 28920 11704 28948
rect 9640 28908 9646 28920
rect 11698 28908 11704 28920
rect 11756 28908 11762 28960
rect 12084 28948 12112 28988
rect 12161 28985 12173 29019
rect 12207 29016 12219 29019
rect 12434 29016 12440 29028
rect 12207 28988 12440 29016
rect 12207 28985 12219 28988
rect 12161 28979 12219 28985
rect 12434 28976 12440 28988
rect 12492 28976 12498 29028
rect 12544 29016 12572 29056
rect 12621 29053 12633 29087
rect 12667 29084 12679 29087
rect 12802 29084 12808 29096
rect 12667 29056 12808 29084
rect 12667 29053 12679 29056
rect 12621 29047 12679 29053
rect 12802 29044 12808 29056
rect 12860 29044 12866 29096
rect 12912 29016 12940 29112
rect 13170 29044 13176 29096
rect 13228 29044 13234 29096
rect 13446 29044 13452 29096
rect 13504 29044 13510 29096
rect 13556 29084 13584 29124
rect 13630 29112 13636 29164
rect 13688 29112 13694 29164
rect 14001 29155 14059 29161
rect 14001 29121 14013 29155
rect 14047 29152 14059 29155
rect 14182 29152 14188 29164
rect 14047 29124 14188 29152
rect 14047 29121 14059 29124
rect 14001 29115 14059 29121
rect 13814 29084 13820 29096
rect 13556 29056 13820 29084
rect 13814 29044 13820 29056
rect 13872 29084 13878 29096
rect 13909 29087 13967 29093
rect 13909 29084 13921 29087
rect 13872 29056 13921 29084
rect 13872 29044 13878 29056
rect 13909 29053 13921 29056
rect 13955 29053 13967 29087
rect 13909 29047 13967 29053
rect 14016 29016 14044 29115
rect 14182 29112 14188 29124
rect 14240 29112 14246 29164
rect 14458 29112 14464 29164
rect 14516 29112 14522 29164
rect 15105 29155 15163 29161
rect 15105 29121 15117 29155
rect 15151 29152 15163 29155
rect 15746 29152 15752 29164
rect 15151 29124 15752 29152
rect 15151 29121 15163 29124
rect 15105 29115 15163 29121
rect 15746 29112 15752 29124
rect 15804 29112 15810 29164
rect 16850 29112 16856 29164
rect 16908 29112 16914 29164
rect 17129 29155 17187 29161
rect 17129 29152 17141 29155
rect 16960 29124 17141 29152
rect 14366 29044 14372 29096
rect 14424 29084 14430 29096
rect 14737 29087 14795 29093
rect 14737 29084 14749 29087
rect 14424 29056 14749 29084
rect 14424 29044 14430 29056
rect 14737 29053 14749 29056
rect 14783 29053 14795 29087
rect 14737 29047 14795 29053
rect 15286 29044 15292 29096
rect 15344 29084 15350 29096
rect 15470 29084 15476 29096
rect 15344 29056 15476 29084
rect 15344 29044 15350 29056
rect 15470 29044 15476 29056
rect 15528 29044 15534 29096
rect 15562 29044 15568 29096
rect 15620 29044 15626 29096
rect 15654 29044 15660 29096
rect 15712 29044 15718 29096
rect 15838 29044 15844 29096
rect 15896 29084 15902 29096
rect 16025 29087 16083 29093
rect 16025 29084 16037 29087
rect 15896 29056 16037 29084
rect 15896 29044 15902 29056
rect 16025 29053 16037 29056
rect 16071 29084 16083 29087
rect 16206 29084 16212 29096
rect 16071 29056 16212 29084
rect 16071 29053 16083 29056
rect 16025 29047 16083 29053
rect 16206 29044 16212 29056
rect 16264 29044 16270 29096
rect 16960 29084 16988 29124
rect 17129 29121 17141 29124
rect 17175 29152 17187 29155
rect 17218 29152 17224 29164
rect 17175 29124 17224 29152
rect 17175 29121 17187 29124
rect 17129 29115 17187 29121
rect 17218 29112 17224 29124
rect 17276 29112 17282 29164
rect 17313 29155 17325 29189
rect 17359 29155 17371 29189
rect 17313 29149 17371 29155
rect 17589 29155 17647 29161
rect 17589 29121 17601 29155
rect 17635 29152 17647 29155
rect 17770 29152 17776 29164
rect 17635 29124 17776 29152
rect 17635 29121 17647 29124
rect 17589 29115 17647 29121
rect 17770 29112 17776 29124
rect 17828 29112 17834 29164
rect 17865 29155 17923 29161
rect 17865 29121 17877 29155
rect 17911 29152 17923 29155
rect 17972 29152 18000 29260
rect 18506 29248 18512 29300
rect 18564 29288 18570 29300
rect 18785 29291 18843 29297
rect 18785 29288 18797 29291
rect 18564 29260 18797 29288
rect 18564 29248 18570 29260
rect 18785 29257 18797 29260
rect 18831 29257 18843 29291
rect 18785 29251 18843 29257
rect 19058 29248 19064 29300
rect 19116 29288 19122 29300
rect 20165 29291 20223 29297
rect 20165 29288 20177 29291
rect 19116 29260 20177 29288
rect 19116 29248 19122 29260
rect 20165 29257 20177 29260
rect 20211 29257 20223 29291
rect 21634 29288 21640 29300
rect 20165 29251 20223 29257
rect 20456 29260 21640 29288
rect 20254 29220 20260 29232
rect 18524 29192 20260 29220
rect 17911 29124 18000 29152
rect 17911 29121 17923 29124
rect 17865 29115 17923 29121
rect 18046 29112 18052 29164
rect 18104 29152 18110 29164
rect 18524 29161 18552 29192
rect 20254 29180 20260 29192
rect 20312 29180 20318 29232
rect 18417 29155 18475 29161
rect 18417 29152 18429 29155
rect 18104 29124 18429 29152
rect 18104 29112 18110 29124
rect 18417 29121 18429 29124
rect 18463 29121 18475 29155
rect 18417 29115 18475 29121
rect 18509 29155 18567 29161
rect 18509 29121 18521 29155
rect 18555 29121 18567 29155
rect 18509 29115 18567 29121
rect 18601 29155 18659 29161
rect 18601 29121 18613 29155
rect 18647 29152 18659 29155
rect 18966 29152 18972 29164
rect 18647 29124 18972 29152
rect 18647 29121 18659 29124
rect 18601 29115 18659 29121
rect 18966 29112 18972 29124
rect 19024 29112 19030 29164
rect 20456 29161 20484 29260
rect 21634 29248 21640 29260
rect 21692 29248 21698 29300
rect 21818 29248 21824 29300
rect 21876 29288 21882 29300
rect 21876 29260 22600 29288
rect 21876 29248 21882 29260
rect 20901 29223 20959 29229
rect 20901 29220 20913 29223
rect 20548 29192 20913 29220
rect 20548 29161 20576 29192
rect 20901 29189 20913 29192
rect 20947 29189 20959 29223
rect 22281 29223 22339 29229
rect 22281 29220 22293 29223
rect 20901 29183 20959 29189
rect 21100 29192 22293 29220
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29121 20499 29155
rect 20441 29115 20499 29121
rect 20533 29155 20591 29161
rect 20533 29121 20545 29155
rect 20579 29121 20591 29155
rect 20533 29115 20591 29121
rect 20622 29112 20628 29164
rect 20680 29112 20686 29164
rect 20806 29112 20812 29164
rect 20864 29112 20870 29164
rect 20990 29112 20996 29164
rect 21048 29152 21054 29164
rect 21100 29161 21128 29192
rect 22281 29189 22293 29192
rect 22327 29189 22339 29223
rect 22281 29183 22339 29189
rect 21085 29155 21143 29161
rect 21085 29152 21097 29155
rect 21048 29124 21097 29152
rect 21048 29112 21054 29124
rect 21085 29121 21097 29124
rect 21131 29121 21143 29155
rect 21085 29115 21143 29121
rect 21174 29112 21180 29164
rect 21232 29112 21238 29164
rect 21450 29112 21456 29164
rect 21508 29112 21514 29164
rect 21634 29112 21640 29164
rect 21692 29152 21698 29164
rect 22572 29161 22600 29260
rect 22646 29248 22652 29300
rect 22704 29248 22710 29300
rect 22738 29248 22744 29300
rect 22796 29288 22802 29300
rect 23382 29288 23388 29300
rect 22796 29260 23388 29288
rect 22796 29248 22802 29260
rect 23382 29248 23388 29260
rect 23440 29248 23446 29300
rect 24946 29288 24952 29300
rect 23768 29260 24952 29288
rect 22005 29155 22063 29161
rect 22005 29152 22017 29155
rect 21692 29124 22017 29152
rect 21692 29112 21698 29124
rect 22005 29121 22017 29124
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 22557 29155 22615 29161
rect 22557 29121 22569 29155
rect 22603 29121 22615 29155
rect 22557 29115 22615 29121
rect 22830 29112 22836 29164
rect 22888 29112 22894 29164
rect 23201 29155 23259 29161
rect 23201 29121 23213 29155
rect 23247 29152 23259 29155
rect 23290 29152 23296 29164
rect 23247 29124 23296 29152
rect 23247 29121 23259 29124
rect 23201 29115 23259 29121
rect 23290 29112 23296 29124
rect 23348 29112 23354 29164
rect 23768 29161 23796 29260
rect 24946 29248 24952 29260
rect 25004 29248 25010 29300
rect 25547 29291 25605 29297
rect 25547 29257 25559 29291
rect 25593 29288 25605 29291
rect 26602 29288 26608 29300
rect 25593 29260 26608 29288
rect 25593 29257 25605 29260
rect 25547 29251 25605 29257
rect 26602 29248 26608 29260
rect 26660 29248 26666 29300
rect 26786 29248 26792 29300
rect 26844 29288 26850 29300
rect 29178 29288 29184 29300
rect 26844 29260 29184 29288
rect 26844 29248 26850 29260
rect 29178 29248 29184 29260
rect 29236 29248 29242 29300
rect 29457 29291 29515 29297
rect 29457 29257 29469 29291
rect 29503 29288 29515 29291
rect 32674 29288 32680 29300
rect 29503 29260 32680 29288
rect 29503 29257 29515 29260
rect 29457 29251 29515 29257
rect 32674 29248 32680 29260
rect 32732 29248 32738 29300
rect 24486 29180 24492 29232
rect 24544 29180 24550 29232
rect 28166 29180 28172 29232
rect 28224 29220 28230 29232
rect 28224 29192 28580 29220
rect 28224 29180 28230 29192
rect 23753 29155 23811 29161
rect 23753 29121 23765 29155
rect 23799 29121 23811 29155
rect 23753 29115 23811 29121
rect 16316 29056 16988 29084
rect 12544 28988 12940 29016
rect 13004 28988 14044 29016
rect 13004 28948 13032 28988
rect 14274 28976 14280 29028
rect 14332 28976 14338 29028
rect 14918 28976 14924 29028
rect 14976 28976 14982 29028
rect 15378 28976 15384 29028
rect 15436 28976 15442 29028
rect 15672 29016 15700 29044
rect 16316 29016 16344 29056
rect 17034 29044 17040 29096
rect 17092 29044 17098 29096
rect 17144 29056 17632 29084
rect 15672 28988 16344 29016
rect 16945 29019 17003 29025
rect 16945 28985 16957 29019
rect 16991 29016 17003 29019
rect 17144 29016 17172 29056
rect 16991 28988 17172 29016
rect 16991 28985 17003 28988
rect 16945 28979 17003 28985
rect 17218 28976 17224 29028
rect 17276 29016 17282 29028
rect 17405 29019 17463 29025
rect 17405 29016 17417 29019
rect 17276 28988 17417 29016
rect 17276 28976 17282 28988
rect 17405 28985 17417 28988
rect 17451 28985 17463 29019
rect 17604 29016 17632 29056
rect 17678 29044 17684 29096
rect 17736 29084 17742 29096
rect 21468 29084 21496 29112
rect 22189 29087 22247 29093
rect 17736 29056 22094 29084
rect 17736 29044 17742 29056
rect 17788 29025 17816 29056
rect 17773 29019 17831 29025
rect 17604 28988 17724 29016
rect 17405 28979 17463 28985
rect 12084 28920 13032 28948
rect 14645 28951 14703 28957
rect 14645 28917 14657 28951
rect 14691 28948 14703 28951
rect 14826 28948 14832 28960
rect 14691 28920 14832 28948
rect 14691 28917 14703 28920
rect 14645 28911 14703 28917
rect 14826 28908 14832 28920
rect 14884 28908 14890 28960
rect 16574 28908 16580 28960
rect 16632 28948 16638 28960
rect 16669 28951 16727 28957
rect 16669 28948 16681 28951
rect 16632 28920 16681 28948
rect 16632 28908 16638 28920
rect 16669 28917 16681 28920
rect 16715 28917 16727 28951
rect 17696 28948 17724 28988
rect 17773 28985 17785 29019
rect 17819 28985 17831 29019
rect 18046 29016 18052 29028
rect 17773 28979 17831 28985
rect 17880 28988 18052 29016
rect 17880 28948 17908 28988
rect 18046 28976 18052 28988
rect 18104 28976 18110 29028
rect 18233 29019 18291 29025
rect 18233 28985 18245 29019
rect 18279 29016 18291 29019
rect 20162 29016 20168 29028
rect 18279 28988 20168 29016
rect 18279 28985 18291 28988
rect 18233 28979 18291 28985
rect 20162 28976 20168 28988
rect 20220 28976 20226 29028
rect 21358 28976 21364 29028
rect 21416 28976 21422 29028
rect 22066 29016 22094 29056
rect 22189 29053 22201 29087
rect 22235 29084 22247 29087
rect 22278 29084 22284 29096
rect 22235 29056 22284 29084
rect 22235 29053 22247 29056
rect 22189 29047 22247 29053
rect 22278 29044 22284 29056
rect 22336 29084 22342 29096
rect 22922 29084 22928 29096
rect 22336 29056 22928 29084
rect 22336 29044 22342 29056
rect 22922 29044 22928 29056
rect 22980 29044 22986 29096
rect 23198 29016 23204 29028
rect 22066 28988 23204 29016
rect 23198 28976 23204 28988
rect 23256 28976 23262 29028
rect 23290 28976 23296 29028
rect 23348 29016 23354 29028
rect 23569 29019 23627 29025
rect 23569 29016 23581 29019
rect 23348 28988 23581 29016
rect 23348 28976 23354 28988
rect 23569 28985 23581 28988
rect 23615 28985 23627 29019
rect 23569 28979 23627 28985
rect 17696 28920 17908 28948
rect 16669 28911 16727 28917
rect 21818 28908 21824 28960
rect 21876 28908 21882 28960
rect 21910 28908 21916 28960
rect 21968 28948 21974 28960
rect 22005 28951 22063 28957
rect 22005 28948 22017 28951
rect 21968 28920 22017 28948
rect 21968 28908 21974 28920
rect 22005 28917 22017 28920
rect 22051 28917 22063 28951
rect 22005 28911 22063 28917
rect 23382 28908 23388 28960
rect 23440 28948 23446 28960
rect 23768 28948 23796 29115
rect 26142 29112 26148 29164
rect 26200 29152 26206 29164
rect 26513 29155 26571 29161
rect 26513 29152 26525 29155
rect 26200 29124 26525 29152
rect 26200 29112 26206 29124
rect 26513 29121 26525 29124
rect 26559 29121 26571 29155
rect 26513 29115 26571 29121
rect 26694 29112 26700 29164
rect 26752 29152 26758 29164
rect 27522 29152 27528 29164
rect 26752 29124 27528 29152
rect 26752 29112 26758 29124
rect 27522 29112 27528 29124
rect 27580 29112 27586 29164
rect 27798 29112 27804 29164
rect 27856 29152 27862 29164
rect 28258 29152 28264 29164
rect 27856 29124 28264 29152
rect 27856 29112 27862 29124
rect 28258 29112 28264 29124
rect 28316 29112 28322 29164
rect 28552 29161 28580 29192
rect 29564 29192 29960 29220
rect 29564 29164 29592 29192
rect 28537 29155 28595 29161
rect 28537 29121 28549 29155
rect 28583 29121 28595 29155
rect 28537 29115 28595 29121
rect 28721 29155 28779 29161
rect 28721 29121 28733 29155
rect 28767 29121 28779 29155
rect 28721 29115 28779 29121
rect 28905 29155 28963 29161
rect 28905 29121 28917 29155
rect 28951 29152 28963 29155
rect 28994 29152 29000 29164
rect 28951 29124 29000 29152
rect 28951 29121 28963 29124
rect 28905 29115 28963 29121
rect 24121 29087 24179 29093
rect 24121 29053 24133 29087
rect 24167 29084 24179 29087
rect 25590 29084 25596 29096
rect 24167 29056 25596 29084
rect 24167 29053 24179 29056
rect 24121 29047 24179 29053
rect 25590 29044 25596 29056
rect 25648 29044 25654 29096
rect 26237 29087 26295 29093
rect 26237 29053 26249 29087
rect 26283 29084 26295 29087
rect 26602 29084 26608 29096
rect 26283 29056 26608 29084
rect 26283 29053 26295 29056
rect 26237 29047 26295 29053
rect 26602 29044 26608 29056
rect 26660 29044 26666 29096
rect 26878 29044 26884 29096
rect 26936 29084 26942 29096
rect 27065 29087 27123 29093
rect 27065 29084 27077 29087
rect 26936 29056 27077 29084
rect 26936 29044 26942 29056
rect 27065 29053 27077 29056
rect 27111 29053 27123 29087
rect 27065 29047 27123 29053
rect 27157 29087 27215 29093
rect 27157 29053 27169 29087
rect 27203 29084 27215 29087
rect 28736 29084 28764 29115
rect 28994 29112 29000 29124
rect 29052 29152 29058 29164
rect 29365 29155 29423 29161
rect 29365 29152 29377 29155
rect 29052 29124 29377 29152
rect 29052 29112 29058 29124
rect 29365 29121 29377 29124
rect 29411 29121 29423 29155
rect 29365 29115 29423 29121
rect 29546 29112 29552 29164
rect 29604 29112 29610 29164
rect 29932 29161 29960 29192
rect 30374 29180 30380 29232
rect 30432 29180 30438 29232
rect 30742 29180 30748 29232
rect 30800 29220 30806 29232
rect 30926 29220 30932 29232
rect 30800 29192 30932 29220
rect 30800 29180 30806 29192
rect 30926 29180 30932 29192
rect 30984 29180 30990 29232
rect 36170 29220 36176 29232
rect 31036 29192 31340 29220
rect 29825 29155 29883 29161
rect 29825 29121 29837 29155
rect 29871 29121 29883 29155
rect 29825 29115 29883 29121
rect 29917 29155 29975 29161
rect 29917 29121 29929 29155
rect 29963 29121 29975 29155
rect 29917 29115 29975 29121
rect 29840 29084 29868 29115
rect 30650 29112 30656 29164
rect 30708 29152 30714 29164
rect 31036 29152 31064 29192
rect 30708 29124 31064 29152
rect 31205 29155 31263 29161
rect 30708 29112 30714 29124
rect 31205 29121 31217 29155
rect 31251 29121 31263 29155
rect 31205 29115 31263 29121
rect 27203 29056 30144 29084
rect 27203 29053 27215 29056
rect 27157 29047 27215 29053
rect 27080 29016 27108 29047
rect 27706 29016 27712 29028
rect 27080 28988 27712 29016
rect 27706 28976 27712 28988
rect 27764 29016 27770 29028
rect 28353 29019 28411 29025
rect 28353 29016 28365 29019
rect 27764 28988 28365 29016
rect 27764 28976 27770 28988
rect 28353 28985 28365 28988
rect 28399 28985 28411 29019
rect 28353 28979 28411 28985
rect 28442 28976 28448 29028
rect 28500 29016 28506 29028
rect 28500 28988 29224 29016
rect 28500 28976 28506 28988
rect 23440 28920 23796 28948
rect 23440 28908 23446 28920
rect 26510 28908 26516 28960
rect 26568 28948 26574 28960
rect 26878 28948 26884 28960
rect 26568 28920 26884 28948
rect 26568 28908 26574 28920
rect 26878 28908 26884 28920
rect 26936 28908 26942 28960
rect 28074 28908 28080 28960
rect 28132 28908 28138 28960
rect 28534 28908 28540 28960
rect 28592 28948 28598 28960
rect 28721 28951 28779 28957
rect 28721 28948 28733 28951
rect 28592 28920 28733 28948
rect 28592 28908 28598 28920
rect 28721 28917 28733 28920
rect 28767 28917 28779 28951
rect 29196 28948 29224 28988
rect 30006 28976 30012 29028
rect 30064 28976 30070 29028
rect 30116 29016 30144 29056
rect 30466 29044 30472 29096
rect 30524 29084 30530 29096
rect 30837 29087 30895 29093
rect 30837 29084 30849 29087
rect 30524 29056 30849 29084
rect 30524 29044 30530 29056
rect 30837 29053 30849 29056
rect 30883 29084 30895 29087
rect 31220 29084 31248 29115
rect 30883 29056 31248 29084
rect 31312 29084 31340 29192
rect 31588 29192 36176 29220
rect 31478 29112 31484 29164
rect 31536 29152 31542 29164
rect 31588 29161 31616 29192
rect 36170 29180 36176 29192
rect 36228 29180 36234 29232
rect 31573 29155 31631 29161
rect 31573 29152 31585 29155
rect 31536 29124 31585 29152
rect 31536 29112 31542 29124
rect 31573 29121 31585 29124
rect 31619 29121 31631 29155
rect 31573 29115 31631 29121
rect 31662 29112 31668 29164
rect 31720 29152 31726 29164
rect 33778 29152 33784 29164
rect 31720 29124 33784 29152
rect 31720 29112 31726 29124
rect 33778 29112 33784 29124
rect 33836 29112 33842 29164
rect 35802 29112 35808 29164
rect 35860 29112 35866 29164
rect 31312 29056 32076 29084
rect 30883 29053 30895 29056
rect 30837 29047 30895 29053
rect 31938 29016 31944 29028
rect 30116 28988 31944 29016
rect 31938 28976 31944 28988
rect 31996 28976 32002 29028
rect 30650 28948 30656 28960
rect 29196 28920 30656 28948
rect 28721 28911 28779 28917
rect 30650 28908 30656 28920
rect 30708 28908 30714 28960
rect 30834 28908 30840 28960
rect 30892 28948 30898 28960
rect 31021 28951 31079 28957
rect 31021 28948 31033 28951
rect 30892 28920 31033 28948
rect 30892 28908 30898 28920
rect 31021 28917 31033 28920
rect 31067 28917 31079 28951
rect 32048 28948 32076 29056
rect 34514 29044 34520 29096
rect 34572 29084 34578 29096
rect 34701 29087 34759 29093
rect 34701 29084 34713 29087
rect 34572 29056 34713 29084
rect 34572 29044 34578 29056
rect 34701 29053 34713 29056
rect 34747 29053 34759 29087
rect 34701 29047 34759 29053
rect 34790 29044 34796 29096
rect 34848 29084 34854 29096
rect 34977 29087 35035 29093
rect 34977 29084 34989 29087
rect 34848 29056 34989 29084
rect 34848 29044 34854 29056
rect 34977 29053 34989 29056
rect 35023 29053 35035 29087
rect 34977 29047 35035 29053
rect 35618 28976 35624 29028
rect 35676 28976 35682 29028
rect 35802 28948 35808 28960
rect 32048 28920 35808 28948
rect 31021 28911 31079 28917
rect 35802 28908 35808 28920
rect 35860 28908 35866 28960
rect 1104 28858 36432 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 36432 28858
rect 1104 28784 36432 28806
rect 5810 28744 5816 28756
rect 4172 28716 5816 28744
rect 1302 28568 1308 28620
rect 1360 28608 1366 28620
rect 1581 28611 1639 28617
rect 1581 28608 1593 28611
rect 1360 28580 1593 28608
rect 1360 28568 1366 28580
rect 1581 28577 1593 28580
rect 1627 28577 1639 28611
rect 1581 28571 1639 28577
rect 1596 28404 1624 28571
rect 3602 28568 3608 28620
rect 3660 28568 3666 28620
rect 3973 28543 4031 28549
rect 3973 28509 3985 28543
rect 4019 28540 4031 28543
rect 4172 28540 4200 28716
rect 5810 28704 5816 28716
rect 5868 28704 5874 28756
rect 6914 28704 6920 28756
rect 6972 28744 6978 28756
rect 7929 28747 7987 28753
rect 7929 28744 7941 28747
rect 6972 28716 7941 28744
rect 6972 28704 6978 28716
rect 7929 28713 7941 28716
rect 7975 28713 7987 28747
rect 7929 28707 7987 28713
rect 8297 28747 8355 28753
rect 8297 28713 8309 28747
rect 8343 28744 8355 28747
rect 8570 28744 8576 28756
rect 8343 28716 8576 28744
rect 8343 28713 8355 28716
rect 8297 28707 8355 28713
rect 8570 28704 8576 28716
rect 8628 28704 8634 28756
rect 9493 28747 9551 28753
rect 9493 28713 9505 28747
rect 9539 28744 9551 28747
rect 9950 28744 9956 28756
rect 9539 28716 9956 28744
rect 9539 28713 9551 28716
rect 9493 28707 9551 28713
rect 9950 28704 9956 28716
rect 10008 28704 10014 28756
rect 10134 28704 10140 28756
rect 10192 28744 10198 28756
rect 11146 28744 11152 28756
rect 10192 28716 11152 28744
rect 10192 28704 10198 28716
rect 11146 28704 11152 28716
rect 11204 28704 11210 28756
rect 15010 28704 15016 28756
rect 15068 28744 15074 28756
rect 15286 28744 15292 28756
rect 15068 28716 15292 28744
rect 15068 28704 15074 28716
rect 15286 28704 15292 28716
rect 15344 28704 15350 28756
rect 15746 28704 15752 28756
rect 15804 28704 15810 28756
rect 16482 28704 16488 28756
rect 16540 28744 16546 28756
rect 19242 28744 19248 28756
rect 16540 28716 19248 28744
rect 16540 28704 16546 28716
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 20809 28747 20867 28753
rect 20809 28713 20821 28747
rect 20855 28744 20867 28747
rect 21174 28744 21180 28756
rect 20855 28716 21180 28744
rect 20855 28713 20867 28716
rect 20809 28707 20867 28713
rect 21174 28704 21180 28716
rect 21232 28704 21238 28756
rect 21545 28747 21603 28753
rect 21545 28713 21557 28747
rect 21591 28744 21603 28747
rect 22278 28744 22284 28756
rect 21591 28716 22284 28744
rect 21591 28713 21603 28716
rect 21545 28707 21603 28713
rect 22278 28704 22284 28716
rect 22336 28704 22342 28756
rect 24394 28744 24400 28756
rect 23400 28716 24400 28744
rect 5537 28679 5595 28685
rect 5537 28645 5549 28679
rect 5583 28645 5595 28679
rect 5537 28639 5595 28645
rect 4985 28611 5043 28617
rect 4985 28577 4997 28611
rect 5031 28608 5043 28611
rect 5350 28608 5356 28620
rect 5031 28580 5356 28608
rect 5031 28577 5043 28580
rect 4985 28571 5043 28577
rect 5350 28568 5356 28580
rect 5408 28568 5414 28620
rect 5552 28608 5580 28639
rect 6270 28636 6276 28688
rect 6328 28636 6334 28688
rect 7098 28636 7104 28688
rect 7156 28676 7162 28688
rect 7466 28676 7472 28688
rect 7156 28648 7472 28676
rect 7156 28636 7162 28648
rect 7466 28636 7472 28648
rect 7524 28676 7530 28688
rect 7524 28648 7696 28676
rect 7524 28636 7530 28648
rect 5552 28580 5856 28608
rect 4019 28512 4200 28540
rect 4249 28543 4307 28549
rect 4019 28509 4031 28512
rect 3973 28503 4031 28509
rect 4249 28509 4261 28543
rect 4295 28509 4307 28543
rect 4249 28503 4307 28509
rect 5629 28543 5687 28549
rect 5629 28509 5641 28543
rect 5675 28509 5687 28543
rect 5629 28503 5687 28509
rect 2774 28432 2780 28484
rect 2832 28432 2838 28484
rect 3329 28475 3387 28481
rect 3329 28441 3341 28475
rect 3375 28472 3387 28475
rect 3789 28475 3847 28481
rect 3789 28472 3801 28475
rect 3375 28444 3801 28472
rect 3375 28441 3387 28444
rect 3329 28435 3387 28441
rect 3789 28441 3801 28444
rect 3835 28441 3847 28475
rect 3789 28435 3847 28441
rect 4062 28432 4068 28484
rect 4120 28472 4126 28484
rect 4264 28472 4292 28503
rect 4120 28444 4292 28472
rect 5169 28475 5227 28481
rect 4120 28432 4126 28444
rect 5169 28441 5181 28475
rect 5215 28472 5227 28475
rect 5258 28472 5264 28484
rect 5215 28444 5264 28472
rect 5215 28441 5227 28444
rect 5169 28435 5227 28441
rect 5258 28432 5264 28444
rect 5316 28432 5322 28484
rect 5644 28472 5672 28503
rect 5718 28500 5724 28552
rect 5776 28500 5782 28552
rect 5828 28540 5856 28580
rect 7558 28568 7564 28620
rect 7616 28568 7622 28620
rect 7668 28608 7696 28648
rect 7742 28636 7748 28688
rect 7800 28676 7806 28688
rect 8113 28679 8171 28685
rect 8113 28676 8125 28679
rect 7800 28648 8125 28676
rect 7800 28636 7806 28648
rect 8113 28645 8125 28648
rect 8159 28645 8171 28679
rect 8113 28639 8171 28645
rect 9214 28636 9220 28688
rect 9272 28676 9278 28688
rect 9272 28648 9628 28676
rect 9272 28636 9278 28648
rect 7837 28611 7895 28617
rect 7837 28608 7849 28611
rect 7668 28580 7849 28608
rect 7837 28577 7849 28580
rect 7883 28577 7895 28611
rect 7837 28571 7895 28577
rect 7926 28568 7932 28620
rect 7984 28608 7990 28620
rect 7984 28580 9352 28608
rect 7984 28568 7990 28580
rect 6031 28543 6089 28549
rect 6031 28540 6043 28543
rect 5828 28512 6043 28540
rect 6031 28509 6043 28512
rect 6077 28509 6089 28543
rect 6031 28503 6089 28509
rect 6454 28500 6460 28552
rect 6512 28500 6518 28552
rect 6549 28543 6607 28549
rect 6549 28509 6561 28543
rect 6595 28540 6607 28543
rect 7006 28540 7012 28552
rect 6595 28512 7012 28540
rect 6595 28509 6607 28512
rect 6549 28503 6607 28509
rect 7006 28500 7012 28512
rect 7064 28500 7070 28552
rect 7282 28500 7288 28552
rect 7340 28500 7346 28552
rect 7374 28500 7380 28552
rect 7432 28500 7438 28552
rect 8496 28549 8524 28580
rect 7653 28543 7711 28549
rect 7653 28509 7665 28543
rect 7699 28540 7711 28543
rect 7745 28543 7803 28549
rect 7745 28540 7757 28543
rect 7699 28512 7757 28540
rect 7699 28509 7711 28512
rect 7653 28503 7711 28509
rect 7745 28509 7757 28512
rect 7791 28540 7803 28543
rect 8205 28543 8263 28549
rect 8205 28540 8217 28543
rect 7791 28512 8217 28540
rect 7791 28509 7803 28512
rect 7745 28503 7803 28509
rect 8205 28509 8217 28512
rect 8251 28509 8263 28543
rect 8205 28503 8263 28509
rect 8481 28543 8539 28549
rect 8481 28509 8493 28543
rect 8527 28509 8539 28543
rect 8481 28503 8539 28509
rect 8573 28543 8631 28549
rect 8573 28509 8585 28543
rect 8619 28540 8631 28543
rect 8662 28540 8668 28552
rect 8619 28512 8668 28540
rect 8619 28509 8631 28512
rect 8573 28503 8631 28509
rect 7392 28472 7420 28500
rect 7926 28472 7932 28484
rect 5644 28444 6776 28472
rect 7392 28444 7932 28472
rect 6748 28416 6776 28444
rect 7926 28432 7932 28444
rect 7984 28432 7990 28484
rect 8220 28472 8248 28503
rect 8662 28500 8668 28512
rect 8720 28500 8726 28552
rect 9214 28500 9220 28552
rect 9272 28500 9278 28552
rect 9232 28472 9260 28500
rect 8220 28444 9260 28472
rect 9324 28472 9352 28580
rect 9398 28500 9404 28552
rect 9456 28500 9462 28552
rect 9600 28472 9628 28648
rect 9766 28636 9772 28688
rect 9824 28676 9830 28688
rect 10226 28676 10232 28688
rect 9824 28648 10232 28676
rect 9824 28636 9830 28648
rect 9968 28617 9996 28648
rect 10226 28636 10232 28648
rect 10284 28636 10290 28688
rect 10318 28636 10324 28688
rect 10376 28676 10382 28688
rect 14093 28679 14151 28685
rect 14093 28676 14105 28679
rect 10376 28648 14105 28676
rect 10376 28636 10382 28648
rect 14093 28645 14105 28648
rect 14139 28676 14151 28679
rect 15194 28676 15200 28688
rect 14139 28648 15200 28676
rect 14139 28645 14151 28648
rect 14093 28639 14151 28645
rect 15194 28636 15200 28648
rect 15252 28636 15258 28688
rect 16577 28679 16635 28685
rect 16577 28645 16589 28679
rect 16623 28676 16635 28679
rect 16850 28676 16856 28688
rect 16623 28648 16856 28676
rect 16623 28645 16635 28648
rect 16577 28639 16635 28645
rect 16850 28636 16856 28648
rect 16908 28636 16914 28688
rect 21683 28679 21741 28685
rect 18524 28648 21036 28676
rect 9953 28611 10011 28617
rect 9953 28577 9965 28611
rect 9999 28577 10011 28611
rect 12710 28608 12716 28620
rect 9953 28571 10011 28577
rect 10060 28580 12716 28608
rect 9674 28500 9680 28552
rect 9732 28500 9738 28552
rect 9766 28500 9772 28552
rect 9824 28500 9830 28552
rect 10060 28549 10088 28580
rect 10045 28543 10103 28549
rect 10045 28509 10057 28543
rect 10091 28509 10103 28543
rect 10045 28503 10103 28509
rect 10318 28500 10324 28552
rect 10376 28500 10382 28552
rect 10413 28543 10471 28549
rect 10413 28509 10425 28543
rect 10459 28540 10471 28543
rect 10594 28540 10600 28552
rect 10459 28512 10600 28540
rect 10459 28509 10471 28512
rect 10413 28503 10471 28509
rect 10594 28500 10600 28512
rect 10652 28500 10658 28552
rect 10888 28549 10916 28580
rect 12710 28568 12716 28580
rect 12768 28568 12774 28620
rect 12894 28568 12900 28620
rect 12952 28568 12958 28620
rect 16758 28608 16764 28620
rect 14660 28580 15240 28608
rect 10873 28543 10931 28549
rect 10873 28509 10885 28543
rect 10919 28509 10931 28543
rect 10873 28503 10931 28509
rect 10962 28500 10968 28552
rect 11020 28540 11026 28552
rect 11057 28543 11115 28549
rect 11057 28540 11069 28543
rect 11020 28512 11069 28540
rect 11020 28500 11026 28512
rect 11057 28509 11069 28512
rect 11103 28509 11115 28543
rect 11057 28503 11115 28509
rect 11790 28500 11796 28552
rect 11848 28540 11854 28552
rect 12069 28543 12127 28549
rect 12069 28540 12081 28543
rect 11848 28512 12081 28540
rect 11848 28500 11854 28512
rect 12069 28509 12081 28512
rect 12115 28509 12127 28543
rect 12069 28503 12127 28509
rect 10137 28475 10195 28481
rect 10137 28472 10149 28475
rect 9324 28444 9444 28472
rect 9600 28444 10149 28472
rect 4157 28407 4215 28413
rect 4157 28404 4169 28407
rect 1596 28376 4169 28404
rect 4157 28373 4169 28376
rect 4203 28373 4215 28407
rect 4157 28367 4215 28373
rect 4798 28364 4804 28416
rect 4856 28404 4862 28416
rect 5077 28407 5135 28413
rect 5077 28404 5089 28407
rect 4856 28376 5089 28404
rect 4856 28364 4862 28376
rect 5077 28373 5089 28376
rect 5123 28373 5135 28407
rect 5077 28367 5135 28373
rect 6730 28364 6736 28416
rect 6788 28364 6794 28416
rect 7101 28407 7159 28413
rect 7101 28373 7113 28407
rect 7147 28404 7159 28407
rect 7282 28404 7288 28416
rect 7147 28376 7288 28404
rect 7147 28373 7159 28376
rect 7101 28367 7159 28373
rect 7282 28364 7288 28376
rect 7340 28364 7346 28416
rect 8757 28407 8815 28413
rect 8757 28373 8769 28407
rect 8803 28404 8815 28407
rect 9122 28404 9128 28416
rect 8803 28376 9128 28404
rect 8803 28373 8815 28376
rect 8757 28367 8815 28373
rect 9122 28364 9128 28376
rect 9180 28364 9186 28416
rect 9306 28364 9312 28416
rect 9364 28364 9370 28416
rect 9416 28404 9444 28444
rect 10137 28441 10149 28444
rect 10183 28441 10195 28475
rect 10137 28435 10195 28441
rect 10226 28432 10232 28484
rect 10284 28472 10290 28484
rect 11609 28475 11667 28481
rect 11609 28472 11621 28475
rect 10284 28444 11621 28472
rect 10284 28432 10290 28444
rect 11609 28441 11621 28444
rect 11655 28472 11667 28475
rect 12084 28472 12112 28503
rect 12342 28500 12348 28552
rect 12400 28500 12406 28552
rect 12989 28543 13047 28549
rect 12989 28509 13001 28543
rect 13035 28540 13047 28543
rect 13078 28540 13084 28552
rect 13035 28512 13084 28540
rect 13035 28509 13047 28512
rect 12989 28503 13047 28509
rect 13078 28500 13084 28512
rect 13136 28500 13142 28552
rect 13262 28500 13268 28552
rect 13320 28540 13326 28552
rect 13357 28543 13415 28549
rect 13357 28540 13369 28543
rect 13320 28512 13369 28540
rect 13320 28500 13326 28512
rect 13357 28509 13369 28512
rect 13403 28540 13415 28543
rect 13538 28540 13544 28552
rect 13403 28512 13544 28540
rect 13403 28509 13415 28512
rect 13357 28503 13415 28509
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 13722 28500 13728 28552
rect 13780 28500 13786 28552
rect 14553 28543 14611 28549
rect 14553 28540 14565 28543
rect 13832 28512 14565 28540
rect 12158 28472 12164 28484
rect 11655 28444 11836 28472
rect 12084 28444 12164 28472
rect 11655 28441 11667 28444
rect 11609 28435 11667 28441
rect 11808 28416 11836 28444
rect 12158 28432 12164 28444
rect 12216 28472 12222 28484
rect 13170 28472 13176 28484
rect 12216 28444 13176 28472
rect 12216 28432 12222 28444
rect 13170 28432 13176 28444
rect 13228 28432 13234 28484
rect 10781 28407 10839 28413
rect 10781 28404 10793 28407
rect 9416 28376 10793 28404
rect 10781 28373 10793 28376
rect 10827 28404 10839 28407
rect 10870 28404 10876 28416
rect 10827 28376 10876 28404
rect 10827 28373 10839 28376
rect 10781 28367 10839 28373
rect 10870 28364 10876 28376
rect 10928 28364 10934 28416
rect 10962 28364 10968 28416
rect 11020 28364 11026 28416
rect 11698 28364 11704 28416
rect 11756 28364 11762 28416
rect 11790 28364 11796 28416
rect 11848 28404 11854 28416
rect 13832 28404 13860 28512
rect 14553 28509 14565 28512
rect 14599 28509 14611 28543
rect 14553 28503 14611 28509
rect 14182 28432 14188 28484
rect 14240 28472 14246 28484
rect 14277 28475 14335 28481
rect 14277 28472 14289 28475
rect 14240 28444 14289 28472
rect 14240 28432 14246 28444
rect 14277 28441 14289 28444
rect 14323 28441 14335 28475
rect 14277 28435 14335 28441
rect 14461 28475 14519 28481
rect 14461 28441 14473 28475
rect 14507 28472 14519 28475
rect 14660 28472 14688 28580
rect 14829 28543 14887 28549
rect 14829 28509 14841 28543
rect 14875 28540 14887 28543
rect 15010 28540 15016 28552
rect 14875 28512 15016 28540
rect 14875 28509 14887 28512
rect 14829 28503 14887 28509
rect 15010 28500 15016 28512
rect 15068 28500 15074 28552
rect 15212 28549 15240 28580
rect 16224 28580 16764 28608
rect 15197 28543 15255 28549
rect 15197 28509 15209 28543
rect 15243 28509 15255 28543
rect 15197 28503 15255 28509
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28540 15347 28543
rect 15378 28540 15384 28552
rect 15335 28512 15384 28540
rect 15335 28509 15347 28512
rect 15289 28503 15347 28509
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 15562 28500 15568 28552
rect 15620 28500 15626 28552
rect 15654 28500 15660 28552
rect 15712 28540 15718 28552
rect 15933 28543 15991 28549
rect 15933 28540 15945 28543
rect 15712 28512 15945 28540
rect 15712 28500 15718 28512
rect 15933 28509 15945 28512
rect 15979 28509 15991 28543
rect 15933 28503 15991 28509
rect 16022 28500 16028 28552
rect 16080 28500 16086 28552
rect 16224 28549 16252 28580
rect 16758 28568 16764 28580
rect 16816 28568 16822 28620
rect 16209 28543 16267 28549
rect 16209 28509 16221 28543
rect 16255 28509 16267 28543
rect 16209 28503 16267 28509
rect 16301 28543 16359 28549
rect 16301 28509 16313 28543
rect 16347 28509 16359 28543
rect 16301 28503 16359 28509
rect 14507 28444 14688 28472
rect 14921 28475 14979 28481
rect 14507 28441 14519 28444
rect 14461 28435 14519 28441
rect 14921 28441 14933 28475
rect 14967 28472 14979 28475
rect 15473 28475 15531 28481
rect 15473 28472 15485 28475
rect 14967 28444 15485 28472
rect 14967 28441 14979 28444
rect 14921 28435 14979 28441
rect 15473 28441 15485 28444
rect 15519 28441 15531 28475
rect 16316 28472 16344 28503
rect 16390 28500 16396 28552
rect 16448 28500 16454 28552
rect 16574 28500 16580 28552
rect 16632 28500 16638 28552
rect 16666 28500 16672 28552
rect 16724 28540 16730 28552
rect 18524 28540 18552 28648
rect 18598 28568 18604 28620
rect 18656 28608 18662 28620
rect 20165 28611 20223 28617
rect 18656 28580 19012 28608
rect 18656 28568 18662 28580
rect 18984 28552 19012 28580
rect 20165 28577 20177 28611
rect 20211 28608 20223 28611
rect 20714 28608 20720 28620
rect 20211 28580 20720 28608
rect 20211 28577 20223 28580
rect 20165 28571 20223 28577
rect 20714 28568 20720 28580
rect 20772 28568 20778 28620
rect 21008 28608 21036 28648
rect 21683 28645 21695 28679
rect 21729 28676 21741 28679
rect 22373 28679 22431 28685
rect 22373 28676 22385 28679
rect 21729 28648 22385 28676
rect 21729 28645 21741 28648
rect 21683 28639 21741 28645
rect 22373 28645 22385 28648
rect 22419 28676 22431 28679
rect 22554 28676 22560 28688
rect 22419 28648 22560 28676
rect 22419 28645 22431 28648
rect 22373 28639 22431 28645
rect 22554 28636 22560 28648
rect 22612 28676 22618 28688
rect 22830 28676 22836 28688
rect 22612 28648 22836 28676
rect 22612 28636 22618 28648
rect 22830 28636 22836 28648
rect 22888 28636 22894 28688
rect 22462 28608 22468 28620
rect 21008 28580 21588 28608
rect 16724 28512 18552 28540
rect 16724 28500 16730 28512
rect 18782 28500 18788 28552
rect 18840 28500 18846 28552
rect 18966 28500 18972 28552
rect 19024 28500 19030 28552
rect 20254 28500 20260 28552
rect 20312 28540 20318 28552
rect 20530 28540 20536 28552
rect 20312 28512 20536 28540
rect 20312 28500 20318 28512
rect 20530 28500 20536 28512
rect 20588 28500 20594 28552
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28540 20959 28543
rect 20990 28540 20996 28552
rect 20947 28512 20996 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 20990 28500 20996 28512
rect 21048 28500 21054 28552
rect 21082 28500 21088 28552
rect 21140 28500 21146 28552
rect 21358 28500 21364 28552
rect 21416 28500 21422 28552
rect 17126 28472 17132 28484
rect 16316 28444 17132 28472
rect 15473 28435 15531 28441
rect 11848 28376 13860 28404
rect 11848 28364 11854 28376
rect 13906 28364 13912 28416
rect 13964 28404 13970 28416
rect 14476 28404 14504 28435
rect 17126 28432 17132 28444
rect 17184 28472 17190 28484
rect 17402 28472 17408 28484
rect 17184 28444 17408 28472
rect 17184 28432 17190 28444
rect 17402 28432 17408 28444
rect 17460 28432 17466 28484
rect 20162 28432 20168 28484
rect 20220 28472 20226 28484
rect 20441 28475 20499 28481
rect 20441 28472 20453 28475
rect 20220 28444 20453 28472
rect 20220 28432 20226 28444
rect 20441 28441 20453 28444
rect 20487 28441 20499 28475
rect 20441 28435 20499 28441
rect 20650 28475 20708 28481
rect 20650 28441 20662 28475
rect 20696 28472 20708 28475
rect 21560 28472 21588 28580
rect 21829 28580 22468 28608
rect 21829 28549 21857 28580
rect 22462 28568 22468 28580
rect 22520 28568 22526 28620
rect 22646 28568 22652 28620
rect 22704 28608 22710 28620
rect 23400 28617 23428 28716
rect 24394 28704 24400 28716
rect 24452 28704 24458 28756
rect 25590 28704 25596 28756
rect 25648 28744 25654 28756
rect 25869 28747 25927 28753
rect 25869 28744 25881 28747
rect 25648 28716 25881 28744
rect 25648 28704 25654 28716
rect 25869 28713 25881 28716
rect 25915 28713 25927 28747
rect 25869 28707 25927 28713
rect 26694 28704 26700 28756
rect 26752 28744 26758 28756
rect 27062 28744 27068 28756
rect 26752 28716 27068 28744
rect 26752 28704 26758 28716
rect 27062 28704 27068 28716
rect 27120 28704 27126 28756
rect 27617 28747 27675 28753
rect 27617 28713 27629 28747
rect 27663 28744 27675 28747
rect 27706 28744 27712 28756
rect 27663 28716 27712 28744
rect 27663 28713 27675 28716
rect 27617 28707 27675 28713
rect 27706 28704 27712 28716
rect 27764 28704 27770 28756
rect 28258 28704 28264 28756
rect 28316 28704 28322 28756
rect 28445 28747 28503 28753
rect 28445 28713 28457 28747
rect 28491 28744 28503 28747
rect 29546 28744 29552 28756
rect 28491 28716 29552 28744
rect 28491 28713 28503 28716
rect 28445 28707 28503 28713
rect 29546 28704 29552 28716
rect 29604 28704 29610 28756
rect 29914 28704 29920 28756
rect 29972 28744 29978 28756
rect 34149 28747 34207 28753
rect 34149 28744 34161 28747
rect 29972 28716 34161 28744
rect 29972 28704 29978 28716
rect 34149 28713 34161 28716
rect 34195 28713 34207 28747
rect 34149 28707 34207 28713
rect 34882 28704 34888 28756
rect 34940 28744 34946 28756
rect 35345 28747 35403 28753
rect 35345 28744 35357 28747
rect 34940 28716 35357 28744
rect 34940 28704 34946 28716
rect 35345 28713 35357 28716
rect 35391 28713 35403 28747
rect 35345 28707 35403 28713
rect 24578 28676 24584 28688
rect 24136 28648 24584 28676
rect 22741 28611 22799 28617
rect 22741 28608 22753 28611
rect 22704 28580 22753 28608
rect 22704 28568 22710 28580
rect 22741 28577 22753 28580
rect 22787 28577 22799 28611
rect 23385 28611 23443 28617
rect 23385 28608 23397 28611
rect 22741 28571 22799 28577
rect 22940 28580 23397 28608
rect 21821 28543 21879 28549
rect 21821 28509 21833 28543
rect 21867 28509 21879 28543
rect 21821 28503 21879 28509
rect 22005 28543 22063 28549
rect 22005 28509 22017 28543
rect 22051 28540 22063 28543
rect 22940 28540 22968 28580
rect 23385 28577 23397 28580
rect 23431 28577 23443 28611
rect 24136 28594 24164 28648
rect 24578 28636 24584 28648
rect 24636 28636 24642 28688
rect 24762 28636 24768 28688
rect 24820 28676 24826 28688
rect 25130 28676 25136 28688
rect 24820 28648 25136 28676
rect 24820 28636 24826 28648
rect 25130 28636 25136 28648
rect 25188 28636 25194 28688
rect 25774 28636 25780 28688
rect 25832 28676 25838 28688
rect 28074 28676 28080 28688
rect 25832 28648 26924 28676
rect 25832 28636 25838 28648
rect 23385 28571 23443 28577
rect 24486 28568 24492 28620
rect 24544 28608 24550 28620
rect 24544 28580 25360 28608
rect 24544 28568 24550 28580
rect 22051 28512 22968 28540
rect 22051 28509 22063 28512
rect 22005 28503 22063 28509
rect 23014 28500 23020 28552
rect 23072 28540 23078 28552
rect 23201 28543 23259 28549
rect 23201 28540 23213 28543
rect 23072 28512 23213 28540
rect 23072 28500 23078 28512
rect 23201 28509 23213 28512
rect 23247 28509 23259 28543
rect 23201 28503 23259 28509
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28509 24087 28543
rect 24029 28503 24087 28509
rect 24397 28543 24455 28549
rect 24397 28509 24409 28543
rect 24443 28540 24455 28543
rect 24854 28540 24860 28552
rect 24443 28512 24860 28540
rect 24443 28509 24455 28512
rect 24397 28503 24455 28509
rect 20696 28444 21496 28472
rect 21560 28444 21864 28472
rect 20696 28441 20708 28444
rect 20650 28435 20708 28441
rect 13964 28376 14504 28404
rect 15013 28407 15071 28413
rect 13964 28364 13970 28376
rect 15013 28373 15025 28407
rect 15059 28404 15071 28407
rect 15562 28404 15568 28416
rect 15059 28376 15568 28404
rect 15059 28373 15071 28376
rect 15013 28367 15071 28373
rect 15562 28364 15568 28376
rect 15620 28364 15626 28416
rect 16390 28364 16396 28416
rect 16448 28404 16454 28416
rect 16574 28404 16580 28416
rect 16448 28376 16580 28404
rect 16448 28364 16454 28376
rect 16574 28364 16580 28376
rect 16632 28364 16638 28416
rect 18874 28364 18880 28416
rect 18932 28364 18938 28416
rect 20806 28364 20812 28416
rect 20864 28404 20870 28416
rect 20993 28407 21051 28413
rect 20993 28404 21005 28407
rect 20864 28376 21005 28404
rect 20864 28364 20870 28376
rect 20993 28373 21005 28376
rect 21039 28373 21051 28407
rect 20993 28367 21051 28373
rect 21358 28364 21364 28416
rect 21416 28364 21422 28416
rect 21468 28404 21496 28444
rect 21726 28404 21732 28416
rect 21468 28376 21732 28404
rect 21726 28364 21732 28376
rect 21784 28364 21790 28416
rect 21836 28404 21864 28444
rect 22370 28432 22376 28484
rect 22428 28472 22434 28484
rect 23566 28472 23572 28484
rect 22428 28444 23572 28472
rect 22428 28432 22434 28444
rect 23566 28432 23572 28444
rect 23624 28472 23630 28484
rect 24044 28472 24072 28503
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 24946 28500 24952 28552
rect 25004 28500 25010 28552
rect 25038 28500 25044 28552
rect 25096 28540 25102 28552
rect 25225 28543 25283 28549
rect 25225 28540 25237 28543
rect 25096 28512 25237 28540
rect 25096 28500 25102 28512
rect 25225 28509 25237 28512
rect 25271 28509 25283 28543
rect 25332 28540 25360 28580
rect 25682 28568 25688 28620
rect 25740 28608 25746 28620
rect 26694 28608 26700 28620
rect 25740 28580 26280 28608
rect 25740 28568 25746 28580
rect 26252 28549 26280 28580
rect 26436 28580 26700 28608
rect 26436 28549 26464 28580
rect 26694 28568 26700 28580
rect 26752 28568 26758 28620
rect 26053 28543 26111 28549
rect 26053 28540 26065 28543
rect 25332 28512 26065 28540
rect 25225 28503 25283 28509
rect 26053 28509 26065 28512
rect 26099 28509 26111 28543
rect 26053 28503 26111 28509
rect 26237 28543 26295 28549
rect 26237 28509 26249 28543
rect 26283 28509 26295 28543
rect 26237 28503 26295 28509
rect 26421 28543 26479 28549
rect 26421 28509 26433 28543
rect 26467 28509 26479 28543
rect 26421 28503 26479 28509
rect 26510 28500 26516 28552
rect 26568 28500 26574 28552
rect 26602 28500 26608 28552
rect 26660 28500 26666 28552
rect 24762 28472 24768 28484
rect 23624 28444 24768 28472
rect 23624 28432 23630 28444
rect 24762 28432 24768 28444
rect 24820 28432 24826 28484
rect 22186 28404 22192 28416
rect 21836 28376 22192 28404
rect 22186 28364 22192 28376
rect 22244 28364 22250 28416
rect 22649 28407 22707 28413
rect 22649 28373 22661 28407
rect 22695 28404 22707 28407
rect 23198 28404 23204 28416
rect 22695 28376 23204 28404
rect 22695 28373 22707 28376
rect 22649 28367 22707 28373
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 23750 28364 23756 28416
rect 23808 28413 23814 28416
rect 23808 28407 23837 28413
rect 23825 28373 23837 28407
rect 23808 28367 23837 28373
rect 23808 28364 23814 28367
rect 24118 28364 24124 28416
rect 24176 28404 24182 28416
rect 24581 28407 24639 28413
rect 24581 28404 24593 28407
rect 24176 28376 24593 28404
rect 24176 28364 24182 28376
rect 24581 28373 24593 28376
rect 24627 28404 24639 28407
rect 24670 28404 24676 28416
rect 24627 28376 24676 28404
rect 24627 28373 24639 28376
rect 24581 28367 24639 28373
rect 24670 28364 24676 28376
rect 24728 28364 24734 28416
rect 24964 28404 24992 28500
rect 26145 28475 26203 28481
rect 26145 28441 26157 28475
rect 26191 28472 26203 28475
rect 26326 28472 26332 28484
rect 26191 28444 26332 28472
rect 26191 28441 26203 28444
rect 26145 28435 26203 28441
rect 26326 28432 26332 28444
rect 26384 28432 26390 28484
rect 26789 28407 26847 28413
rect 26789 28404 26801 28407
rect 24964 28376 26801 28404
rect 26789 28373 26801 28376
rect 26835 28373 26847 28407
rect 26896 28404 26924 28648
rect 27816 28648 28080 28676
rect 27522 28608 27528 28620
rect 26988 28580 27528 28608
rect 26988 28540 27016 28580
rect 27522 28568 27528 28580
rect 27580 28568 27586 28620
rect 27816 28617 27844 28648
rect 28074 28636 28080 28648
rect 28132 28636 28138 28688
rect 28626 28636 28632 28688
rect 28684 28676 28690 28688
rect 28902 28676 28908 28688
rect 28684 28648 28908 28676
rect 28684 28636 28690 28648
rect 28902 28636 28908 28648
rect 28960 28676 28966 28688
rect 28960 28648 32812 28676
rect 28960 28636 28966 28648
rect 27783 28611 27844 28617
rect 27783 28577 27795 28611
rect 27829 28580 27844 28611
rect 28537 28611 28595 28617
rect 28537 28608 28549 28611
rect 28000 28580 28549 28608
rect 27829 28577 27841 28580
rect 27783 28571 27841 28577
rect 27065 28543 27123 28549
rect 27065 28540 27077 28543
rect 26988 28512 27077 28540
rect 27065 28509 27077 28512
rect 27111 28509 27123 28543
rect 27065 28503 27123 28509
rect 27433 28543 27491 28549
rect 27433 28509 27445 28543
rect 27479 28540 27491 28543
rect 27614 28540 27620 28552
rect 27479 28512 27620 28540
rect 27479 28509 27501 28512
rect 27433 28506 27501 28509
rect 27433 28503 27491 28506
rect 27614 28500 27620 28512
rect 27672 28540 27678 28552
rect 27893 28543 27951 28549
rect 27893 28540 27905 28543
rect 27672 28534 27752 28540
rect 27872 28534 27905 28540
rect 27672 28512 27905 28534
rect 27672 28500 27678 28512
rect 27724 28509 27905 28512
rect 27939 28509 27951 28543
rect 27724 28506 27951 28509
rect 27893 28503 27951 28506
rect 27246 28432 27252 28484
rect 27304 28432 27310 28484
rect 27338 28432 27344 28484
rect 27396 28432 27402 28484
rect 28000 28404 28028 28580
rect 28537 28577 28549 28580
rect 28583 28577 28595 28611
rect 28537 28571 28595 28577
rect 28810 28568 28816 28620
rect 28868 28568 28874 28620
rect 30098 28568 30104 28620
rect 30156 28608 30162 28620
rect 32217 28611 32275 28617
rect 30156 28580 31984 28608
rect 30156 28568 30162 28580
rect 28258 28500 28264 28552
rect 28316 28540 28322 28552
rect 28718 28540 28724 28552
rect 28316 28512 28724 28540
rect 28316 28500 28322 28512
rect 28718 28500 28724 28512
rect 28776 28500 28782 28552
rect 29914 28540 29920 28552
rect 29748 28512 29920 28540
rect 28626 28432 28632 28484
rect 28684 28472 28690 28484
rect 29546 28472 29552 28484
rect 28684 28444 29552 28472
rect 28684 28432 28690 28444
rect 29546 28432 29552 28444
rect 29604 28472 29610 28484
rect 29748 28472 29776 28512
rect 29914 28500 29920 28512
rect 29972 28500 29978 28552
rect 30190 28500 30196 28552
rect 30248 28540 30254 28552
rect 31757 28543 31815 28549
rect 31757 28540 31769 28543
rect 30248 28512 31769 28540
rect 30248 28500 30254 28512
rect 31757 28509 31769 28512
rect 31803 28509 31815 28543
rect 31757 28503 31815 28509
rect 29604 28444 29776 28472
rect 29604 28432 29610 28444
rect 29822 28432 29828 28484
rect 29880 28472 29886 28484
rect 29880 28444 31800 28472
rect 29880 28432 29886 28444
rect 26896 28376 28028 28404
rect 26789 28367 26847 28373
rect 28442 28364 28448 28416
rect 28500 28404 28506 28416
rect 30834 28404 30840 28416
rect 28500 28376 30840 28404
rect 28500 28364 28506 28376
rect 30834 28364 30840 28376
rect 30892 28364 30898 28416
rect 31573 28407 31631 28413
rect 31573 28373 31585 28407
rect 31619 28404 31631 28407
rect 31662 28404 31668 28416
rect 31619 28376 31668 28404
rect 31619 28373 31631 28376
rect 31573 28367 31631 28373
rect 31662 28364 31668 28376
rect 31720 28364 31726 28416
rect 31772 28404 31800 28444
rect 31846 28432 31852 28484
rect 31904 28432 31910 28484
rect 31956 28481 31984 28580
rect 32217 28577 32229 28611
rect 32263 28608 32275 28611
rect 32674 28608 32680 28620
rect 32263 28580 32680 28608
rect 32263 28577 32275 28580
rect 32217 28571 32275 28577
rect 32674 28568 32680 28580
rect 32732 28568 32738 28620
rect 32784 28608 32812 28648
rect 33318 28636 33324 28688
rect 33376 28676 33382 28688
rect 34333 28679 34391 28685
rect 34333 28676 34345 28679
rect 33376 28648 34345 28676
rect 33376 28636 33382 28648
rect 34333 28645 34345 28648
rect 34379 28645 34391 28679
rect 34333 28639 34391 28645
rect 34422 28636 34428 28688
rect 34480 28676 34486 28688
rect 34480 28648 35204 28676
rect 34480 28636 34486 28648
rect 34701 28611 34759 28617
rect 34701 28608 34713 28611
rect 32784 28580 34713 28608
rect 34701 28577 34713 28580
rect 34747 28577 34759 28611
rect 34701 28571 34759 28577
rect 34790 28568 34796 28620
rect 34848 28608 34854 28620
rect 34848 28580 35112 28608
rect 34848 28568 34854 28580
rect 32030 28500 32036 28552
rect 32088 28549 32094 28552
rect 32088 28543 32117 28549
rect 32105 28509 32117 28543
rect 32088 28503 32117 28509
rect 32088 28500 32094 28503
rect 33778 28500 33784 28552
rect 33836 28500 33842 28552
rect 34808 28540 34836 28568
rect 35084 28549 35112 28580
rect 35176 28549 35204 28648
rect 33888 28512 34836 28540
rect 35069 28543 35127 28549
rect 31941 28475 31999 28481
rect 31941 28441 31953 28475
rect 31987 28472 31999 28475
rect 33888 28472 33916 28512
rect 35069 28509 35081 28543
rect 35115 28509 35127 28543
rect 35069 28503 35127 28509
rect 35161 28543 35219 28549
rect 35161 28509 35173 28543
rect 35207 28509 35219 28543
rect 35161 28503 35219 28509
rect 31987 28444 33916 28472
rect 31987 28441 31999 28444
rect 31941 28435 31999 28441
rect 34698 28432 34704 28484
rect 34756 28472 34762 28484
rect 34839 28475 34897 28481
rect 34839 28472 34851 28475
rect 34756 28444 34851 28472
rect 34756 28432 34762 28444
rect 34839 28441 34851 28444
rect 34885 28441 34897 28475
rect 34839 28435 34897 28441
rect 34977 28475 35035 28481
rect 34977 28441 34989 28475
rect 35023 28472 35035 28475
rect 35618 28472 35624 28484
rect 35023 28444 35624 28472
rect 35023 28441 35035 28444
rect 34977 28435 35035 28441
rect 34158 28407 34216 28413
rect 34158 28404 34170 28407
rect 31772 28376 34170 28404
rect 34158 28373 34170 28376
rect 34204 28373 34216 28407
rect 34158 28367 34216 28373
rect 34606 28364 34612 28416
rect 34664 28404 34670 28416
rect 34992 28404 35020 28435
rect 35618 28432 35624 28444
rect 35676 28432 35682 28484
rect 34664 28376 35020 28404
rect 34664 28364 34670 28376
rect 1104 28314 36432 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 36432 28314
rect 1104 28240 36432 28262
rect 2774 28200 2780 28212
rect 2746 28160 2780 28200
rect 2832 28160 2838 28212
rect 3510 28160 3516 28212
rect 3568 28200 3574 28212
rect 4341 28203 4399 28209
rect 4341 28200 4353 28203
rect 3568 28172 4353 28200
rect 3568 28160 3574 28172
rect 4341 28169 4353 28172
rect 4387 28200 4399 28203
rect 5718 28200 5724 28212
rect 4387 28172 5724 28200
rect 4387 28169 4399 28172
rect 4341 28163 4399 28169
rect 5718 28160 5724 28172
rect 5776 28160 5782 28212
rect 7190 28160 7196 28212
rect 7248 28200 7254 28212
rect 7377 28203 7435 28209
rect 7377 28200 7389 28203
rect 7248 28172 7389 28200
rect 7248 28160 7254 28172
rect 7377 28169 7389 28172
rect 7423 28169 7435 28203
rect 7377 28163 7435 28169
rect 9217 28203 9275 28209
rect 9217 28169 9229 28203
rect 9263 28200 9275 28203
rect 9674 28200 9680 28212
rect 9263 28172 9680 28200
rect 9263 28169 9275 28172
rect 9217 28163 9275 28169
rect 2746 28132 2774 28160
rect 5994 28132 6000 28144
rect 2714 28104 2774 28132
rect 4724 28104 6000 28132
rect 3418 28024 3424 28076
rect 3476 28064 3482 28076
rect 3602 28064 3608 28076
rect 3476 28036 3608 28064
rect 3476 28024 3482 28036
rect 3602 28024 3608 28036
rect 3660 28024 3666 28076
rect 4338 28067 4396 28073
rect 4338 28033 4350 28067
rect 4384 28064 4396 28067
rect 4724 28064 4752 28104
rect 5994 28092 6000 28104
rect 6052 28092 6058 28144
rect 6914 28092 6920 28144
rect 6972 28092 6978 28144
rect 7006 28092 7012 28144
rect 7064 28132 7070 28144
rect 7101 28135 7159 28141
rect 7101 28132 7113 28135
rect 7064 28104 7113 28132
rect 7064 28092 7070 28104
rect 7101 28101 7113 28104
rect 7147 28132 7159 28135
rect 7469 28135 7527 28141
rect 7469 28132 7481 28135
rect 7147 28104 7481 28132
rect 7147 28101 7159 28104
rect 7101 28095 7159 28101
rect 7469 28101 7481 28104
rect 7515 28101 7527 28135
rect 7742 28132 7748 28144
rect 7469 28095 7527 28101
rect 7576 28104 7748 28132
rect 4384 28036 4752 28064
rect 4801 28067 4859 28073
rect 4384 28033 4396 28036
rect 4338 28027 4396 28033
rect 4801 28033 4813 28067
rect 4847 28064 4859 28067
rect 5258 28064 5264 28076
rect 4847 28036 5264 28064
rect 4847 28033 4859 28036
rect 4801 28027 4859 28033
rect 5258 28024 5264 28036
rect 5316 28024 5322 28076
rect 5813 28067 5871 28073
rect 5813 28033 5825 28067
rect 5859 28064 5871 28067
rect 5902 28064 5908 28076
rect 5859 28036 5908 28064
rect 5859 28033 5871 28036
rect 5813 28027 5871 28033
rect 5902 28024 5908 28036
rect 5960 28024 5966 28076
rect 6089 28067 6147 28073
rect 6089 28033 6101 28067
rect 6135 28064 6147 28067
rect 6730 28064 6736 28076
rect 6135 28036 6736 28064
rect 6135 28033 6147 28036
rect 6089 28027 6147 28033
rect 6730 28024 6736 28036
rect 6788 28064 6794 28076
rect 7377 28067 7435 28073
rect 6788 28036 7328 28064
rect 6788 28024 6794 28036
rect 1394 27956 1400 28008
rect 1452 27956 1458 28008
rect 3142 27956 3148 28008
rect 3200 27956 3206 28008
rect 4982 28005 4988 28008
rect 4709 27999 4767 28005
rect 4709 27965 4721 27999
rect 4755 27996 4767 27999
rect 4939 27999 4988 28005
rect 4755 27968 4844 27996
rect 4755 27965 4767 27968
rect 4709 27959 4767 27965
rect 4816 27928 4844 27968
rect 4939 27965 4951 27999
rect 4985 27965 4988 27999
rect 4939 27959 4988 27965
rect 4982 27956 4988 27959
rect 5040 27956 5046 28008
rect 7190 27956 7196 28008
rect 7248 27956 7254 28008
rect 7300 27996 7328 28036
rect 7377 28033 7389 28067
rect 7423 28064 7435 28067
rect 7576 28064 7604 28104
rect 7742 28092 7748 28104
rect 7800 28092 7806 28144
rect 9232 28132 9260 28163
rect 9674 28160 9680 28172
rect 9732 28160 9738 28212
rect 9766 28160 9772 28212
rect 9824 28200 9830 28212
rect 10410 28200 10416 28212
rect 9824 28172 10416 28200
rect 9824 28160 9830 28172
rect 10410 28160 10416 28172
rect 10468 28160 10474 28212
rect 13170 28160 13176 28212
rect 13228 28160 13234 28212
rect 15378 28160 15384 28212
rect 15436 28200 15442 28212
rect 17862 28200 17868 28212
rect 15436 28172 17868 28200
rect 15436 28160 15442 28172
rect 17862 28160 17868 28172
rect 17920 28160 17926 28212
rect 19150 28200 19156 28212
rect 18984 28172 19156 28200
rect 8772 28104 9260 28132
rect 7423 28036 7604 28064
rect 7653 28067 7711 28073
rect 7423 28033 7435 28036
rect 7377 28027 7435 28033
rect 7653 28033 7665 28067
rect 7699 28064 7711 28067
rect 8110 28064 8116 28076
rect 7699 28036 8116 28064
rect 7699 28033 7711 28036
rect 7653 28027 7711 28033
rect 8110 28024 8116 28036
rect 8168 28024 8174 28076
rect 8772 28073 8800 28104
rect 9306 28092 9312 28144
rect 9364 28132 9370 28144
rect 10962 28132 10968 28144
rect 9364 28104 10088 28132
rect 9364 28092 9370 28104
rect 8296 28067 8354 28073
rect 8296 28033 8308 28067
rect 8342 28064 8354 28067
rect 8573 28067 8631 28073
rect 8573 28064 8585 28067
rect 8342 28036 8585 28064
rect 8342 28033 8354 28036
rect 8296 28027 8354 28033
rect 8573 28033 8585 28036
rect 8619 28033 8631 28067
rect 8573 28027 8631 28033
rect 8757 28067 8815 28073
rect 8757 28033 8769 28067
rect 8803 28033 8815 28067
rect 8757 28027 8815 28033
rect 8846 28024 8852 28076
rect 8904 28024 8910 28076
rect 9030 28024 9036 28076
rect 9088 28064 9094 28076
rect 9125 28067 9183 28073
rect 9125 28064 9137 28067
rect 9088 28036 9137 28064
rect 9088 28024 9094 28036
rect 9125 28033 9137 28036
rect 9171 28033 9183 28067
rect 9125 28027 9183 28033
rect 9214 28024 9220 28076
rect 9272 28024 9278 28076
rect 9401 28067 9459 28073
rect 9401 28033 9413 28067
rect 9447 28064 9459 28067
rect 9582 28064 9588 28076
rect 9447 28036 9588 28064
rect 9447 28033 9459 28036
rect 9401 28027 9459 28033
rect 9582 28024 9588 28036
rect 9640 28024 9646 28076
rect 9766 28024 9772 28076
rect 9824 28024 9830 28076
rect 10060 28073 10088 28104
rect 10152 28104 10968 28132
rect 10152 28073 10180 28104
rect 10962 28092 10968 28104
rect 11020 28092 11026 28144
rect 11698 28092 11704 28144
rect 11756 28132 11762 28144
rect 11756 28104 12480 28132
rect 11756 28092 11762 28104
rect 9953 28067 10011 28073
rect 9953 28033 9965 28067
rect 9999 28033 10011 28067
rect 9953 28027 10011 28033
rect 10045 28067 10103 28073
rect 10045 28033 10057 28067
rect 10091 28033 10103 28067
rect 10045 28027 10103 28033
rect 10137 28067 10195 28073
rect 10137 28033 10149 28067
rect 10183 28033 10195 28067
rect 10137 28027 10195 28033
rect 7837 27999 7895 28005
rect 7837 27996 7849 27999
rect 7300 27968 7849 27996
rect 7837 27965 7849 27968
rect 7883 27965 7895 27999
rect 7837 27959 7895 27965
rect 7929 27999 7987 28005
rect 7929 27965 7941 27999
rect 7975 27996 7987 27999
rect 8018 27996 8024 28008
rect 7975 27968 8024 27996
rect 7975 27965 7987 27968
rect 7929 27959 7987 27965
rect 5258 27928 5264 27940
rect 4080 27900 4752 27928
rect 4816 27900 5264 27928
rect 2498 27820 2504 27872
rect 2556 27860 2562 27872
rect 4080 27860 4108 27900
rect 2556 27832 4108 27860
rect 4157 27863 4215 27869
rect 2556 27820 2562 27832
rect 4157 27829 4169 27863
rect 4203 27860 4215 27863
rect 4614 27860 4620 27872
rect 4203 27832 4620 27860
rect 4203 27829 4215 27832
rect 4157 27823 4215 27829
rect 4614 27820 4620 27832
rect 4672 27820 4678 27872
rect 4724 27860 4752 27900
rect 5258 27888 5264 27900
rect 5316 27888 5322 27940
rect 5353 27931 5411 27937
rect 5353 27897 5365 27931
rect 5399 27928 5411 27931
rect 7852 27928 7880 27959
rect 8018 27956 8024 27968
rect 8076 27956 8082 28008
rect 8481 27999 8539 28005
rect 8481 27965 8493 27999
rect 8527 27996 8539 27999
rect 9674 27996 9680 28008
rect 8527 27968 9680 27996
rect 8527 27965 8539 27968
rect 8481 27959 8539 27965
rect 9674 27956 9680 27968
rect 9732 27956 9738 28008
rect 9784 27928 9812 28024
rect 9968 27996 9996 28027
rect 10226 28024 10232 28076
rect 10284 28024 10290 28076
rect 10318 28024 10324 28076
rect 10376 28064 10382 28076
rect 10505 28067 10563 28073
rect 10505 28064 10517 28067
rect 10376 28036 10517 28064
rect 10376 28024 10382 28036
rect 10505 28033 10517 28036
rect 10551 28033 10563 28067
rect 10505 28027 10563 28033
rect 10594 28024 10600 28076
rect 10652 28024 10658 28076
rect 10778 28024 10784 28076
rect 10836 28064 10842 28076
rect 11057 28067 11115 28073
rect 11057 28064 11069 28067
rect 10836 28036 11069 28064
rect 10836 28024 10842 28036
rect 11057 28033 11069 28036
rect 11103 28033 11115 28067
rect 11057 28027 11115 28033
rect 11238 28024 11244 28076
rect 11296 28024 11302 28076
rect 11885 28067 11943 28073
rect 11885 28033 11897 28067
rect 11931 28064 11943 28067
rect 12250 28064 12256 28076
rect 11931 28036 12256 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 12250 28024 12256 28036
rect 12308 28024 12314 28076
rect 12342 28024 12348 28076
rect 12400 28024 12406 28076
rect 12452 28073 12480 28104
rect 13078 28092 13084 28144
rect 13136 28132 13142 28144
rect 13136 28104 13584 28132
rect 13136 28092 13142 28104
rect 13556 28076 13584 28104
rect 18230 28092 18236 28144
rect 18288 28132 18294 28144
rect 18984 28132 19012 28172
rect 19150 28160 19156 28172
rect 19208 28160 19214 28212
rect 19242 28160 19248 28212
rect 19300 28200 19306 28212
rect 20993 28203 21051 28209
rect 19300 28160 19334 28200
rect 20993 28169 21005 28203
rect 21039 28200 21051 28203
rect 21818 28200 21824 28212
rect 21039 28172 21824 28200
rect 21039 28169 21051 28172
rect 20993 28163 21051 28169
rect 21818 28160 21824 28172
rect 21876 28160 21882 28212
rect 24578 28160 24584 28212
rect 24636 28200 24642 28212
rect 24636 28172 25084 28200
rect 24636 28160 24642 28172
rect 18288 28104 19012 28132
rect 19306 28132 19334 28160
rect 25056 28144 25084 28172
rect 25130 28160 25136 28212
rect 25188 28200 25194 28212
rect 25501 28203 25559 28209
rect 25501 28200 25513 28203
rect 25188 28172 25513 28200
rect 25188 28160 25194 28172
rect 25501 28169 25513 28172
rect 25547 28169 25559 28203
rect 25501 28163 25559 28169
rect 25961 28203 26019 28209
rect 25961 28169 25973 28203
rect 26007 28200 26019 28203
rect 26510 28200 26516 28212
rect 26007 28172 26516 28200
rect 26007 28169 26019 28172
rect 25961 28163 26019 28169
rect 26510 28160 26516 28172
rect 26568 28160 26574 28212
rect 27157 28203 27215 28209
rect 27157 28200 27169 28203
rect 26620 28172 27169 28200
rect 19306 28104 20760 28132
rect 18288 28092 18294 28104
rect 12437 28067 12495 28073
rect 12437 28033 12449 28067
rect 12483 28033 12495 28067
rect 12437 28027 12495 28033
rect 13357 28067 13415 28073
rect 13357 28033 13369 28067
rect 13403 28033 13415 28067
rect 13357 28027 13415 28033
rect 10612 27996 10640 28024
rect 9968 27968 10640 27996
rect 10965 27999 11023 28005
rect 10060 27940 10088 27968
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11149 27999 11207 28005
rect 11011 27968 11100 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 11072 27940 11100 27968
rect 11149 27965 11161 27999
rect 11195 27996 11207 27999
rect 12069 27999 12127 28005
rect 12069 27996 12081 27999
rect 11195 27968 12081 27996
rect 11195 27965 11207 27968
rect 11149 27959 11207 27965
rect 12069 27965 12081 27968
rect 12115 27965 12127 27999
rect 13372 27996 13400 28027
rect 13538 28024 13544 28076
rect 13596 28024 13602 28076
rect 14093 28067 14151 28073
rect 14093 28033 14105 28067
rect 14139 28064 14151 28067
rect 14458 28064 14464 28076
rect 14139 28036 14464 28064
rect 14139 28033 14151 28036
rect 14093 28027 14151 28033
rect 14458 28024 14464 28036
rect 14516 28024 14522 28076
rect 14737 28067 14795 28073
rect 14737 28033 14749 28067
rect 14783 28064 14795 28067
rect 14826 28064 14832 28076
rect 14783 28036 14832 28064
rect 14783 28033 14795 28036
rect 14737 28027 14795 28033
rect 14826 28024 14832 28036
rect 14884 28024 14890 28076
rect 15470 28024 15476 28076
rect 15528 28024 15534 28076
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16298 28064 16304 28076
rect 16163 28036 16304 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 16298 28024 16304 28036
rect 16356 28024 16362 28076
rect 16666 28024 16672 28076
rect 16724 28064 16730 28076
rect 16942 28064 16948 28076
rect 16724 28036 16948 28064
rect 16724 28024 16730 28036
rect 16942 28024 16948 28036
rect 17000 28064 17006 28076
rect 17129 28067 17187 28073
rect 17129 28064 17141 28067
rect 17000 28036 17141 28064
rect 17000 28024 17006 28036
rect 17129 28033 17141 28036
rect 17175 28033 17187 28067
rect 17129 28027 17187 28033
rect 17310 28024 17316 28076
rect 17368 28024 17374 28076
rect 17494 28024 17500 28076
rect 17552 28064 17558 28076
rect 17678 28064 17684 28076
rect 17552 28036 17684 28064
rect 17552 28024 17558 28036
rect 17678 28024 17684 28036
rect 17736 28064 17742 28076
rect 18984 28073 19012 28104
rect 18509 28067 18567 28073
rect 18509 28064 18521 28067
rect 17736 28036 18521 28064
rect 17736 28024 17742 28036
rect 18509 28033 18521 28036
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 18785 28067 18843 28073
rect 18785 28033 18797 28067
rect 18831 28064 18843 28067
rect 18969 28067 19027 28073
rect 18831 28036 18920 28064
rect 18831 28033 18843 28036
rect 18785 28027 18843 28033
rect 13446 27996 13452 28008
rect 13372 27968 13452 27996
rect 12069 27959 12127 27965
rect 13446 27956 13452 27968
rect 13504 27996 13510 28008
rect 13722 27996 13728 28008
rect 13504 27968 13728 27996
rect 13504 27956 13510 27968
rect 13722 27956 13728 27968
rect 13780 27996 13786 28008
rect 14921 27999 14979 28005
rect 14921 27996 14933 27999
rect 13780 27968 14933 27996
rect 13780 27956 13786 27968
rect 14921 27965 14933 27968
rect 14967 27965 14979 27999
rect 14921 27959 14979 27965
rect 15654 27956 15660 28008
rect 15712 27996 15718 28008
rect 16482 27996 16488 28008
rect 15712 27968 16488 27996
rect 15712 27956 15718 27968
rect 16482 27956 16488 27968
rect 16540 27996 16546 28008
rect 16761 27999 16819 28005
rect 16761 27996 16773 27999
rect 16540 27968 16773 27996
rect 16540 27956 16546 27968
rect 16761 27965 16773 27968
rect 16807 27965 16819 27999
rect 18892 27996 18920 28036
rect 18969 28033 18981 28067
rect 19015 28033 19027 28067
rect 18969 28027 19027 28033
rect 19150 28024 19156 28076
rect 19208 28054 19214 28076
rect 20732 28073 20760 28104
rect 20898 28092 20904 28144
rect 20956 28132 20962 28144
rect 21174 28132 21180 28144
rect 20956 28104 21180 28132
rect 20956 28092 20962 28104
rect 21174 28092 21180 28104
rect 21232 28092 21238 28144
rect 22186 28092 22192 28144
rect 22244 28132 22250 28144
rect 23750 28132 23756 28144
rect 22244 28104 23756 28132
rect 22244 28092 22250 28104
rect 23750 28092 23756 28104
rect 23808 28092 23814 28144
rect 25038 28092 25044 28144
rect 25096 28132 25102 28144
rect 25593 28135 25651 28141
rect 25593 28132 25605 28135
rect 25096 28104 25605 28132
rect 25096 28092 25102 28104
rect 25593 28101 25605 28104
rect 25639 28101 25651 28135
rect 25593 28095 25651 28101
rect 26418 28092 26424 28144
rect 26476 28092 26482 28144
rect 26620 28132 26648 28172
rect 27157 28169 27169 28172
rect 27203 28169 27215 28203
rect 27157 28163 27215 28169
rect 27338 28160 27344 28212
rect 27396 28200 27402 28212
rect 27522 28200 27528 28212
rect 27396 28172 27528 28200
rect 27396 28160 27402 28172
rect 27522 28160 27528 28172
rect 27580 28160 27586 28212
rect 27614 28160 27620 28212
rect 27672 28160 27678 28212
rect 27706 28160 27712 28212
rect 27764 28200 27770 28212
rect 28813 28203 28871 28209
rect 28813 28200 28825 28203
rect 27764 28172 28825 28200
rect 27764 28160 27770 28172
rect 28813 28169 28825 28172
rect 28859 28169 28871 28203
rect 36354 28200 36360 28212
rect 28813 28163 28871 28169
rect 30668 28172 36360 28200
rect 26528 28104 26648 28132
rect 19705 28067 19763 28073
rect 19705 28064 19717 28067
rect 19260 28054 19717 28064
rect 19208 28036 19717 28054
rect 19208 28026 19288 28036
rect 19705 28033 19717 28036
rect 19751 28033 19763 28067
rect 19705 28027 19763 28033
rect 20717 28067 20775 28073
rect 20717 28033 20729 28067
rect 20763 28033 20775 28067
rect 20717 28027 20775 28033
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22281 28067 22339 28073
rect 22281 28033 22293 28067
rect 22327 28064 22339 28067
rect 22327 28033 22340 28064
rect 22281 28027 22340 28033
rect 19208 28024 19214 28026
rect 19061 27999 19119 28005
rect 19061 27996 19073 27999
rect 18892 27968 19073 27996
rect 16761 27959 16819 27965
rect 19061 27965 19073 27968
rect 19107 27996 19119 27999
rect 19426 27996 19432 28008
rect 19107 27968 19432 27996
rect 19107 27965 19119 27968
rect 19061 27959 19119 27965
rect 19426 27956 19432 27968
rect 19484 27956 19490 28008
rect 19518 27956 19524 28008
rect 19576 27956 19582 28008
rect 21910 27956 21916 28008
rect 21968 27996 21974 28008
rect 22020 27996 22048 28027
rect 21968 27968 22048 27996
rect 21968 27956 21974 27968
rect 5399 27900 7144 27928
rect 7852 27900 9812 27928
rect 5399 27897 5411 27900
rect 5353 27891 5411 27897
rect 6641 27863 6699 27869
rect 6641 27860 6653 27863
rect 4724 27832 6653 27860
rect 6641 27829 6653 27832
rect 6687 27829 6699 27863
rect 7116 27860 7144 27900
rect 10042 27888 10048 27940
rect 10100 27888 10106 27940
rect 11054 27888 11060 27940
rect 11112 27888 11118 27940
rect 11514 27888 11520 27940
rect 11572 27888 11578 27940
rect 18966 27888 18972 27940
rect 19024 27928 19030 27940
rect 19153 27931 19211 27937
rect 19153 27928 19165 27931
rect 19024 27900 19165 27928
rect 19024 27888 19030 27900
rect 19153 27897 19165 27900
rect 19199 27897 19211 27931
rect 19153 27891 19211 27897
rect 19610 27888 19616 27940
rect 19668 27928 19674 27940
rect 19889 27931 19947 27937
rect 19889 27928 19901 27931
rect 19668 27900 19901 27928
rect 19668 27888 19674 27900
rect 19889 27897 19901 27900
rect 19935 27928 19947 27931
rect 19978 27928 19984 27940
rect 19935 27900 19984 27928
rect 19935 27897 19947 27900
rect 19889 27891 19947 27897
rect 19978 27888 19984 27900
rect 20036 27888 20042 27940
rect 22312 27928 22340 28027
rect 22370 28024 22376 28076
rect 22428 28024 22434 28076
rect 22922 28024 22928 28076
rect 22980 28024 22986 28076
rect 23106 28024 23112 28076
rect 23164 28024 23170 28076
rect 23382 28024 23388 28076
rect 23440 28024 23446 28076
rect 24762 28024 24768 28076
rect 24820 28024 24826 28076
rect 26234 28024 26240 28076
rect 26292 28064 26298 28076
rect 26528 28064 26556 28104
rect 26878 28092 26884 28144
rect 26936 28132 26942 28144
rect 26973 28135 27031 28141
rect 26973 28132 26985 28135
rect 26936 28104 26985 28132
rect 26936 28092 26942 28104
rect 26973 28101 26985 28104
rect 27019 28101 27031 28135
rect 26973 28095 27031 28101
rect 28258 28092 28264 28144
rect 28316 28132 28322 28144
rect 29779 28135 29837 28141
rect 29779 28132 29791 28135
rect 28316 28104 29791 28132
rect 28316 28092 28322 28104
rect 29779 28101 29791 28104
rect 29825 28101 29837 28135
rect 29779 28095 29837 28101
rect 30006 28092 30012 28144
rect 30064 28132 30070 28144
rect 30668 28132 30696 28172
rect 36354 28160 36360 28172
rect 36412 28160 36418 28212
rect 30064 28104 30696 28132
rect 30064 28092 30070 28104
rect 26292 28036 26556 28064
rect 26292 28024 26298 28036
rect 27062 28024 27068 28076
rect 27120 28064 27126 28076
rect 27525 28067 27583 28073
rect 27525 28064 27537 28067
rect 27120 28036 27537 28064
rect 27120 28024 27126 28036
rect 27525 28033 27537 28036
rect 27571 28033 27583 28067
rect 27525 28027 27583 28033
rect 27709 28067 27767 28073
rect 27709 28033 27721 28067
rect 27755 28064 27767 28067
rect 27755 28036 27844 28064
rect 27755 28033 27767 28036
rect 27709 28027 27767 28033
rect 22830 27956 22836 28008
rect 22888 27956 22894 28008
rect 23017 27999 23075 28005
rect 23017 27965 23029 27999
rect 23063 27965 23075 27999
rect 23017 27959 23075 27965
rect 22922 27928 22928 27940
rect 22312 27900 22928 27928
rect 22922 27888 22928 27900
rect 22980 27888 22986 27940
rect 7834 27860 7840 27872
rect 7116 27832 7840 27860
rect 6641 27823 6699 27829
rect 7834 27820 7840 27832
rect 7892 27820 7898 27872
rect 8110 27820 8116 27872
rect 8168 27860 8174 27872
rect 9033 27863 9091 27869
rect 9033 27860 9045 27863
rect 8168 27832 9045 27860
rect 8168 27820 8174 27832
rect 9033 27829 9045 27832
rect 9079 27860 9091 27863
rect 9582 27860 9588 27872
rect 9079 27832 9588 27860
rect 9079 27829 9091 27832
rect 9033 27823 9091 27829
rect 9582 27820 9588 27832
rect 9640 27820 9646 27872
rect 9674 27820 9680 27872
rect 9732 27860 9738 27872
rect 9769 27863 9827 27869
rect 9769 27860 9781 27863
rect 9732 27832 9781 27860
rect 9732 27820 9738 27832
rect 9769 27829 9781 27832
rect 9815 27829 9827 27863
rect 9769 27823 9827 27829
rect 10778 27820 10784 27872
rect 10836 27820 10842 27872
rect 11606 27820 11612 27872
rect 11664 27860 11670 27872
rect 12894 27860 12900 27872
rect 11664 27832 12900 27860
rect 11664 27820 11670 27832
rect 12894 27820 12900 27832
rect 12952 27820 12958 27872
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 18325 27863 18383 27869
rect 18325 27860 18337 27863
rect 18012 27832 18337 27860
rect 18012 27820 18018 27832
rect 18325 27829 18337 27832
rect 18371 27829 18383 27863
rect 18325 27823 18383 27829
rect 20990 27820 20996 27872
rect 21048 27820 21054 27872
rect 22554 27820 22560 27872
rect 22612 27820 22618 27872
rect 22646 27820 22652 27872
rect 22704 27820 22710 27872
rect 23032 27860 23060 27959
rect 23290 27956 23296 28008
rect 23348 27996 23354 28008
rect 23661 27999 23719 28005
rect 23661 27996 23673 27999
rect 23348 27968 23673 27996
rect 23348 27956 23354 27968
rect 23661 27965 23673 27968
rect 23707 27965 23719 27999
rect 23661 27959 23719 27965
rect 24670 27956 24676 28008
rect 24728 27996 24734 28008
rect 25409 27999 25467 28005
rect 25409 27996 25421 27999
rect 24728 27968 25421 27996
rect 24728 27956 24734 27968
rect 25409 27965 25421 27968
rect 25455 27996 25467 27999
rect 26326 27996 26332 28008
rect 25455 27968 26332 27996
rect 25455 27965 25467 27968
rect 25409 27959 25467 27965
rect 26326 27956 26332 27968
rect 26384 27956 26390 28008
rect 25866 27888 25872 27940
rect 25924 27928 25930 27940
rect 26053 27931 26111 27937
rect 26053 27928 26065 27931
rect 25924 27900 26065 27928
rect 25924 27888 25930 27900
rect 26053 27897 26065 27900
rect 26099 27897 26111 27931
rect 26053 27891 26111 27897
rect 26970 27888 26976 27940
rect 27028 27928 27034 27940
rect 27816 27928 27844 28036
rect 28442 28024 28448 28076
rect 28500 28024 28506 28076
rect 29638 28024 29644 28076
rect 29696 28024 29702 28076
rect 29914 28024 29920 28076
rect 29972 28024 29978 28076
rect 30101 28067 30159 28073
rect 30101 28033 30113 28067
rect 30147 28064 30159 28067
rect 30190 28064 30196 28076
rect 30147 28036 30196 28064
rect 30147 28033 30159 28036
rect 30101 28027 30159 28033
rect 30190 28024 30196 28036
rect 30248 28024 30254 28076
rect 30300 28036 30512 28064
rect 28534 27956 28540 28008
rect 28592 27996 28598 28008
rect 28721 27999 28779 28005
rect 28721 27996 28733 27999
rect 28592 27968 28733 27996
rect 28592 27956 28598 27968
rect 28721 27965 28733 27968
rect 28767 27965 28779 27999
rect 28721 27959 28779 27965
rect 28930 27999 28988 28005
rect 28930 27965 28942 27999
rect 28976 27996 28988 27999
rect 28976 27965 28994 27996
rect 28930 27959 28994 27965
rect 27028 27900 27200 27928
rect 27028 27888 27034 27900
rect 23106 27860 23112 27872
rect 23032 27832 23112 27860
rect 23106 27820 23112 27832
rect 23164 27820 23170 27872
rect 26234 27820 26240 27872
rect 26292 27860 26298 27872
rect 26421 27863 26479 27869
rect 26421 27860 26433 27863
rect 26292 27832 26433 27860
rect 26292 27820 26298 27832
rect 26421 27829 26433 27832
rect 26467 27829 26479 27863
rect 26421 27823 26479 27829
rect 26605 27863 26663 27869
rect 26605 27829 26617 27863
rect 26651 27860 26663 27863
rect 27062 27860 27068 27872
rect 26651 27832 27068 27860
rect 26651 27829 26663 27832
rect 26605 27823 26663 27829
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 27172 27869 27200 27900
rect 27356 27900 27844 27928
rect 28966 27940 28994 27959
rect 30006 27956 30012 28008
rect 30064 27996 30070 28008
rect 30300 27996 30328 28036
rect 30064 27968 30328 27996
rect 30064 27956 30070 27968
rect 30374 27956 30380 28008
rect 30432 27956 30438 28008
rect 30484 27996 30512 28036
rect 30558 28024 30564 28076
rect 30616 28024 30622 28076
rect 30668 28073 30696 28104
rect 31386 28092 31392 28144
rect 31444 28132 31450 28144
rect 31573 28135 31631 28141
rect 31573 28132 31585 28135
rect 31444 28104 31585 28132
rect 31444 28092 31450 28104
rect 31573 28101 31585 28104
rect 31619 28132 31631 28135
rect 31846 28132 31852 28144
rect 31619 28104 31852 28132
rect 31619 28101 31631 28104
rect 31573 28095 31631 28101
rect 31846 28092 31852 28104
rect 31904 28092 31910 28144
rect 32585 28135 32643 28141
rect 32585 28101 32597 28135
rect 32631 28132 32643 28135
rect 33318 28132 33324 28144
rect 32631 28104 33324 28132
rect 32631 28101 32643 28104
rect 32585 28095 32643 28101
rect 33318 28092 33324 28104
rect 33376 28092 33382 28144
rect 30653 28067 30711 28073
rect 30653 28033 30665 28067
rect 30699 28033 30711 28067
rect 30653 28027 30711 28033
rect 30745 28067 30803 28073
rect 30745 28033 30757 28067
rect 30791 28033 30803 28067
rect 30745 28027 30803 28033
rect 31481 28067 31539 28073
rect 31481 28033 31493 28067
rect 31527 28033 31539 28067
rect 31481 28027 31539 28033
rect 31757 28067 31815 28073
rect 31757 28033 31769 28067
rect 31803 28064 31815 28067
rect 32306 28064 32312 28076
rect 31803 28036 32312 28064
rect 31803 28033 31815 28036
rect 31757 28027 31815 28033
rect 30760 27996 30788 28027
rect 30484 27968 30788 27996
rect 30837 27999 30895 28005
rect 30837 27965 30849 27999
rect 30883 27965 30895 27999
rect 30837 27959 30895 27965
rect 31496 27996 31524 28027
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 32398 28024 32404 28076
rect 32456 28024 32462 28076
rect 32674 28024 32680 28076
rect 32732 28024 32738 28076
rect 32769 28067 32827 28073
rect 32769 28033 32781 28067
rect 32815 28033 32827 28067
rect 32769 28027 32827 28033
rect 32784 27996 32812 28027
rect 31496 27968 32812 27996
rect 28966 27900 29000 27940
rect 27356 27872 27384 27900
rect 28994 27888 29000 27900
rect 29052 27928 29058 27940
rect 29730 27928 29736 27940
rect 29052 27900 29736 27928
rect 29052 27888 29058 27900
rect 29730 27888 29736 27900
rect 29788 27888 29794 27940
rect 30285 27931 30343 27937
rect 30285 27897 30297 27931
rect 30331 27928 30343 27931
rect 30466 27928 30472 27940
rect 30331 27900 30472 27928
rect 30331 27897 30343 27900
rect 30285 27891 30343 27897
rect 30466 27888 30472 27900
rect 30524 27928 30530 27940
rect 30852 27928 30880 27959
rect 30524 27900 30880 27928
rect 30524 27888 30530 27900
rect 27157 27863 27215 27869
rect 27157 27829 27169 27863
rect 27203 27829 27215 27863
rect 27157 27823 27215 27829
rect 27338 27820 27344 27872
rect 27396 27820 27402 27872
rect 29086 27820 29092 27872
rect 29144 27820 29150 27872
rect 29362 27820 29368 27872
rect 29420 27860 29426 27872
rect 31496 27860 31524 27968
rect 29420 27832 31524 27860
rect 29420 27820 29426 27832
rect 31846 27820 31852 27872
rect 31904 27860 31910 27872
rect 31941 27863 31999 27869
rect 31941 27860 31953 27863
rect 31904 27832 31953 27860
rect 31904 27820 31910 27832
rect 31941 27829 31953 27832
rect 31987 27829 31999 27863
rect 31941 27823 31999 27829
rect 32950 27820 32956 27872
rect 33008 27820 33014 27872
rect 1104 27770 36432 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 36432 27770
rect 1104 27696 36432 27718
rect 2130 27616 2136 27668
rect 2188 27656 2194 27668
rect 4709 27659 4767 27665
rect 4709 27656 4721 27659
rect 2188 27628 4721 27656
rect 2188 27616 2194 27628
rect 4709 27625 4721 27628
rect 4755 27625 4767 27659
rect 4709 27619 4767 27625
rect 4893 27659 4951 27665
rect 4893 27625 4905 27659
rect 4939 27656 4951 27659
rect 4982 27656 4988 27668
rect 4939 27628 4988 27656
rect 4939 27625 4951 27628
rect 4893 27619 4951 27625
rect 4982 27616 4988 27628
rect 5040 27616 5046 27668
rect 5258 27616 5264 27668
rect 5316 27656 5322 27668
rect 6273 27659 6331 27665
rect 6273 27656 6285 27659
rect 5316 27628 6285 27656
rect 5316 27616 5322 27628
rect 6273 27625 6285 27628
rect 6319 27625 6331 27659
rect 6273 27619 6331 27625
rect 7377 27659 7435 27665
rect 7377 27625 7389 27659
rect 7423 27656 7435 27659
rect 7466 27656 7472 27668
rect 7423 27628 7472 27656
rect 7423 27625 7435 27628
rect 7377 27619 7435 27625
rect 2225 27591 2283 27597
rect 2225 27557 2237 27591
rect 2271 27588 2283 27591
rect 3142 27588 3148 27600
rect 2271 27560 3148 27588
rect 2271 27557 2283 27560
rect 2225 27551 2283 27557
rect 3142 27548 3148 27560
rect 3200 27548 3206 27600
rect 6288 27588 6316 27619
rect 7466 27616 7472 27628
rect 7524 27616 7530 27668
rect 7742 27616 7748 27668
rect 7800 27656 7806 27668
rect 10042 27656 10048 27668
rect 7800 27628 10048 27656
rect 7800 27616 7806 27628
rect 10042 27616 10048 27628
rect 10100 27616 10106 27668
rect 10226 27616 10232 27668
rect 10284 27656 10290 27668
rect 10321 27659 10379 27665
rect 10321 27656 10333 27659
rect 10284 27628 10333 27656
rect 10284 27616 10290 27628
rect 10321 27625 10333 27628
rect 10367 27625 10379 27659
rect 10321 27619 10379 27625
rect 11054 27616 11060 27668
rect 11112 27656 11118 27668
rect 11517 27659 11575 27665
rect 11517 27656 11529 27659
rect 11112 27628 11529 27656
rect 11112 27616 11118 27628
rect 11517 27625 11529 27628
rect 11563 27656 11575 27659
rect 11563 27628 12434 27656
rect 11563 27625 11575 27628
rect 11517 27619 11575 27625
rect 9030 27588 9036 27600
rect 6288 27560 7604 27588
rect 4522 27480 4528 27532
rect 4580 27480 4586 27532
rect 5350 27480 5356 27532
rect 5408 27520 5414 27532
rect 5445 27523 5503 27529
rect 5445 27520 5457 27523
rect 5408 27492 5457 27520
rect 5408 27480 5414 27492
rect 5445 27489 5457 27492
rect 5491 27489 5503 27523
rect 5445 27483 5503 27489
rect 5736 27492 6408 27520
rect 2406 27412 2412 27464
rect 2464 27412 2470 27464
rect 2685 27455 2743 27461
rect 2685 27421 2697 27455
rect 2731 27452 2743 27455
rect 4062 27452 4068 27464
rect 2731 27424 4068 27452
rect 2731 27421 2743 27424
rect 2685 27415 2743 27421
rect 4062 27412 4068 27424
rect 4120 27412 4126 27464
rect 4433 27455 4491 27461
rect 4433 27421 4445 27455
rect 4479 27452 4491 27455
rect 4614 27452 4620 27464
rect 4479 27424 4620 27452
rect 4479 27421 4491 27424
rect 4433 27415 4491 27421
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 5261 27455 5319 27461
rect 5261 27421 5273 27455
rect 5307 27452 5319 27455
rect 5736 27452 5764 27492
rect 5307 27424 5764 27452
rect 5902 27455 5960 27461
rect 5307 27421 5319 27424
rect 5261 27415 5319 27421
rect 5902 27421 5914 27455
rect 5948 27452 5960 27455
rect 5994 27452 6000 27464
rect 5948 27424 6000 27452
rect 5948 27421 5960 27424
rect 5902 27415 5960 27421
rect 5994 27412 6000 27424
rect 6052 27412 6058 27464
rect 6380 27461 6408 27492
rect 7374 27480 7380 27532
rect 7432 27520 7438 27532
rect 7576 27529 7604 27560
rect 7760 27560 9036 27588
rect 7561 27523 7619 27529
rect 7561 27520 7573 27523
rect 7432 27492 7573 27520
rect 7432 27480 7438 27492
rect 7561 27489 7573 27492
rect 7607 27489 7619 27523
rect 7561 27483 7619 27489
rect 6365 27455 6423 27461
rect 6365 27421 6377 27455
rect 6411 27452 6423 27455
rect 6454 27452 6460 27464
rect 6411 27424 6460 27452
rect 6411 27421 6423 27424
rect 6365 27415 6423 27421
rect 6454 27412 6460 27424
rect 6512 27412 6518 27464
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27452 7711 27455
rect 7760 27452 7788 27560
rect 9030 27548 9036 27560
rect 9088 27588 9094 27600
rect 12253 27591 12311 27597
rect 12253 27588 12265 27591
rect 9088 27560 12265 27588
rect 9088 27548 9094 27560
rect 12253 27557 12265 27560
rect 12299 27557 12311 27591
rect 12406 27588 12434 27628
rect 15194 27616 15200 27668
rect 15252 27656 15258 27668
rect 15400 27659 15458 27665
rect 15400 27656 15412 27659
rect 15252 27628 15412 27656
rect 15252 27616 15258 27628
rect 15400 27625 15412 27628
rect 15446 27625 15458 27659
rect 22186 27656 22192 27668
rect 15400 27619 15458 27625
rect 21376 27628 22192 27656
rect 13633 27591 13691 27597
rect 12406 27560 13584 27588
rect 12253 27551 12311 27557
rect 8757 27523 8815 27529
rect 8757 27489 8769 27523
rect 8803 27520 8815 27523
rect 9214 27520 9220 27532
rect 8803 27492 9220 27520
rect 8803 27489 8815 27492
rect 8757 27483 8815 27489
rect 9214 27480 9220 27492
rect 9272 27520 9278 27532
rect 9309 27523 9367 27529
rect 9309 27520 9321 27523
rect 9272 27492 9321 27520
rect 9272 27480 9278 27492
rect 9309 27489 9321 27492
rect 9355 27520 9367 27523
rect 11609 27523 11667 27529
rect 9355 27492 9628 27520
rect 9355 27489 9367 27492
rect 9309 27483 9367 27489
rect 9600 27464 9628 27492
rect 11609 27489 11621 27523
rect 11655 27520 11667 27523
rect 12342 27520 12348 27532
rect 11655 27492 12348 27520
rect 11655 27489 11667 27492
rect 11609 27483 11667 27489
rect 12342 27480 12348 27492
rect 12400 27480 12406 27532
rect 12710 27480 12716 27532
rect 12768 27520 12774 27532
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 12768 27492 13277 27520
rect 12768 27480 12774 27492
rect 13265 27489 13277 27492
rect 13311 27489 13323 27523
rect 13556 27520 13584 27560
rect 13633 27557 13645 27591
rect 13679 27588 13691 27591
rect 14274 27588 14280 27600
rect 13679 27560 14280 27588
rect 13679 27557 13691 27560
rect 13633 27551 13691 27557
rect 14274 27548 14280 27560
rect 14332 27548 14338 27600
rect 15289 27591 15347 27597
rect 15289 27557 15301 27591
rect 15335 27588 15347 27591
rect 16942 27588 16948 27600
rect 15335 27560 16948 27588
rect 15335 27557 15347 27560
rect 15289 27551 15347 27557
rect 16942 27548 16948 27560
rect 17000 27548 17006 27600
rect 17129 27591 17187 27597
rect 17129 27557 17141 27591
rect 17175 27588 17187 27591
rect 17494 27588 17500 27600
rect 17175 27560 17500 27588
rect 17175 27557 17187 27560
rect 17129 27551 17187 27557
rect 17494 27548 17500 27560
rect 17552 27548 17558 27600
rect 20714 27548 20720 27600
rect 20772 27588 20778 27600
rect 21376 27588 21404 27628
rect 22186 27616 22192 27628
rect 22244 27616 22250 27668
rect 23290 27616 23296 27668
rect 23348 27656 23354 27668
rect 23385 27659 23443 27665
rect 23385 27656 23397 27659
rect 23348 27628 23397 27656
rect 23348 27616 23354 27628
rect 23385 27625 23397 27628
rect 23431 27625 23443 27659
rect 23385 27619 23443 27625
rect 25866 27616 25872 27668
rect 25924 27656 25930 27668
rect 26053 27659 26111 27665
rect 26053 27656 26065 27659
rect 25924 27628 26065 27656
rect 25924 27616 25930 27628
rect 26053 27625 26065 27628
rect 26099 27625 26111 27659
rect 26053 27619 26111 27625
rect 26605 27659 26663 27665
rect 26605 27625 26617 27659
rect 26651 27656 26663 27659
rect 26694 27656 26700 27668
rect 26651 27628 26700 27656
rect 26651 27625 26663 27628
rect 26605 27619 26663 27625
rect 26694 27616 26700 27628
rect 26752 27616 26758 27668
rect 26881 27659 26939 27665
rect 26881 27625 26893 27659
rect 26927 27656 26939 27659
rect 27246 27656 27252 27668
rect 26927 27628 27252 27656
rect 26927 27625 26939 27628
rect 26881 27619 26939 27625
rect 27246 27616 27252 27628
rect 27304 27616 27310 27668
rect 28994 27656 29000 27668
rect 27356 27628 29000 27656
rect 20772 27560 21404 27588
rect 20772 27548 20778 27560
rect 26326 27548 26332 27600
rect 26384 27588 26390 27600
rect 27356 27588 27384 27628
rect 28994 27616 29000 27628
rect 29052 27616 29058 27668
rect 30190 27656 30196 27668
rect 29104 27628 30196 27656
rect 26384 27560 27384 27588
rect 26384 27548 26390 27560
rect 28810 27548 28816 27600
rect 28868 27588 28874 27600
rect 29104 27588 29132 27628
rect 30190 27616 30196 27628
rect 30248 27616 30254 27668
rect 30745 27659 30803 27665
rect 30745 27625 30757 27659
rect 30791 27656 30803 27659
rect 31018 27656 31024 27668
rect 30791 27628 31024 27656
rect 30791 27625 30803 27628
rect 30745 27619 30803 27625
rect 31018 27616 31024 27628
rect 31076 27616 31082 27668
rect 31662 27616 31668 27668
rect 31720 27616 31726 27668
rect 28868 27560 29132 27588
rect 28868 27548 28874 27560
rect 29178 27548 29184 27600
rect 29236 27588 29242 27600
rect 31110 27588 31116 27600
rect 29236 27560 29960 27588
rect 29236 27548 29242 27560
rect 14829 27523 14887 27529
rect 14829 27520 14841 27523
rect 13556 27492 14841 27520
rect 13265 27483 13323 27489
rect 14829 27489 14841 27492
rect 14875 27489 14887 27523
rect 14829 27483 14887 27489
rect 15197 27523 15255 27529
rect 15197 27489 15209 27523
rect 15243 27520 15255 27523
rect 15378 27520 15384 27532
rect 15243 27492 15384 27520
rect 15243 27489 15255 27492
rect 15197 27483 15255 27489
rect 15378 27480 15384 27492
rect 15436 27480 15442 27532
rect 18966 27480 18972 27532
rect 19024 27520 19030 27532
rect 19521 27523 19579 27529
rect 19521 27520 19533 27523
rect 19024 27492 19533 27520
rect 19024 27480 19030 27492
rect 19521 27489 19533 27492
rect 19567 27520 19579 27523
rect 21174 27520 21180 27532
rect 19567 27492 21180 27520
rect 19567 27489 19579 27492
rect 19521 27483 19579 27489
rect 21174 27480 21180 27492
rect 21232 27480 21238 27532
rect 23382 27520 23388 27532
rect 21284 27492 23388 27520
rect 21284 27464 21312 27492
rect 23382 27480 23388 27492
rect 23440 27480 23446 27532
rect 25130 27480 25136 27532
rect 25188 27480 25194 27532
rect 26234 27480 26240 27532
rect 26292 27480 26298 27532
rect 26602 27480 26608 27532
rect 26660 27520 26666 27532
rect 27338 27520 27344 27532
rect 26660 27492 27344 27520
rect 26660 27480 26666 27492
rect 27338 27480 27344 27492
rect 27396 27520 27402 27532
rect 29822 27520 29828 27532
rect 27396 27492 29828 27520
rect 27396 27480 27402 27492
rect 29822 27480 29828 27492
rect 29880 27480 29886 27532
rect 8573 27455 8631 27461
rect 8573 27452 8585 27455
rect 7699 27424 7788 27452
rect 7852 27424 8585 27452
rect 7699 27421 7711 27424
rect 7653 27415 7711 27421
rect 1394 27344 1400 27396
rect 1452 27384 1458 27396
rect 2593 27387 2651 27393
rect 2593 27384 2605 27387
rect 1452 27356 2605 27384
rect 1452 27344 1458 27356
rect 2593 27353 2605 27356
rect 2639 27353 2651 27387
rect 2593 27347 2651 27353
rect 4798 27344 4804 27396
rect 4856 27344 4862 27396
rect 5350 27276 5356 27328
rect 5408 27276 5414 27328
rect 5718 27276 5724 27328
rect 5776 27276 5782 27328
rect 5902 27276 5908 27328
rect 5960 27276 5966 27328
rect 6012 27316 6040 27412
rect 6086 27344 6092 27396
rect 6144 27384 6150 27396
rect 7852 27384 7880 27424
rect 8573 27421 8585 27424
rect 8619 27421 8631 27455
rect 8573 27415 8631 27421
rect 9122 27412 9128 27464
rect 9180 27412 9186 27464
rect 9490 27412 9496 27464
rect 9548 27412 9554 27464
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 10229 27455 10287 27461
rect 10229 27452 10241 27455
rect 9640 27424 10241 27452
rect 9640 27412 9646 27424
rect 10229 27421 10241 27424
rect 10275 27421 10287 27455
rect 10229 27415 10287 27421
rect 10410 27412 10416 27464
rect 10468 27412 10474 27464
rect 10778 27412 10784 27464
rect 10836 27452 10842 27464
rect 11090 27455 11148 27461
rect 11090 27452 11102 27455
rect 10836 27424 11102 27452
rect 10836 27412 10842 27424
rect 11090 27421 11102 27424
rect 11136 27421 11148 27455
rect 11090 27415 11148 27421
rect 11701 27455 11759 27461
rect 11701 27421 11713 27455
rect 11747 27421 11759 27455
rect 11701 27415 11759 27421
rect 6144 27356 7880 27384
rect 7929 27387 7987 27393
rect 6144 27344 6150 27356
rect 7929 27353 7941 27387
rect 7975 27353 7987 27387
rect 7929 27347 7987 27353
rect 7944 27316 7972 27347
rect 8018 27344 8024 27396
rect 8076 27344 8082 27396
rect 8110 27344 8116 27396
rect 8168 27384 8174 27396
rect 9401 27387 9459 27393
rect 9401 27384 9413 27387
rect 8168 27356 9413 27384
rect 8168 27344 8174 27356
rect 9401 27353 9413 27356
rect 9447 27353 9459 27387
rect 9401 27347 9459 27353
rect 11330 27344 11336 27396
rect 11388 27384 11394 27396
rect 11716 27384 11744 27415
rect 11790 27412 11796 27464
rect 11848 27452 11854 27464
rect 11848 27424 11893 27452
rect 11848 27412 11854 27424
rect 12158 27412 12164 27464
rect 12216 27412 12222 27464
rect 12434 27412 12440 27464
rect 12492 27412 12498 27464
rect 12621 27455 12679 27461
rect 12621 27421 12633 27455
rect 12667 27452 12679 27455
rect 12894 27452 12900 27464
rect 12667 27424 12900 27452
rect 12667 27421 12679 27424
rect 12621 27415 12679 27421
rect 12894 27412 12900 27424
rect 12952 27412 12958 27464
rect 12989 27455 13047 27461
rect 12989 27421 13001 27455
rect 13035 27421 13047 27455
rect 12989 27415 13047 27421
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27452 13231 27455
rect 13446 27452 13452 27464
rect 13219 27424 13452 27452
rect 13219 27421 13231 27424
rect 13173 27415 13231 27421
rect 11388 27356 11744 27384
rect 12069 27387 12127 27393
rect 11388 27344 11394 27356
rect 12069 27353 12081 27387
rect 12115 27384 12127 27387
rect 12250 27384 12256 27396
rect 12115 27356 12256 27384
rect 12115 27353 12127 27356
rect 12069 27347 12127 27353
rect 12250 27344 12256 27356
rect 12308 27344 12314 27396
rect 12526 27344 12532 27396
rect 12584 27384 12590 27396
rect 13004 27384 13032 27415
rect 13446 27412 13452 27424
rect 13504 27412 13510 27464
rect 13538 27412 13544 27464
rect 13596 27412 13602 27464
rect 13725 27455 13783 27461
rect 13725 27421 13737 27455
rect 13771 27452 13783 27455
rect 14090 27452 14096 27464
rect 13771 27424 14096 27452
rect 13771 27421 13783 27424
rect 13725 27415 13783 27421
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 14737 27455 14795 27461
rect 14737 27421 14749 27455
rect 14783 27452 14795 27455
rect 16298 27452 16304 27464
rect 14783 27424 16304 27452
rect 14783 27421 14795 27424
rect 14737 27415 14795 27421
rect 12584 27356 13032 27384
rect 13556 27384 13584 27412
rect 14185 27387 14243 27393
rect 14185 27384 14197 27387
rect 13556 27356 14197 27384
rect 12584 27344 12590 27356
rect 14185 27353 14197 27356
rect 14231 27353 14243 27387
rect 14660 27384 14688 27415
rect 16298 27412 16304 27424
rect 16356 27412 16362 27464
rect 17126 27412 17132 27464
rect 17184 27452 17190 27464
rect 18877 27455 18935 27461
rect 17184 27424 17526 27452
rect 17184 27412 17190 27424
rect 18877 27421 18889 27455
rect 18923 27421 18935 27455
rect 18877 27415 18935 27421
rect 19245 27455 19303 27461
rect 19245 27421 19257 27455
rect 19291 27452 19303 27455
rect 19426 27452 19432 27464
rect 19291 27424 19432 27452
rect 19291 27421 19303 27424
rect 19245 27415 19303 27421
rect 15470 27384 15476 27396
rect 14660 27356 15476 27384
rect 14185 27347 14243 27353
rect 15470 27344 15476 27356
rect 15528 27344 15534 27396
rect 15562 27344 15568 27396
rect 15620 27384 15626 27396
rect 17034 27384 17040 27396
rect 15620 27356 17040 27384
rect 15620 27344 15626 27356
rect 17034 27344 17040 27356
rect 17092 27344 17098 27396
rect 18598 27344 18604 27396
rect 18656 27344 18662 27396
rect 18690 27344 18696 27396
rect 18748 27384 18754 27396
rect 18892 27384 18920 27415
rect 19426 27412 19432 27424
rect 19484 27452 19490 27464
rect 19610 27452 19616 27464
rect 19484 27424 19616 27452
rect 19484 27412 19490 27424
rect 19610 27412 19616 27424
rect 19668 27412 19674 27464
rect 19978 27412 19984 27464
rect 20036 27452 20042 27464
rect 20717 27455 20775 27461
rect 20717 27452 20729 27455
rect 20036 27424 20729 27452
rect 20036 27412 20042 27424
rect 20717 27421 20729 27424
rect 20763 27421 20775 27455
rect 20717 27415 20775 27421
rect 21266 27412 21272 27464
rect 21324 27412 21330 27464
rect 23566 27412 23572 27464
rect 23624 27412 23630 27464
rect 23750 27412 23756 27464
rect 23808 27412 23814 27464
rect 23934 27412 23940 27464
rect 23992 27412 23998 27464
rect 25866 27412 25872 27464
rect 25924 27452 25930 27464
rect 25961 27455 26019 27461
rect 25961 27452 25973 27455
rect 25924 27424 25973 27452
rect 25924 27412 25930 27424
rect 25961 27421 25973 27424
rect 26007 27421 26019 27455
rect 26881 27455 26939 27461
rect 26881 27452 26893 27455
rect 25961 27415 26019 27421
rect 26252 27424 26893 27452
rect 18748 27356 18920 27384
rect 18748 27344 18754 27356
rect 21542 27344 21548 27396
rect 21600 27344 21606 27396
rect 23106 27384 23112 27396
rect 22770 27356 23112 27384
rect 23106 27344 23112 27356
rect 23164 27344 23170 27396
rect 26252 27393 26280 27424
rect 26881 27421 26893 27424
rect 26927 27421 26939 27455
rect 26881 27415 26939 27421
rect 27062 27412 27068 27464
rect 27120 27452 27126 27464
rect 27157 27455 27215 27461
rect 27157 27452 27169 27455
rect 27120 27424 27169 27452
rect 27120 27412 27126 27424
rect 27157 27421 27169 27424
rect 27203 27421 27215 27455
rect 27157 27415 27215 27421
rect 27522 27412 27528 27464
rect 27580 27452 27586 27464
rect 29932 27461 29960 27560
rect 30668 27560 31116 27588
rect 30668 27532 30696 27560
rect 31110 27548 31116 27560
rect 31168 27548 31174 27600
rect 31202 27548 31208 27600
rect 31260 27588 31266 27600
rect 31389 27591 31447 27597
rect 31389 27588 31401 27591
rect 31260 27560 31401 27588
rect 31260 27548 31266 27560
rect 31389 27557 31401 27560
rect 31435 27557 31447 27591
rect 31389 27551 31447 27557
rect 31478 27548 31484 27600
rect 31536 27588 31542 27600
rect 34606 27588 34612 27600
rect 31536 27560 34612 27588
rect 31536 27548 31542 27560
rect 34606 27548 34612 27560
rect 34664 27548 34670 27600
rect 30009 27523 30067 27529
rect 30009 27489 30021 27523
rect 30055 27520 30067 27523
rect 30098 27520 30104 27532
rect 30055 27492 30104 27520
rect 30055 27489 30067 27492
rect 30009 27483 30067 27489
rect 30098 27480 30104 27492
rect 30156 27480 30162 27532
rect 30377 27523 30435 27529
rect 30377 27489 30389 27523
rect 30423 27520 30435 27523
rect 30650 27520 30656 27532
rect 30423 27492 30656 27520
rect 30423 27489 30435 27492
rect 30377 27483 30435 27489
rect 30650 27480 30656 27492
rect 30708 27480 30714 27532
rect 30926 27480 30932 27532
rect 30984 27520 30990 27532
rect 30984 27492 31248 27520
rect 30984 27480 30990 27492
rect 29733 27455 29791 27461
rect 29733 27452 29745 27455
rect 27580 27424 29745 27452
rect 27580 27412 27586 27424
rect 29733 27421 29745 27424
rect 29779 27421 29791 27455
rect 29733 27415 29791 27421
rect 29917 27455 29975 27461
rect 29917 27421 29929 27455
rect 29963 27452 29975 27455
rect 31018 27452 31024 27464
rect 29963 27424 31024 27452
rect 29963 27421 29975 27424
rect 29917 27415 29975 27421
rect 31018 27412 31024 27424
rect 31076 27412 31082 27464
rect 31220 27461 31248 27492
rect 31205 27455 31263 27461
rect 31205 27421 31217 27455
rect 31251 27421 31263 27455
rect 31205 27415 31263 27421
rect 31665 27455 31723 27461
rect 31665 27421 31677 27455
rect 31711 27421 31723 27455
rect 31665 27415 31723 27421
rect 23293 27387 23351 27393
rect 23293 27353 23305 27387
rect 23339 27353 23351 27387
rect 23293 27347 23351 27353
rect 23661 27387 23719 27393
rect 23661 27353 23673 27387
rect 23707 27353 23719 27387
rect 23661 27347 23719 27353
rect 26237 27387 26295 27393
rect 26237 27353 26249 27387
rect 26283 27353 26295 27387
rect 26789 27387 26847 27393
rect 26237 27347 26295 27353
rect 26436 27356 26740 27384
rect 10778 27316 10784 27328
rect 6012 27288 10784 27316
rect 10778 27276 10784 27288
rect 10836 27276 10842 27328
rect 10962 27276 10968 27328
rect 11020 27276 11026 27328
rect 11149 27319 11207 27325
rect 11149 27285 11161 27319
rect 11195 27316 11207 27319
rect 11238 27316 11244 27328
rect 11195 27288 11244 27316
rect 11195 27285 11207 27288
rect 11149 27279 11207 27285
rect 11238 27276 11244 27288
rect 11296 27316 11302 27328
rect 11698 27316 11704 27328
rect 11296 27288 11704 27316
rect 11296 27276 11302 27288
rect 11698 27276 11704 27288
rect 11756 27276 11762 27328
rect 16298 27276 16304 27328
rect 16356 27316 16362 27328
rect 18322 27316 18328 27328
rect 16356 27288 18328 27316
rect 16356 27276 16362 27288
rect 18322 27276 18328 27288
rect 18380 27276 18386 27328
rect 18506 27276 18512 27328
rect 18564 27316 18570 27328
rect 20165 27319 20223 27325
rect 20165 27316 20177 27319
rect 18564 27288 20177 27316
rect 18564 27276 18570 27288
rect 20165 27285 20177 27288
rect 20211 27285 20223 27319
rect 20165 27279 20223 27285
rect 20898 27276 20904 27328
rect 20956 27316 20962 27328
rect 21910 27316 21916 27328
rect 20956 27288 21916 27316
rect 20956 27276 20962 27288
rect 21910 27276 21916 27288
rect 21968 27316 21974 27328
rect 22830 27316 22836 27328
rect 21968 27288 22836 27316
rect 21968 27276 21974 27288
rect 22830 27276 22836 27288
rect 22888 27316 22894 27328
rect 23308 27316 23336 27347
rect 22888 27288 23336 27316
rect 23676 27316 23704 27347
rect 24489 27319 24547 27325
rect 24489 27316 24501 27319
rect 23676 27288 24501 27316
rect 22888 27276 22894 27288
rect 24489 27285 24501 27288
rect 24535 27285 24547 27319
rect 24489 27279 24547 27285
rect 26050 27276 26056 27328
rect 26108 27316 26114 27328
rect 26252 27316 26280 27347
rect 26436 27325 26464 27356
rect 26108 27288 26280 27316
rect 26421 27319 26479 27325
rect 26108 27276 26114 27288
rect 26421 27285 26433 27319
rect 26467 27285 26479 27319
rect 26421 27279 26479 27285
rect 26602 27276 26608 27328
rect 26660 27276 26666 27328
rect 26712 27316 26740 27356
rect 26789 27353 26801 27387
rect 26835 27384 26847 27387
rect 27246 27384 27252 27396
rect 26835 27356 27252 27384
rect 26835 27353 26847 27356
rect 26789 27347 26847 27353
rect 27246 27344 27252 27356
rect 27304 27344 27310 27396
rect 29086 27344 29092 27396
rect 29144 27384 29150 27396
rect 31680 27384 31708 27415
rect 31846 27412 31852 27464
rect 31904 27412 31910 27464
rect 29144 27356 31708 27384
rect 29144 27344 29150 27356
rect 26878 27316 26884 27328
rect 26712 27288 26884 27316
rect 26878 27276 26884 27288
rect 26936 27276 26942 27328
rect 27065 27319 27123 27325
rect 27065 27285 27077 27319
rect 27111 27316 27123 27319
rect 27798 27316 27804 27328
rect 27111 27288 27804 27316
rect 27111 27285 27123 27288
rect 27065 27279 27123 27285
rect 27798 27276 27804 27288
rect 27856 27276 27862 27328
rect 29549 27319 29607 27325
rect 29549 27285 29561 27319
rect 29595 27316 29607 27319
rect 30098 27316 30104 27328
rect 29595 27288 30104 27316
rect 29595 27285 29607 27288
rect 29549 27279 29607 27285
rect 30098 27276 30104 27288
rect 30156 27276 30162 27328
rect 30742 27276 30748 27328
rect 30800 27276 30806 27328
rect 30926 27276 30932 27328
rect 30984 27276 30990 27328
rect 32033 27319 32091 27325
rect 32033 27285 32045 27319
rect 32079 27316 32091 27319
rect 33502 27316 33508 27328
rect 32079 27288 33508 27316
rect 32079 27285 32091 27288
rect 32033 27279 32091 27285
rect 33502 27276 33508 27288
rect 33560 27276 33566 27328
rect 1104 27226 36432 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 36432 27226
rect 1104 27152 36432 27174
rect 2866 27112 2872 27124
rect 2240 27084 2872 27112
rect 2240 26985 2268 27084
rect 2866 27072 2872 27084
rect 2924 27112 2930 27124
rect 3418 27112 3424 27124
rect 2924 27084 3424 27112
rect 2924 27072 2930 27084
rect 3418 27072 3424 27084
rect 3476 27072 3482 27124
rect 4614 27072 4620 27124
rect 4672 27112 4678 27124
rect 7926 27112 7932 27124
rect 4672 27084 7932 27112
rect 4672 27072 4678 27084
rect 7926 27072 7932 27084
rect 7984 27112 7990 27124
rect 8110 27112 8116 27124
rect 7984 27084 8116 27112
rect 7984 27072 7990 27084
rect 8110 27072 8116 27084
rect 8168 27072 8174 27124
rect 9309 27115 9367 27121
rect 9309 27081 9321 27115
rect 9355 27112 9367 27115
rect 9490 27112 9496 27124
rect 9355 27084 9496 27112
rect 9355 27081 9367 27084
rect 9309 27075 9367 27081
rect 9490 27072 9496 27084
rect 9548 27072 9554 27124
rect 10870 27072 10876 27124
rect 10928 27112 10934 27124
rect 10928 27084 12434 27112
rect 10928 27072 10934 27084
rect 2774 27004 2780 27056
rect 2832 27044 2838 27056
rect 5169 27047 5227 27053
rect 2832 27016 2990 27044
rect 2832 27004 2838 27016
rect 5169 27013 5181 27047
rect 5215 27044 5227 27047
rect 5350 27044 5356 27056
rect 5215 27016 5356 27044
rect 5215 27013 5227 27016
rect 5169 27007 5227 27013
rect 5350 27004 5356 27016
rect 5408 27004 5414 27056
rect 6454 27004 6460 27056
rect 6512 27044 6518 27056
rect 12253 27047 12311 27053
rect 12253 27044 12265 27047
rect 6512 27016 12265 27044
rect 6512 27004 6518 27016
rect 12253 27013 12265 27016
rect 12299 27013 12311 27047
rect 12406 27044 12434 27084
rect 12986 27072 12992 27124
rect 13044 27112 13050 27124
rect 13354 27112 13360 27124
rect 13044 27084 13360 27112
rect 13044 27072 13050 27084
rect 13354 27072 13360 27084
rect 13412 27072 13418 27124
rect 14734 27072 14740 27124
rect 14792 27072 14798 27124
rect 16482 27112 16488 27124
rect 14844 27084 16488 27112
rect 12526 27044 12532 27056
rect 12406 27016 12532 27044
rect 12253 27007 12311 27013
rect 12526 27004 12532 27016
rect 12584 27004 12590 27056
rect 12710 27004 12716 27056
rect 12768 27044 12774 27056
rect 14752 27044 14780 27072
rect 12768 27016 14780 27044
rect 12768 27004 12774 27016
rect 2225 26979 2283 26985
rect 2225 26945 2237 26979
rect 2271 26945 2283 26979
rect 2225 26939 2283 26945
rect 4801 26979 4859 26985
rect 4801 26945 4813 26979
rect 4847 26976 4859 26979
rect 5718 26976 5724 26988
rect 4847 26948 5724 26976
rect 4847 26945 4859 26948
rect 4801 26939 4859 26945
rect 5718 26936 5724 26948
rect 5776 26936 5782 26988
rect 7101 26979 7159 26985
rect 7101 26945 7113 26979
rect 7147 26976 7159 26979
rect 7190 26976 7196 26988
rect 7147 26948 7196 26976
rect 7147 26945 7159 26948
rect 7101 26939 7159 26945
rect 7190 26936 7196 26948
rect 7248 26936 7254 26988
rect 7282 26936 7288 26988
rect 7340 26936 7346 26988
rect 7650 26936 7656 26988
rect 7708 26976 7714 26988
rect 7745 26979 7803 26985
rect 7745 26976 7757 26979
rect 7708 26948 7757 26976
rect 7708 26936 7714 26948
rect 7745 26945 7757 26948
rect 7791 26945 7803 26979
rect 7745 26939 7803 26945
rect 8941 26979 8999 26985
rect 8941 26945 8953 26979
rect 8987 26976 8999 26979
rect 9122 26976 9128 26988
rect 8987 26948 9128 26976
rect 8987 26945 8999 26948
rect 8941 26939 8999 26945
rect 9122 26936 9128 26948
rect 9180 26936 9186 26988
rect 10965 26979 11023 26985
rect 10965 26945 10977 26979
rect 11011 26945 11023 26979
rect 10965 26939 11023 26945
rect 2501 26911 2559 26917
rect 2501 26877 2513 26911
rect 2547 26908 2559 26911
rect 3694 26908 3700 26920
rect 2547 26880 3700 26908
rect 2547 26877 2559 26880
rect 2501 26871 2559 26877
rect 3694 26868 3700 26880
rect 3752 26868 3758 26920
rect 4522 26868 4528 26920
rect 4580 26908 4586 26920
rect 4982 26908 4988 26920
rect 4580 26880 4988 26908
rect 4580 26868 4586 26880
rect 4982 26868 4988 26880
rect 5040 26868 5046 26920
rect 7466 26908 7472 26920
rect 5092 26880 7472 26908
rect 3973 26843 4031 26849
rect 3973 26809 3985 26843
rect 4019 26840 4031 26843
rect 4062 26840 4068 26852
rect 4019 26812 4068 26840
rect 4019 26809 4031 26812
rect 3973 26803 4031 26809
rect 4062 26800 4068 26812
rect 4120 26840 4126 26852
rect 5092 26840 5120 26880
rect 7466 26868 7472 26880
rect 7524 26868 7530 26920
rect 9033 26911 9091 26917
rect 9033 26877 9045 26911
rect 9079 26877 9091 26911
rect 9033 26871 9091 26877
rect 10781 26911 10839 26917
rect 10781 26877 10793 26911
rect 10827 26877 10839 26911
rect 10781 26871 10839 26877
rect 4120 26812 5120 26840
rect 4120 26800 4126 26812
rect 5258 26800 5264 26852
rect 5316 26840 5322 26852
rect 7745 26843 7803 26849
rect 7745 26840 7757 26843
rect 5316 26812 7757 26840
rect 5316 26800 5322 26812
rect 7745 26809 7757 26812
rect 7791 26809 7803 26843
rect 7745 26803 7803 26809
rect 9048 26784 9076 26871
rect 9582 26800 9588 26852
rect 9640 26840 9646 26852
rect 10796 26840 10824 26871
rect 10980 26852 11008 26939
rect 11330 26936 11336 26988
rect 11388 26936 11394 26988
rect 12158 26936 12164 26988
rect 12216 26936 12222 26988
rect 12621 26979 12679 26985
rect 12621 26945 12633 26979
rect 12667 26976 12679 26979
rect 12894 26976 12900 26988
rect 12667 26948 12900 26976
rect 12667 26945 12679 26948
rect 12621 26939 12679 26945
rect 12894 26936 12900 26948
rect 12952 26936 12958 26988
rect 13004 26985 13032 27016
rect 12989 26979 13047 26985
rect 12989 26945 13001 26979
rect 13035 26945 13047 26979
rect 12989 26939 13047 26945
rect 13173 26979 13231 26985
rect 13173 26945 13185 26979
rect 13219 26976 13231 26979
rect 13446 26976 13452 26988
rect 13219 26948 13452 26976
rect 13219 26945 13231 26948
rect 13173 26939 13231 26945
rect 13446 26936 13452 26948
rect 13504 26936 13510 26988
rect 14182 26936 14188 26988
rect 14240 26976 14246 26988
rect 14645 26979 14703 26985
rect 14645 26976 14657 26979
rect 14240 26948 14657 26976
rect 14240 26936 14246 26948
rect 14645 26945 14657 26948
rect 14691 26945 14703 26979
rect 14645 26939 14703 26945
rect 14737 26979 14795 26985
rect 14737 26945 14749 26979
rect 14783 26976 14795 26979
rect 14844 26976 14872 27084
rect 16482 27072 16488 27084
rect 16540 27072 16546 27124
rect 17773 27115 17831 27121
rect 17773 27081 17785 27115
rect 17819 27112 17831 27115
rect 18598 27112 18604 27124
rect 17819 27084 18604 27112
rect 17819 27081 17831 27084
rect 17773 27075 17831 27081
rect 18598 27072 18604 27084
rect 18656 27072 18662 27124
rect 21177 27115 21235 27121
rect 21177 27081 21189 27115
rect 21223 27112 21235 27115
rect 21542 27112 21548 27124
rect 21223 27084 21548 27112
rect 21223 27081 21235 27084
rect 21177 27075 21235 27081
rect 21542 27072 21548 27084
rect 21600 27072 21606 27124
rect 23106 27112 23112 27124
rect 22388 27084 23112 27112
rect 18506 27044 18512 27056
rect 18064 27016 18512 27044
rect 14783 26948 14872 26976
rect 14921 26979 14979 26985
rect 14783 26945 14795 26948
rect 14737 26939 14795 26945
rect 14921 26945 14933 26979
rect 14967 26976 14979 26979
rect 16390 26976 16396 26988
rect 14967 26948 16396 26976
rect 14967 26945 14979 26948
rect 14921 26939 14979 26945
rect 12713 26911 12771 26917
rect 12713 26877 12725 26911
rect 12759 26877 12771 26911
rect 12713 26871 12771 26877
rect 9640 26812 10824 26840
rect 9640 26800 9646 26812
rect 10962 26800 10968 26852
rect 11020 26800 11026 26852
rect 11146 26800 11152 26852
rect 11204 26800 11210 26852
rect 12728 26840 12756 26871
rect 14366 26868 14372 26920
rect 14424 26868 14430 26920
rect 14660 26908 14688 26939
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 16574 26936 16580 26988
rect 16632 26976 16638 26988
rect 16669 26979 16727 26985
rect 16669 26976 16681 26979
rect 16632 26948 16681 26976
rect 16632 26936 16638 26948
rect 16669 26945 16681 26948
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 16945 26979 17003 26985
rect 16945 26945 16957 26979
rect 16991 26976 17003 26979
rect 16991 26948 17172 26976
rect 16991 26945 17003 26948
rect 16945 26939 17003 26945
rect 14829 26911 14887 26917
rect 14829 26908 14841 26911
rect 14660 26880 14841 26908
rect 14829 26877 14841 26880
rect 14875 26877 14887 26911
rect 14829 26871 14887 26877
rect 16022 26868 16028 26920
rect 16080 26908 16086 26920
rect 17037 26911 17095 26917
rect 17037 26908 17049 26911
rect 16080 26880 17049 26908
rect 16080 26868 16086 26880
rect 17037 26877 17049 26880
rect 17083 26877 17095 26911
rect 17144 26908 17172 26948
rect 17218 26936 17224 26988
rect 17276 26936 17282 26988
rect 17402 26936 17408 26988
rect 17460 26936 17466 26988
rect 17494 26936 17500 26988
rect 17552 26976 17558 26988
rect 17681 26979 17739 26985
rect 17681 26976 17693 26979
rect 17552 26948 17693 26976
rect 17552 26936 17558 26948
rect 17681 26945 17693 26948
rect 17727 26945 17739 26979
rect 17681 26939 17739 26945
rect 17865 26979 17923 26985
rect 17865 26945 17877 26979
rect 17911 26976 17923 26979
rect 17954 26976 17960 26988
rect 17911 26948 17960 26976
rect 17911 26945 17923 26948
rect 17865 26939 17923 26945
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 18064 26985 18092 27016
rect 18506 27004 18512 27016
rect 18564 27004 18570 27056
rect 18966 27044 18972 27056
rect 18616 27016 18972 27044
rect 18616 26988 18644 27016
rect 18966 27004 18972 27016
rect 19024 27004 19030 27056
rect 22388 27044 22416 27084
rect 23106 27072 23112 27084
rect 23164 27112 23170 27124
rect 24473 27115 24531 27121
rect 23164 27084 23612 27112
rect 23164 27072 23170 27084
rect 20194 27016 22416 27044
rect 22465 27047 22523 27053
rect 22465 27013 22477 27047
rect 22511 27044 22523 27047
rect 22554 27044 22560 27056
rect 22511 27016 22560 27044
rect 22511 27013 22523 27016
rect 22465 27007 22523 27013
rect 22554 27004 22560 27016
rect 22612 27004 22618 27056
rect 18049 26979 18107 26985
rect 18049 26945 18061 26979
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 18138 26936 18144 26988
rect 18196 26976 18202 26988
rect 18233 26979 18291 26985
rect 18233 26976 18245 26979
rect 18196 26948 18245 26976
rect 18196 26936 18202 26948
rect 18233 26945 18245 26948
rect 18279 26945 18291 26979
rect 18233 26939 18291 26945
rect 18325 26979 18383 26985
rect 18325 26945 18337 26979
rect 18371 26945 18383 26979
rect 18325 26939 18383 26945
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26976 18475 26979
rect 18598 26976 18604 26988
rect 18463 26948 18604 26976
rect 18463 26945 18475 26948
rect 18417 26939 18475 26945
rect 17310 26908 17316 26920
rect 17144 26880 17316 26908
rect 17037 26871 17095 26877
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 14734 26840 14740 26852
rect 12728 26812 14740 26840
rect 14734 26800 14740 26812
rect 14792 26800 14798 26852
rect 5077 26775 5135 26781
rect 5077 26741 5089 26775
rect 5123 26772 5135 26775
rect 5442 26772 5448 26784
rect 5123 26744 5448 26772
rect 5123 26741 5135 26744
rect 5077 26735 5135 26741
rect 5442 26732 5448 26744
rect 5500 26732 5506 26784
rect 7282 26732 7288 26784
rect 7340 26772 7346 26784
rect 8941 26775 8999 26781
rect 8941 26772 8953 26775
rect 7340 26744 8953 26772
rect 7340 26732 7346 26744
rect 8941 26741 8953 26744
rect 8987 26741 8999 26775
rect 8941 26735 8999 26741
rect 9030 26732 9036 26784
rect 9088 26772 9094 26784
rect 13354 26772 13360 26784
rect 9088 26744 13360 26772
rect 9088 26732 9094 26744
rect 13354 26732 13360 26744
rect 13412 26732 13418 26784
rect 13722 26732 13728 26784
rect 13780 26772 13786 26784
rect 16942 26772 16948 26784
rect 13780 26744 16948 26772
rect 13780 26732 13786 26744
rect 16942 26732 16948 26744
rect 17000 26732 17006 26784
rect 18340 26772 18368 26939
rect 18598 26936 18604 26948
rect 18656 26936 18662 26988
rect 18690 26936 18696 26988
rect 18748 26936 18754 26988
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26945 20683 26979
rect 20625 26939 20683 26945
rect 18969 26911 19027 26917
rect 18969 26908 18981 26911
rect 18616 26880 18981 26908
rect 18616 26849 18644 26880
rect 18969 26877 18981 26880
rect 19015 26877 19027 26911
rect 20640 26908 20668 26939
rect 20714 26936 20720 26988
rect 20772 26976 20778 26988
rect 20809 26979 20867 26985
rect 20809 26976 20821 26979
rect 20772 26948 20821 26976
rect 20772 26936 20778 26948
rect 20809 26945 20821 26948
rect 20855 26945 20867 26979
rect 20809 26939 20867 26945
rect 20898 26936 20904 26988
rect 20956 26936 20962 26988
rect 20993 26979 21051 26985
rect 20993 26945 21005 26979
rect 21039 26976 21051 26979
rect 21082 26976 21088 26988
rect 21039 26948 21088 26976
rect 21039 26945 21051 26948
rect 20993 26939 21051 26945
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26976 21327 26979
rect 23584 26976 23612 27084
rect 24473 27081 24485 27115
rect 24519 27112 24531 27115
rect 24946 27112 24952 27124
rect 24519 27084 24952 27112
rect 24519 27081 24531 27084
rect 24473 27075 24531 27081
rect 24946 27072 24952 27084
rect 25004 27072 25010 27124
rect 25038 27072 25044 27124
rect 25096 27112 25102 27124
rect 31478 27112 31484 27124
rect 25096 27084 31484 27112
rect 25096 27072 25102 27084
rect 31478 27072 31484 27084
rect 31536 27072 31542 27124
rect 24673 27047 24731 27053
rect 24673 27013 24685 27047
rect 24719 27044 24731 27047
rect 25130 27044 25136 27056
rect 24719 27016 25136 27044
rect 24719 27013 24731 27016
rect 24673 27007 24731 27013
rect 25130 27004 25136 27016
rect 25188 27004 25194 27056
rect 26145 27047 26203 27053
rect 26145 27013 26157 27047
rect 26191 27044 26203 27047
rect 26191 27016 26556 27044
rect 26191 27013 26203 27016
rect 26145 27007 26203 27013
rect 24762 26976 24768 26988
rect 21315 26948 22140 26976
rect 23584 26962 24768 26976
rect 23598 26948 24768 26962
rect 21315 26945 21327 26948
rect 21269 26939 21327 26945
rect 21450 26908 21456 26920
rect 20640 26880 21456 26908
rect 18969 26871 19027 26877
rect 21450 26868 21456 26880
rect 21508 26868 21514 26920
rect 21545 26911 21603 26917
rect 21545 26877 21557 26911
rect 21591 26908 21603 26911
rect 21818 26908 21824 26920
rect 21591 26880 21824 26908
rect 21591 26877 21603 26880
rect 21545 26871 21603 26877
rect 21818 26868 21824 26880
rect 21876 26868 21882 26920
rect 18601 26843 18659 26849
rect 18601 26809 18613 26843
rect 18647 26809 18659 26843
rect 18601 26803 18659 26809
rect 20346 26800 20352 26852
rect 20404 26840 20410 26852
rect 21269 26843 21327 26849
rect 21269 26840 21281 26843
rect 20404 26812 21281 26840
rect 20404 26800 20410 26812
rect 21269 26809 21281 26812
rect 21315 26809 21327 26843
rect 21269 26803 21327 26809
rect 21361 26843 21419 26849
rect 21361 26809 21373 26843
rect 21407 26840 21419 26843
rect 22002 26840 22008 26852
rect 21407 26812 22008 26840
rect 21407 26809 21419 26812
rect 21361 26803 21419 26809
rect 22002 26800 22008 26812
rect 22060 26800 22066 26852
rect 19518 26772 19524 26784
rect 18340 26744 19524 26772
rect 19518 26732 19524 26744
rect 19576 26732 19582 26784
rect 19978 26732 19984 26784
rect 20036 26772 20042 26784
rect 20441 26775 20499 26781
rect 20441 26772 20453 26775
rect 20036 26744 20453 26772
rect 20036 26732 20042 26744
rect 20441 26741 20453 26744
rect 20487 26741 20499 26775
rect 22112 26772 22140 26948
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 26050 26936 26056 26988
rect 26108 26936 26114 26988
rect 26234 26936 26240 26988
rect 26292 26936 26298 26988
rect 26418 26985 26424 26988
rect 26375 26979 26424 26985
rect 26375 26945 26387 26979
rect 26421 26945 26424 26979
rect 26375 26939 26424 26945
rect 26418 26936 26424 26939
rect 26476 26936 26482 26988
rect 26528 26976 26556 27016
rect 27154 27004 27160 27056
rect 27212 27044 27218 27056
rect 32674 27044 32680 27056
rect 27212 27016 32680 27044
rect 27212 27004 27218 27016
rect 32674 27004 32680 27016
rect 32732 27004 32738 27056
rect 34422 27004 34428 27056
rect 34480 27044 34486 27056
rect 34480 27016 35020 27044
rect 34480 27004 34486 27016
rect 27430 26976 27436 26988
rect 26528 26948 27436 26976
rect 27430 26936 27436 26948
rect 27488 26936 27494 26988
rect 27522 26936 27528 26988
rect 27580 26936 27586 26988
rect 31662 26936 31668 26988
rect 31720 26976 31726 26988
rect 33134 26976 33140 26988
rect 31720 26948 33140 26976
rect 31720 26936 31726 26948
rect 33134 26936 33140 26948
rect 33192 26936 33198 26988
rect 33962 26936 33968 26988
rect 34020 26976 34026 26988
rect 34517 26979 34575 26985
rect 34517 26976 34529 26979
rect 34020 26948 34529 26976
rect 34020 26936 34026 26948
rect 34517 26945 34529 26948
rect 34563 26945 34575 26979
rect 34517 26939 34575 26945
rect 34610 26979 34668 26985
rect 34610 26945 34622 26979
rect 34656 26976 34668 26979
rect 34698 26976 34704 26988
rect 34656 26948 34704 26976
rect 34656 26945 34668 26948
rect 34610 26939 34668 26945
rect 22186 26868 22192 26920
rect 22244 26868 22250 26920
rect 22554 26868 22560 26920
rect 22612 26908 22618 26920
rect 22922 26908 22928 26920
rect 22612 26880 22928 26908
rect 22612 26868 22618 26880
rect 22922 26868 22928 26880
rect 22980 26908 22986 26920
rect 23934 26908 23940 26920
rect 22980 26880 23940 26908
rect 22980 26868 22986 26880
rect 23934 26868 23940 26880
rect 23992 26908 23998 26920
rect 24213 26911 24271 26917
rect 24213 26908 24225 26911
rect 23992 26880 24225 26908
rect 23992 26868 23998 26880
rect 24213 26877 24225 26880
rect 24259 26877 24271 26911
rect 24213 26871 24271 26877
rect 26513 26911 26571 26917
rect 26513 26877 26525 26911
rect 26559 26908 26571 26911
rect 27540 26908 27568 26936
rect 26559 26880 27568 26908
rect 26559 26877 26571 26880
rect 26513 26871 26571 26877
rect 27614 26868 27620 26920
rect 27672 26908 27678 26920
rect 27672 26880 28672 26908
rect 27672 26868 27678 26880
rect 24762 26800 24768 26852
rect 24820 26840 24826 26852
rect 28644 26840 28672 26880
rect 31202 26868 31208 26920
rect 31260 26908 31266 26920
rect 31570 26908 31576 26920
rect 31260 26880 31576 26908
rect 31260 26868 31266 26880
rect 31570 26868 31576 26880
rect 31628 26908 31634 26920
rect 34624 26908 34652 26939
rect 34698 26936 34704 26948
rect 34756 26936 34762 26988
rect 34992 26985 35020 27016
rect 34793 26979 34851 26985
rect 34793 26945 34805 26979
rect 34839 26945 34851 26979
rect 34793 26939 34851 26945
rect 34885 26979 34943 26985
rect 34885 26945 34897 26979
rect 34931 26945 34943 26979
rect 34885 26939 34943 26945
rect 34982 26979 35040 26985
rect 34982 26945 34994 26979
rect 35028 26945 35040 26979
rect 34982 26939 35040 26945
rect 34808 26908 34836 26939
rect 31628 26880 34652 26908
rect 34716 26880 34836 26908
rect 34900 26908 34928 26939
rect 34900 26880 35480 26908
rect 31628 26868 31634 26880
rect 32030 26840 32036 26852
rect 24820 26812 28580 26840
rect 28644 26812 32036 26840
rect 24820 26800 24826 26812
rect 23198 26772 23204 26784
rect 22112 26744 23204 26772
rect 20441 26735 20499 26741
rect 23198 26732 23204 26744
rect 23256 26732 23262 26784
rect 23474 26732 23480 26784
rect 23532 26772 23538 26784
rect 24305 26775 24363 26781
rect 24305 26772 24317 26775
rect 23532 26744 24317 26772
rect 23532 26732 23538 26744
rect 24305 26741 24317 26744
rect 24351 26741 24363 26775
rect 24305 26735 24363 26741
rect 24486 26732 24492 26784
rect 24544 26732 24550 26784
rect 25869 26775 25927 26781
rect 25869 26741 25881 26775
rect 25915 26772 25927 26775
rect 25958 26772 25964 26784
rect 25915 26744 25964 26772
rect 25915 26741 25927 26744
rect 25869 26735 25927 26741
rect 25958 26732 25964 26744
rect 26016 26732 26022 26784
rect 26786 26732 26792 26784
rect 26844 26772 26850 26784
rect 27154 26772 27160 26784
rect 26844 26744 27160 26772
rect 26844 26732 26850 26744
rect 27154 26732 27160 26744
rect 27212 26772 27218 26784
rect 27433 26775 27491 26781
rect 27433 26772 27445 26775
rect 27212 26744 27445 26772
rect 27212 26732 27218 26744
rect 27433 26741 27445 26744
rect 27479 26741 27491 26775
rect 27433 26735 27491 26741
rect 27801 26775 27859 26781
rect 27801 26741 27813 26775
rect 27847 26772 27859 26775
rect 28442 26772 28448 26784
rect 27847 26744 28448 26772
rect 27847 26741 27859 26744
rect 27801 26735 27859 26741
rect 28442 26732 28448 26744
rect 28500 26732 28506 26784
rect 28552 26772 28580 26812
rect 32030 26800 32036 26812
rect 32088 26800 32094 26852
rect 34606 26800 34612 26852
rect 34664 26840 34670 26852
rect 34716 26840 34744 26880
rect 34664 26812 34744 26840
rect 34664 26800 34670 26812
rect 35452 26784 35480 26880
rect 32490 26772 32496 26784
rect 28552 26744 32496 26772
rect 32490 26732 32496 26744
rect 32548 26732 32554 26784
rect 35161 26775 35219 26781
rect 35161 26741 35173 26775
rect 35207 26772 35219 26775
rect 35342 26772 35348 26784
rect 35207 26744 35348 26772
rect 35207 26741 35219 26744
rect 35161 26735 35219 26741
rect 35342 26732 35348 26744
rect 35400 26732 35406 26784
rect 35434 26732 35440 26784
rect 35492 26732 35498 26784
rect 1104 26682 36432 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 36432 26682
rect 1104 26608 36432 26630
rect 1660 26571 1718 26577
rect 1660 26537 1672 26571
rect 1706 26568 1718 26571
rect 1706 26540 2774 26568
rect 1706 26537 1718 26540
rect 1660 26531 1718 26537
rect 2746 26500 2774 26540
rect 3694 26528 3700 26580
rect 3752 26568 3758 26580
rect 3789 26571 3847 26577
rect 3789 26568 3801 26571
rect 3752 26540 3801 26568
rect 3752 26528 3758 26540
rect 3789 26537 3801 26540
rect 3835 26537 3847 26571
rect 3789 26531 3847 26537
rect 5261 26571 5319 26577
rect 5261 26537 5273 26571
rect 5307 26568 5319 26571
rect 5350 26568 5356 26580
rect 5307 26540 5356 26568
rect 5307 26537 5319 26540
rect 5261 26531 5319 26537
rect 5350 26528 5356 26540
rect 5408 26528 5414 26580
rect 5721 26571 5779 26577
rect 5721 26537 5733 26571
rect 5767 26568 5779 26571
rect 5994 26568 6000 26580
rect 5767 26540 6000 26568
rect 5767 26537 5779 26540
rect 5721 26531 5779 26537
rect 5994 26528 6000 26540
rect 6052 26528 6058 26580
rect 6273 26571 6331 26577
rect 6273 26537 6285 26571
rect 6319 26568 6331 26571
rect 6454 26568 6460 26580
rect 6319 26540 6460 26568
rect 6319 26537 6331 26540
rect 6273 26531 6331 26537
rect 6454 26528 6460 26540
rect 6512 26568 6518 26580
rect 7282 26568 7288 26580
rect 6512 26540 7288 26568
rect 6512 26528 6518 26540
rect 7282 26528 7288 26540
rect 7340 26568 7346 26580
rect 7377 26571 7435 26577
rect 7377 26568 7389 26571
rect 7340 26540 7389 26568
rect 7340 26528 7346 26540
rect 7377 26537 7389 26540
rect 7423 26537 7435 26571
rect 7377 26531 7435 26537
rect 7466 26528 7472 26580
rect 7524 26528 7530 26580
rect 7650 26528 7656 26580
rect 7708 26568 7714 26580
rect 7745 26571 7803 26577
rect 7745 26568 7757 26571
rect 7708 26540 7757 26568
rect 7708 26528 7714 26540
rect 7745 26537 7757 26540
rect 7791 26537 7803 26571
rect 7745 26531 7803 26537
rect 11149 26571 11207 26577
rect 11149 26537 11161 26571
rect 11195 26568 11207 26571
rect 11330 26568 11336 26580
rect 11195 26540 11336 26568
rect 11195 26537 11207 26540
rect 11149 26531 11207 26537
rect 11330 26528 11336 26540
rect 11388 26528 11394 26580
rect 11514 26528 11520 26580
rect 11572 26528 11578 26580
rect 12894 26528 12900 26580
rect 12952 26568 12958 26580
rect 16117 26571 16175 26577
rect 16117 26568 16129 26571
rect 12952 26540 16129 26568
rect 12952 26528 12958 26540
rect 16117 26537 16129 26540
rect 16163 26537 16175 26571
rect 16117 26531 16175 26537
rect 16942 26528 16948 26580
rect 17000 26568 17006 26580
rect 17681 26571 17739 26577
rect 17681 26568 17693 26571
rect 17000 26540 17693 26568
rect 17000 26528 17006 26540
rect 17681 26537 17693 26540
rect 17727 26537 17739 26571
rect 17681 26531 17739 26537
rect 18138 26528 18144 26580
rect 18196 26528 18202 26580
rect 21082 26528 21088 26580
rect 21140 26568 21146 26580
rect 22189 26571 22247 26577
rect 22189 26568 22201 26571
rect 21140 26540 22201 26568
rect 21140 26528 21146 26540
rect 22189 26537 22201 26540
rect 22235 26568 22247 26571
rect 22370 26568 22376 26580
rect 22235 26540 22376 26568
rect 22235 26537 22247 26540
rect 22189 26531 22247 26537
rect 22370 26528 22376 26540
rect 22428 26528 22434 26580
rect 22922 26528 22928 26580
rect 22980 26568 22986 26580
rect 24946 26568 24952 26580
rect 22980 26540 24952 26568
rect 22980 26528 22986 26540
rect 24946 26528 24952 26540
rect 25004 26528 25010 26580
rect 25866 26528 25872 26580
rect 25924 26568 25930 26580
rect 26513 26571 26571 26577
rect 26513 26568 26525 26571
rect 25924 26540 26525 26568
rect 25924 26528 25930 26540
rect 26513 26537 26525 26540
rect 26559 26537 26571 26571
rect 26513 26531 26571 26537
rect 4430 26500 4436 26512
rect 2746 26472 4436 26500
rect 4430 26460 4436 26472
rect 4488 26460 4494 26512
rect 4798 26460 4804 26512
rect 4856 26500 4862 26512
rect 5905 26503 5963 26509
rect 5905 26500 5917 26503
rect 4856 26472 5917 26500
rect 4856 26460 4862 26472
rect 5905 26469 5917 26472
rect 5951 26469 5963 26503
rect 7484 26500 7512 26528
rect 8386 26500 8392 26512
rect 7484 26472 8392 26500
rect 5905 26463 5963 26469
rect 8386 26460 8392 26472
rect 8444 26500 8450 26512
rect 13265 26503 13323 26509
rect 8444 26472 12434 26500
rect 8444 26460 8450 26472
rect 1397 26435 1455 26441
rect 1397 26401 1409 26435
rect 1443 26432 1455 26435
rect 2866 26432 2872 26444
rect 1443 26404 2872 26432
rect 1443 26401 1455 26404
rect 1397 26395 1455 26401
rect 2866 26392 2872 26404
rect 2924 26392 2930 26444
rect 2958 26392 2964 26444
rect 3016 26432 3022 26444
rect 3145 26435 3203 26441
rect 3145 26432 3157 26435
rect 3016 26404 3157 26432
rect 3016 26392 3022 26404
rect 3145 26401 3157 26404
rect 3191 26432 3203 26435
rect 3878 26432 3884 26444
rect 3191 26404 3884 26432
rect 3191 26401 3203 26404
rect 3145 26395 3203 26401
rect 3878 26392 3884 26404
rect 3936 26392 3942 26444
rect 4062 26392 4068 26444
rect 4120 26432 4126 26444
rect 4249 26435 4307 26441
rect 4249 26432 4261 26435
rect 4120 26404 4261 26432
rect 4120 26392 4126 26404
rect 4249 26401 4261 26404
rect 4295 26401 4307 26435
rect 4249 26395 4307 26401
rect 4338 26392 4344 26444
rect 4396 26392 4402 26444
rect 5537 26435 5595 26441
rect 5537 26401 5549 26435
rect 5583 26432 5595 26435
rect 5718 26432 5724 26444
rect 5583 26404 5724 26432
rect 5583 26401 5595 26404
rect 5537 26395 5595 26401
rect 5718 26392 5724 26404
rect 5776 26392 5782 26444
rect 7190 26432 7196 26444
rect 5828 26404 7196 26432
rect 2774 26324 2780 26376
rect 2832 26324 2838 26376
rect 4157 26367 4215 26373
rect 4157 26333 4169 26367
rect 4203 26364 4215 26367
rect 4614 26364 4620 26376
rect 4203 26336 4620 26364
rect 4203 26333 4215 26336
rect 4157 26327 4215 26333
rect 4614 26324 4620 26336
rect 4672 26324 4678 26376
rect 4709 26367 4767 26373
rect 4709 26333 4721 26367
rect 4755 26364 4767 26367
rect 4982 26364 4988 26376
rect 4755 26336 4988 26364
rect 4755 26333 4767 26336
rect 4709 26327 4767 26333
rect 4982 26324 4988 26336
rect 5040 26364 5046 26376
rect 5828 26373 5856 26404
rect 7190 26392 7196 26404
rect 7248 26392 7254 26444
rect 7469 26435 7527 26441
rect 7469 26432 7481 26435
rect 7300 26404 7481 26432
rect 5813 26367 5871 26373
rect 5813 26364 5825 26367
rect 5040 26336 5825 26364
rect 5040 26324 5046 26336
rect 5813 26333 5825 26336
rect 5859 26333 5871 26367
rect 5813 26327 5871 26333
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26333 6239 26367
rect 6181 26327 6239 26333
rect 5077 26299 5135 26305
rect 5077 26265 5089 26299
rect 5123 26296 5135 26299
rect 6086 26296 6092 26308
rect 5123 26268 6092 26296
rect 5123 26265 5135 26268
rect 5077 26259 5135 26265
rect 6086 26256 6092 26268
rect 6144 26256 6150 26308
rect 6196 26296 6224 26327
rect 6270 26324 6276 26376
rect 6328 26324 6334 26376
rect 6546 26296 6552 26308
rect 6196 26268 6552 26296
rect 6546 26256 6552 26268
rect 6604 26296 6610 26308
rect 7300 26296 7328 26404
rect 7469 26401 7481 26404
rect 7515 26432 7527 26435
rect 9030 26432 9036 26444
rect 7515 26404 9036 26432
rect 7515 26401 7527 26404
rect 7469 26395 7527 26401
rect 9030 26392 9036 26404
rect 9088 26392 9094 26444
rect 10318 26392 10324 26444
rect 10376 26432 10382 26444
rect 11974 26432 11980 26444
rect 10376 26404 11980 26432
rect 10376 26392 10382 26404
rect 7377 26367 7435 26373
rect 7377 26333 7389 26367
rect 7423 26333 7435 26367
rect 7377 26327 7435 26333
rect 6604 26268 7328 26296
rect 7392 26296 7420 26327
rect 9582 26324 9588 26376
rect 9640 26364 9646 26376
rect 11057 26367 11115 26373
rect 11057 26364 11069 26367
rect 9640 26336 11069 26364
rect 9640 26324 9646 26336
rect 11057 26333 11069 26336
rect 11103 26333 11115 26367
rect 11057 26327 11115 26333
rect 11241 26367 11299 26373
rect 11241 26333 11253 26367
rect 11287 26364 11299 26367
rect 11330 26364 11336 26376
rect 11287 26336 11336 26364
rect 11287 26333 11299 26336
rect 11241 26327 11299 26333
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 11624 26373 11652 26404
rect 11974 26392 11980 26404
rect 12032 26392 12038 26444
rect 11425 26367 11483 26373
rect 11425 26333 11437 26367
rect 11471 26333 11483 26367
rect 11425 26327 11483 26333
rect 11609 26367 11667 26373
rect 11609 26333 11621 26367
rect 11655 26333 11667 26367
rect 11609 26327 11667 26333
rect 8110 26296 8116 26308
rect 7392 26268 8116 26296
rect 6604 26256 6610 26268
rect 8110 26256 8116 26268
rect 8168 26256 8174 26308
rect 11440 26296 11468 26327
rect 12158 26296 12164 26308
rect 9416 26268 11284 26296
rect 11440 26268 12164 26296
rect 2682 26188 2688 26240
rect 2740 26228 2746 26240
rect 4706 26228 4712 26240
rect 2740 26200 4712 26228
rect 2740 26188 2746 26200
rect 4706 26188 4712 26200
rect 4764 26188 4770 26240
rect 5350 26188 5356 26240
rect 5408 26228 5414 26240
rect 9416 26228 9444 26268
rect 11256 26240 11284 26268
rect 12158 26256 12164 26268
rect 12216 26256 12222 26308
rect 12406 26296 12434 26472
rect 13265 26469 13277 26503
rect 13311 26500 13323 26503
rect 13630 26500 13636 26512
rect 13311 26472 13636 26500
rect 13311 26469 13323 26472
rect 13265 26463 13323 26469
rect 13630 26460 13636 26472
rect 13688 26460 13694 26512
rect 15194 26460 15200 26512
rect 15252 26460 15258 26512
rect 17034 26460 17040 26512
rect 17092 26500 17098 26512
rect 17218 26500 17224 26512
rect 17092 26472 17224 26500
rect 17092 26460 17098 26472
rect 17218 26460 17224 26472
rect 17276 26460 17282 26512
rect 20254 26460 20260 26512
rect 20312 26460 20318 26512
rect 23290 26500 23296 26512
rect 20732 26472 23296 26500
rect 13354 26392 13360 26444
rect 13412 26392 13418 26444
rect 15212 26432 15240 26460
rect 14476 26404 15240 26432
rect 16485 26435 16543 26441
rect 12526 26324 12532 26376
rect 12584 26364 12590 26376
rect 12621 26367 12679 26373
rect 12621 26364 12633 26367
rect 12584 26336 12633 26364
rect 12584 26324 12590 26336
rect 12621 26333 12633 26336
rect 12667 26333 12679 26367
rect 12621 26327 12679 26333
rect 12714 26367 12772 26373
rect 12714 26333 12726 26367
rect 12760 26333 12772 26367
rect 12714 26327 12772 26333
rect 12728 26296 12756 26327
rect 12802 26324 12808 26376
rect 12860 26364 12866 26376
rect 13086 26367 13144 26373
rect 13086 26364 13098 26367
rect 12860 26336 13098 26364
rect 12860 26324 12866 26336
rect 13086 26333 13098 26336
rect 13132 26333 13144 26367
rect 13086 26327 13144 26333
rect 13541 26367 13599 26373
rect 13541 26333 13553 26367
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 12406 26268 12756 26296
rect 12894 26256 12900 26308
rect 12952 26256 12958 26308
rect 12986 26256 12992 26308
rect 13044 26256 13050 26308
rect 13556 26296 13584 26327
rect 13722 26324 13728 26376
rect 13780 26324 13786 26376
rect 14476 26373 14504 26404
rect 16485 26401 16497 26435
rect 16531 26432 16543 26435
rect 18138 26432 18144 26444
rect 16531 26404 18144 26432
rect 16531 26401 16543 26404
rect 16485 26395 16543 26401
rect 18138 26392 18144 26404
rect 18196 26392 18202 26444
rect 18506 26392 18512 26444
rect 18564 26432 18570 26444
rect 20732 26432 20760 26472
rect 23290 26460 23296 26472
rect 23348 26460 23354 26512
rect 23382 26460 23388 26512
rect 23440 26500 23446 26512
rect 23477 26503 23535 26509
rect 23477 26500 23489 26503
rect 23440 26472 23489 26500
rect 23440 26460 23446 26472
rect 23477 26469 23489 26472
rect 23523 26469 23535 26503
rect 23477 26463 23535 26469
rect 25590 26460 25596 26512
rect 25648 26500 25654 26512
rect 26528 26500 26556 26531
rect 26694 26528 26700 26580
rect 26752 26568 26758 26580
rect 28810 26568 28816 26580
rect 26752 26540 28816 26568
rect 26752 26528 26758 26540
rect 28810 26528 28816 26540
rect 28868 26528 28874 26580
rect 31570 26568 31576 26580
rect 29840 26540 31576 26568
rect 25648 26472 26004 26500
rect 26528 26472 27384 26500
rect 25648 26460 25654 26472
rect 18564 26404 20760 26432
rect 20809 26435 20867 26441
rect 18564 26392 18570 26404
rect 20809 26401 20821 26435
rect 20855 26432 20867 26435
rect 22094 26432 22100 26444
rect 20855 26404 22100 26432
rect 20855 26401 20867 26404
rect 20809 26395 20867 26401
rect 22094 26392 22100 26404
rect 22152 26432 22158 26444
rect 25038 26432 25044 26444
rect 22152 26404 25044 26432
rect 22152 26392 22158 26404
rect 25038 26392 25044 26404
rect 25096 26392 25102 26444
rect 25501 26435 25559 26441
rect 25501 26401 25513 26435
rect 25547 26432 25559 26435
rect 25774 26432 25780 26444
rect 25547 26404 25780 26432
rect 25547 26401 25559 26404
rect 25501 26395 25559 26401
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26333 14519 26367
rect 14461 26327 14519 26333
rect 15013 26367 15071 26373
rect 15013 26333 15025 26367
rect 15059 26333 15071 26367
rect 15013 26327 15071 26333
rect 15197 26367 15255 26373
rect 15197 26333 15209 26367
rect 15243 26333 15255 26367
rect 15197 26327 15255 26333
rect 13814 26296 13820 26308
rect 13556 26268 13820 26296
rect 13814 26256 13820 26268
rect 13872 26256 13878 26308
rect 14090 26256 14096 26308
rect 14148 26296 14154 26308
rect 14292 26296 14320 26327
rect 14829 26299 14887 26305
rect 14829 26296 14841 26299
rect 14148 26268 14841 26296
rect 14148 26256 14154 26268
rect 14829 26265 14841 26268
rect 14875 26265 14887 26299
rect 14829 26259 14887 26265
rect 5408 26200 9444 26228
rect 5408 26188 5414 26200
rect 9490 26188 9496 26240
rect 9548 26228 9554 26240
rect 10594 26228 10600 26240
rect 9548 26200 10600 26228
rect 9548 26188 9554 26200
rect 10594 26188 10600 26200
rect 10652 26188 10658 26240
rect 10686 26188 10692 26240
rect 10744 26228 10750 26240
rect 10962 26228 10968 26240
rect 10744 26200 10968 26228
rect 10744 26188 10750 26200
rect 10962 26188 10968 26200
rect 11020 26188 11026 26240
rect 11238 26188 11244 26240
rect 11296 26188 11302 26240
rect 11330 26188 11336 26240
rect 11388 26228 11394 26240
rect 11790 26228 11796 26240
rect 11388 26200 11796 26228
rect 11388 26188 11394 26200
rect 11790 26188 11796 26200
rect 11848 26228 11854 26240
rect 12710 26228 12716 26240
rect 11848 26200 12716 26228
rect 11848 26188 11854 26200
rect 12710 26188 12716 26200
rect 12768 26228 12774 26240
rect 12912 26228 12940 26256
rect 12768 26200 12940 26228
rect 12768 26188 12774 26200
rect 13446 26188 13452 26240
rect 13504 26228 13510 26240
rect 14185 26231 14243 26237
rect 14185 26228 14197 26231
rect 13504 26200 14197 26228
rect 13504 26188 13510 26200
rect 14185 26197 14197 26200
rect 14231 26197 14243 26231
rect 15028 26228 15056 26327
rect 15212 26296 15240 26327
rect 15838 26324 15844 26376
rect 15896 26324 15902 26376
rect 16022 26364 16028 26376
rect 15948 26336 16028 26364
rect 15948 26296 15976 26336
rect 16022 26324 16028 26336
rect 16080 26324 16086 26376
rect 16393 26367 16451 26373
rect 16393 26333 16405 26367
rect 16439 26333 16451 26367
rect 16393 26327 16451 26333
rect 16408 26296 16436 26327
rect 16942 26324 16948 26376
rect 17000 26324 17006 26376
rect 18049 26367 18107 26373
rect 18049 26364 18061 26367
rect 17052 26336 18061 26364
rect 17052 26296 17080 26336
rect 18049 26333 18061 26336
rect 18095 26333 18107 26367
rect 18049 26327 18107 26333
rect 18233 26367 18291 26373
rect 18233 26333 18245 26367
rect 18279 26364 18291 26367
rect 18598 26364 18604 26376
rect 18279 26336 18604 26364
rect 18279 26333 18291 26336
rect 18233 26327 18291 26333
rect 18598 26324 18604 26336
rect 18656 26324 18662 26376
rect 20346 26324 20352 26376
rect 20404 26324 20410 26376
rect 20625 26367 20683 26373
rect 20625 26333 20637 26367
rect 20671 26364 20683 26367
rect 22922 26364 22928 26376
rect 20671 26336 22928 26364
rect 20671 26333 20683 26336
rect 20625 26327 20683 26333
rect 15212 26268 15976 26296
rect 16040 26268 16436 26296
rect 16592 26268 17080 26296
rect 16040 26240 16068 26268
rect 15838 26228 15844 26240
rect 15028 26200 15844 26228
rect 14185 26191 14243 26197
rect 15838 26188 15844 26200
rect 15896 26188 15902 26240
rect 16022 26188 16028 26240
rect 16080 26188 16086 26240
rect 16390 26188 16396 26240
rect 16448 26228 16454 26240
rect 16592 26228 16620 26268
rect 17310 26256 17316 26308
rect 17368 26256 17374 26308
rect 17494 26256 17500 26308
rect 17552 26256 17558 26308
rect 19242 26256 19248 26308
rect 19300 26296 19306 26308
rect 19978 26296 19984 26308
rect 19300 26268 19984 26296
rect 19300 26256 19306 26268
rect 19978 26256 19984 26268
rect 20036 26256 20042 26308
rect 20254 26256 20260 26308
rect 20312 26296 20318 26308
rect 20640 26296 20668 26327
rect 22922 26324 22928 26336
rect 22980 26324 22986 26376
rect 23106 26364 23112 26376
rect 23032 26336 23112 26364
rect 20312 26268 20668 26296
rect 20312 26256 20318 26268
rect 20714 26256 20720 26308
rect 20772 26296 20778 26308
rect 21358 26296 21364 26308
rect 20772 26268 21364 26296
rect 20772 26256 20778 26268
rect 21358 26256 21364 26268
rect 21416 26256 21422 26308
rect 21818 26296 21824 26308
rect 21560 26268 21824 26296
rect 16448 26200 16620 26228
rect 16448 26188 16454 26200
rect 16758 26188 16764 26240
rect 16816 26228 16822 26240
rect 19426 26228 19432 26240
rect 16816 26200 19432 26228
rect 16816 26188 16822 26200
rect 19426 26188 19432 26200
rect 19484 26188 19490 26240
rect 19610 26188 19616 26240
rect 19668 26228 19674 26240
rect 21560 26228 21588 26268
rect 21818 26256 21824 26268
rect 21876 26256 21882 26308
rect 21910 26256 21916 26308
rect 21968 26256 21974 26308
rect 22002 26256 22008 26308
rect 22060 26296 22066 26308
rect 22738 26296 22744 26308
rect 22060 26268 22744 26296
rect 22060 26256 22066 26268
rect 22738 26256 22744 26268
rect 22796 26296 22802 26308
rect 23032 26296 23060 26336
rect 23106 26324 23112 26336
rect 23164 26364 23170 26376
rect 23293 26367 23351 26373
rect 23293 26364 23305 26367
rect 23164 26336 23305 26364
rect 23164 26324 23170 26336
rect 23293 26333 23305 26336
rect 23339 26333 23351 26367
rect 23293 26327 23351 26333
rect 25406 26324 25412 26376
rect 25464 26324 25470 26376
rect 25700 26373 25728 26404
rect 25774 26392 25780 26404
rect 25832 26392 25838 26444
rect 25976 26432 26004 26472
rect 26602 26432 26608 26444
rect 25976 26404 26608 26432
rect 25593 26367 25651 26373
rect 25593 26333 25605 26367
rect 25639 26333 25651 26367
rect 25593 26327 25651 26333
rect 25685 26367 25743 26373
rect 25685 26333 25697 26367
rect 25731 26333 25743 26367
rect 25685 26327 25743 26333
rect 22796 26268 23060 26296
rect 25608 26296 25636 26327
rect 25866 26324 25872 26376
rect 25924 26324 25930 26376
rect 25976 26373 26004 26404
rect 26602 26392 26608 26404
rect 26660 26392 26666 26444
rect 26970 26392 26976 26444
rect 27028 26432 27034 26444
rect 27028 26404 27200 26432
rect 27028 26392 27034 26404
rect 25961 26367 26019 26373
rect 25961 26333 25973 26367
rect 26007 26333 26019 26367
rect 25961 26327 26019 26333
rect 26234 26324 26240 26376
rect 26292 26324 26298 26376
rect 26694 26324 26700 26376
rect 26752 26324 26758 26376
rect 27065 26367 27123 26373
rect 27065 26333 27077 26367
rect 27111 26333 27123 26367
rect 27172 26364 27200 26404
rect 27356 26373 27384 26472
rect 27448 26404 28120 26432
rect 27448 26376 27476 26404
rect 27249 26367 27307 26373
rect 27249 26364 27261 26367
rect 27172 26336 27261 26364
rect 27065 26327 27123 26333
rect 27249 26333 27261 26336
rect 27295 26333 27307 26367
rect 27249 26327 27307 26333
rect 27341 26367 27399 26373
rect 27341 26333 27353 26367
rect 27387 26333 27399 26367
rect 27341 26327 27399 26333
rect 25608 26268 25728 26296
rect 22796 26256 22802 26268
rect 19668 26200 21588 26228
rect 19668 26188 19674 26200
rect 21634 26188 21640 26240
rect 21692 26228 21698 26240
rect 23658 26228 23664 26240
rect 21692 26200 23664 26228
rect 21692 26188 21698 26200
rect 23658 26188 23664 26200
rect 23716 26188 23722 26240
rect 25700 26228 25728 26268
rect 25774 26256 25780 26308
rect 25832 26256 25838 26308
rect 26970 26296 26976 26308
rect 25884 26268 26976 26296
rect 25884 26228 25912 26268
rect 26970 26256 26976 26268
rect 27028 26296 27034 26308
rect 27080 26296 27108 26327
rect 27430 26324 27436 26376
rect 27488 26324 27494 26376
rect 27525 26367 27583 26373
rect 27525 26333 27537 26367
rect 27571 26333 27583 26367
rect 27525 26327 27583 26333
rect 27028 26268 27108 26296
rect 27157 26299 27215 26305
rect 27028 26256 27034 26268
rect 27157 26265 27169 26299
rect 27203 26296 27215 26299
rect 27540 26296 27568 26327
rect 27706 26324 27712 26376
rect 27764 26324 27770 26376
rect 27890 26373 27896 26376
rect 27857 26367 27896 26373
rect 27857 26333 27869 26367
rect 27857 26327 27896 26333
rect 27890 26324 27896 26327
rect 27948 26324 27954 26376
rect 27982 26324 27988 26376
rect 28040 26324 28046 26376
rect 28092 26373 28120 26404
rect 28077 26367 28135 26373
rect 28077 26333 28089 26367
rect 28123 26333 28135 26367
rect 28077 26327 28135 26333
rect 28215 26367 28273 26373
rect 28215 26333 28227 26367
rect 28261 26364 28273 26367
rect 28442 26364 28448 26376
rect 28261 26336 28448 26364
rect 28261 26333 28273 26336
rect 28215 26327 28273 26333
rect 28442 26324 28448 26336
rect 28500 26324 28506 26376
rect 29454 26324 29460 26376
rect 29512 26364 29518 26376
rect 29549 26367 29607 26373
rect 29549 26364 29561 26367
rect 29512 26336 29561 26364
rect 29512 26324 29518 26336
rect 29549 26333 29561 26336
rect 29595 26333 29607 26367
rect 29549 26327 29607 26333
rect 29638 26324 29644 26376
rect 29696 26324 29702 26376
rect 29840 26373 29868 26540
rect 31570 26528 31576 26540
rect 31628 26528 31634 26580
rect 31665 26571 31723 26577
rect 31665 26537 31677 26571
rect 31711 26568 31723 26571
rect 31754 26568 31760 26580
rect 31711 26540 31760 26568
rect 31711 26537 31723 26540
rect 31665 26531 31723 26537
rect 31754 26528 31760 26540
rect 31812 26528 31818 26580
rect 31941 26571 31999 26577
rect 31941 26537 31953 26571
rect 31987 26568 31999 26571
rect 32122 26568 32128 26580
rect 31987 26540 32128 26568
rect 31987 26537 31999 26540
rect 31941 26531 31999 26537
rect 32122 26528 32128 26540
rect 32180 26528 32186 26580
rect 32217 26571 32275 26577
rect 32217 26537 32229 26571
rect 32263 26537 32275 26571
rect 32217 26531 32275 26537
rect 30374 26460 30380 26512
rect 30432 26500 30438 26512
rect 30926 26500 30932 26512
rect 30432 26472 30932 26500
rect 30432 26460 30438 26472
rect 30926 26460 30932 26472
rect 30984 26500 30990 26512
rect 32232 26500 32260 26531
rect 30984 26472 32260 26500
rect 30984 26460 30990 26472
rect 31665 26435 31723 26441
rect 31665 26401 31677 26435
rect 31711 26432 31723 26435
rect 32122 26432 32128 26444
rect 31711 26404 32128 26432
rect 31711 26401 31723 26404
rect 31665 26395 31723 26401
rect 32122 26392 32128 26404
rect 32180 26392 32186 26444
rect 32398 26392 32404 26444
rect 32456 26432 32462 26444
rect 32674 26432 32680 26444
rect 32456 26404 32680 26432
rect 32456 26392 32462 26404
rect 32674 26392 32680 26404
rect 32732 26392 32738 26444
rect 29825 26367 29883 26373
rect 29825 26333 29837 26367
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 29914 26324 29920 26376
rect 29972 26324 29978 26376
rect 30101 26367 30159 26373
rect 30101 26333 30113 26367
rect 30147 26364 30159 26367
rect 31757 26367 31815 26373
rect 30147 26336 31616 26364
rect 30147 26333 30159 26336
rect 30101 26327 30159 26333
rect 27614 26296 27620 26308
rect 27203 26268 27620 26296
rect 27203 26265 27215 26268
rect 27157 26259 27215 26265
rect 27614 26256 27620 26268
rect 27672 26256 27678 26308
rect 31481 26299 31539 26305
rect 31481 26296 31493 26299
rect 28368 26268 31493 26296
rect 25700 26200 25912 26228
rect 26237 26231 26295 26237
rect 26237 26197 26249 26231
rect 26283 26228 26295 26231
rect 26418 26228 26424 26240
rect 26283 26200 26424 26228
rect 26283 26197 26295 26200
rect 26237 26191 26295 26197
rect 26418 26188 26424 26200
rect 26476 26188 26482 26240
rect 26786 26188 26792 26240
rect 26844 26228 26850 26240
rect 27246 26228 27252 26240
rect 26844 26200 27252 26228
rect 26844 26188 26850 26200
rect 27246 26188 27252 26200
rect 27304 26188 27310 26240
rect 28368 26237 28396 26268
rect 31481 26265 31493 26268
rect 31527 26265 31539 26299
rect 31588 26296 31616 26336
rect 31757 26333 31769 26367
rect 31803 26364 31815 26367
rect 31846 26364 31852 26376
rect 31803 26336 31852 26364
rect 31803 26333 31815 26336
rect 31757 26327 31815 26333
rect 31846 26324 31852 26336
rect 31904 26324 31910 26376
rect 33962 26364 33968 26376
rect 31956 26336 33968 26364
rect 31956 26296 31984 26336
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 34057 26367 34115 26373
rect 34057 26333 34069 26367
rect 34103 26333 34115 26367
rect 34057 26327 34115 26333
rect 31588 26268 31984 26296
rect 31481 26259 31539 26265
rect 32030 26256 32036 26308
rect 32088 26256 32094 26308
rect 32233 26299 32291 26305
rect 32233 26296 32245 26299
rect 32140 26268 32245 26296
rect 28353 26231 28411 26237
rect 28353 26197 28365 26231
rect 28399 26197 28411 26231
rect 28353 26191 28411 26197
rect 31938 26188 31944 26240
rect 31996 26228 32002 26240
rect 32140 26228 32168 26268
rect 32233 26265 32245 26268
rect 32279 26265 32291 26299
rect 32233 26259 32291 26265
rect 33134 26256 33140 26308
rect 33192 26296 33198 26308
rect 33318 26296 33324 26308
rect 33192 26268 33324 26296
rect 33192 26256 33198 26268
rect 33318 26256 33324 26268
rect 33376 26296 33382 26308
rect 34072 26296 34100 26327
rect 34146 26324 34152 26376
rect 34204 26324 34210 26376
rect 33376 26268 34100 26296
rect 33376 26256 33382 26268
rect 31996 26200 32168 26228
rect 31996 26188 32002 26200
rect 32398 26188 32404 26240
rect 32456 26188 32462 26240
rect 33778 26188 33784 26240
rect 33836 26228 33842 26240
rect 33873 26231 33931 26237
rect 33873 26228 33885 26231
rect 33836 26200 33885 26228
rect 33836 26188 33842 26200
rect 33873 26197 33885 26200
rect 33919 26197 33931 26231
rect 33873 26191 33931 26197
rect 1104 26138 36432 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 36432 26138
rect 1104 26064 36432 26086
rect 2130 25984 2136 26036
rect 2188 25984 2194 26036
rect 3050 25984 3056 26036
rect 3108 26024 3114 26036
rect 4338 26024 4344 26036
rect 3108 25996 4344 26024
rect 3108 25984 3114 25996
rect 4338 25984 4344 25996
rect 4396 25984 4402 26036
rect 4430 25984 4436 26036
rect 4488 25984 4494 26036
rect 4706 25984 4712 26036
rect 4764 26024 4770 26036
rect 4801 26027 4859 26033
rect 4801 26024 4813 26027
rect 4764 25996 4813 26024
rect 4764 25984 4770 25996
rect 4801 25993 4813 25996
rect 4847 26024 4859 26027
rect 5258 26024 5264 26036
rect 4847 25996 5264 26024
rect 4847 25993 4859 25996
rect 4801 25987 4859 25993
rect 5258 25984 5264 25996
rect 5316 25984 5322 26036
rect 6086 25984 6092 26036
rect 6144 25984 6150 26036
rect 6196 25996 9628 26024
rect 3068 25956 3096 25984
rect 2424 25928 3096 25956
rect 2225 25823 2283 25829
rect 2225 25789 2237 25823
rect 2271 25820 2283 25823
rect 2314 25820 2320 25832
rect 2271 25792 2320 25820
rect 2271 25789 2283 25792
rect 2225 25783 2283 25789
rect 2314 25780 2320 25792
rect 2372 25780 2378 25832
rect 2424 25829 2452 25928
rect 4614 25916 4620 25968
rect 4672 25956 4678 25968
rect 6196 25956 6224 25996
rect 4672 25928 6224 25956
rect 7285 25959 7343 25965
rect 4672 25916 4678 25928
rect 7285 25925 7297 25959
rect 7331 25956 7343 25959
rect 7374 25956 7380 25968
rect 7331 25928 7380 25956
rect 7331 25925 7343 25928
rect 7285 25919 7343 25925
rect 7374 25916 7380 25928
rect 7432 25916 7438 25968
rect 7469 25959 7527 25965
rect 7469 25925 7481 25959
rect 7515 25956 7527 25959
rect 7834 25956 7840 25968
rect 7515 25928 7840 25956
rect 7515 25925 7527 25928
rect 7469 25919 7527 25925
rect 7834 25916 7840 25928
rect 7892 25916 7898 25968
rect 9125 25959 9183 25965
rect 8772 25928 8984 25956
rect 3970 25848 3976 25900
rect 4028 25848 4034 25900
rect 4338 25848 4344 25900
rect 4396 25888 4402 25900
rect 5997 25891 6055 25897
rect 4396 25860 5120 25888
rect 4396 25848 4402 25860
rect 2409 25823 2467 25829
rect 2409 25789 2421 25823
rect 2455 25789 2467 25823
rect 2409 25783 2467 25789
rect 2593 25823 2651 25829
rect 2593 25789 2605 25823
rect 2639 25789 2651 25823
rect 2593 25783 2651 25789
rect 2869 25823 2927 25829
rect 2869 25789 2881 25823
rect 2915 25820 2927 25823
rect 4706 25820 4712 25832
rect 2915 25792 4712 25820
rect 2915 25789 2927 25792
rect 2869 25783 2927 25789
rect 1670 25644 1676 25696
rect 1728 25684 1734 25696
rect 1765 25687 1823 25693
rect 1765 25684 1777 25687
rect 1728 25656 1777 25684
rect 1728 25644 1734 25656
rect 1765 25653 1777 25656
rect 1811 25653 1823 25687
rect 2608 25684 2636 25783
rect 4706 25780 4712 25792
rect 4764 25780 4770 25832
rect 4893 25823 4951 25829
rect 4893 25820 4905 25823
rect 4816 25792 4905 25820
rect 3878 25712 3884 25764
rect 3936 25752 3942 25764
rect 4816 25752 4844 25792
rect 4893 25789 4905 25792
rect 4939 25820 4951 25823
rect 4982 25820 4988 25832
rect 4939 25792 4988 25820
rect 4939 25789 4951 25792
rect 4893 25783 4951 25789
rect 4982 25780 4988 25792
rect 5040 25780 5046 25832
rect 5092 25829 5120 25860
rect 5997 25857 6009 25891
rect 6043 25857 6055 25891
rect 5997 25851 6055 25857
rect 6181 25891 6239 25897
rect 6181 25857 6193 25891
rect 6227 25888 6239 25891
rect 6546 25888 6552 25900
rect 6227 25860 6552 25888
rect 6227 25857 6239 25860
rect 6181 25851 6239 25857
rect 5077 25823 5135 25829
rect 5077 25789 5089 25823
rect 5123 25820 5135 25823
rect 5534 25820 5540 25832
rect 5123 25792 5540 25820
rect 5123 25789 5135 25792
rect 5077 25783 5135 25789
rect 5534 25780 5540 25792
rect 5592 25780 5598 25832
rect 5813 25823 5871 25829
rect 5813 25789 5825 25823
rect 5859 25789 5871 25823
rect 6012 25820 6040 25851
rect 6546 25848 6552 25860
rect 6604 25848 6610 25900
rect 7190 25848 7196 25900
rect 7248 25888 7254 25900
rect 7561 25891 7619 25897
rect 7561 25888 7573 25891
rect 7248 25860 7573 25888
rect 7248 25848 7254 25860
rect 7561 25857 7573 25860
rect 7607 25857 7619 25891
rect 7561 25851 7619 25857
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25888 7987 25891
rect 8478 25888 8484 25900
rect 7975 25860 8484 25888
rect 7975 25857 7987 25860
rect 7929 25851 7987 25857
rect 8478 25848 8484 25860
rect 8536 25848 8542 25900
rect 8772 25897 8800 25928
rect 8757 25891 8815 25897
rect 8757 25857 8769 25891
rect 8803 25857 8815 25891
rect 8757 25851 8815 25857
rect 8850 25891 8908 25897
rect 8850 25857 8862 25891
rect 8896 25857 8908 25891
rect 8850 25851 8908 25857
rect 6730 25820 6736 25832
rect 6012 25792 6736 25820
rect 5813 25783 5871 25789
rect 5828 25752 5856 25783
rect 6730 25780 6736 25792
rect 6788 25780 6794 25832
rect 8864 25752 8892 25851
rect 3936 25724 4844 25752
rect 5184 25724 8892 25752
rect 3936 25712 3942 25724
rect 2866 25684 2872 25696
rect 2608 25656 2872 25684
rect 1765 25647 1823 25653
rect 2866 25644 2872 25656
rect 2924 25644 2930 25696
rect 3418 25644 3424 25696
rect 3476 25684 3482 25696
rect 4341 25687 4399 25693
rect 4341 25684 4353 25687
rect 3476 25656 4353 25684
rect 3476 25644 3482 25656
rect 4341 25653 4353 25656
rect 4387 25684 4399 25687
rect 5184 25684 5212 25724
rect 4387 25656 5212 25684
rect 4387 25653 4399 25656
rect 4341 25647 4399 25653
rect 5258 25644 5264 25696
rect 5316 25644 5322 25696
rect 5350 25644 5356 25696
rect 5408 25684 5414 25696
rect 7009 25687 7067 25693
rect 7009 25684 7021 25687
rect 5408 25656 7021 25684
rect 5408 25644 5414 25656
rect 7009 25653 7021 25656
rect 7055 25653 7067 25687
rect 7009 25647 7067 25653
rect 7834 25644 7840 25696
rect 7892 25644 7898 25696
rect 8956 25684 8984 25928
rect 9125 25925 9137 25959
rect 9171 25956 9183 25959
rect 9398 25956 9404 25968
rect 9171 25928 9404 25956
rect 9171 25925 9183 25928
rect 9125 25919 9183 25925
rect 9398 25916 9404 25928
rect 9456 25916 9462 25968
rect 9033 25891 9091 25897
rect 9033 25857 9045 25891
rect 9079 25857 9091 25891
rect 9033 25851 9091 25857
rect 9263 25891 9321 25897
rect 9263 25857 9275 25891
rect 9309 25888 9321 25891
rect 9309 25860 9444 25888
rect 9309 25857 9321 25860
rect 9263 25851 9321 25857
rect 9048 25752 9076 25851
rect 9416 25820 9444 25860
rect 9490 25848 9496 25900
rect 9548 25848 9554 25900
rect 9600 25897 9628 25996
rect 9784 25996 11100 26024
rect 9784 25968 9812 25996
rect 9766 25916 9772 25968
rect 9824 25916 9830 25968
rect 9861 25959 9919 25965
rect 9861 25925 9873 25959
rect 9907 25956 9919 25959
rect 10134 25956 10140 25968
rect 9907 25928 10140 25956
rect 9907 25925 9919 25928
rect 9861 25919 9919 25925
rect 10134 25916 10140 25928
rect 10192 25916 10198 25968
rect 10888 25965 10916 25996
rect 10873 25959 10931 25965
rect 10873 25925 10885 25959
rect 10919 25925 10931 25959
rect 10873 25919 10931 25925
rect 10962 25916 10968 25968
rect 11020 25916 11026 25968
rect 11072 25956 11100 25996
rect 11238 25984 11244 26036
rect 11296 26024 11302 26036
rect 11296 25996 12481 26024
rect 11296 25984 11302 25996
rect 11330 25956 11336 25968
rect 11072 25928 11336 25956
rect 11330 25916 11336 25928
rect 11388 25916 11394 25968
rect 11514 25916 11520 25968
rect 11572 25956 11578 25968
rect 11572 25928 11928 25956
rect 11572 25916 11578 25928
rect 9586 25891 9644 25897
rect 9586 25857 9598 25891
rect 9632 25857 9644 25891
rect 9586 25851 9644 25857
rect 9958 25891 10016 25897
rect 9958 25857 9970 25891
rect 10004 25857 10016 25891
rect 9958 25851 10016 25857
rect 9968 25820 9996 25851
rect 10594 25848 10600 25900
rect 10652 25848 10658 25900
rect 10689 25891 10747 25897
rect 10689 25857 10701 25891
rect 10735 25888 10747 25891
rect 10778 25888 10784 25900
rect 10735 25860 10784 25888
rect 10735 25857 10747 25860
rect 10689 25851 10747 25857
rect 10778 25848 10784 25860
rect 10836 25848 10842 25900
rect 11054 25848 11060 25900
rect 11112 25848 11118 25900
rect 11900 25897 11928 25928
rect 12453 25897 12481 25996
rect 12618 25984 12624 26036
rect 12676 26024 12682 26036
rect 12676 25996 12756 26024
rect 12676 25984 12682 25996
rect 12728 25965 12756 25996
rect 13814 25984 13820 26036
rect 13872 26024 13878 26036
rect 14084 26027 14142 26033
rect 14084 26024 14096 26027
rect 13872 25996 14096 26024
rect 13872 25984 13878 25996
rect 14084 25993 14096 25996
rect 14130 25993 14142 26027
rect 14084 25987 14142 25993
rect 15102 25984 15108 26036
rect 15160 26024 15166 26036
rect 18877 26027 18935 26033
rect 18877 26024 18889 26027
rect 15160 25996 18889 26024
rect 15160 25984 15166 25996
rect 18877 25993 18889 25996
rect 18923 25993 18935 26027
rect 18877 25987 18935 25993
rect 19337 26027 19395 26033
rect 19337 25993 19349 26027
rect 19383 26024 19395 26027
rect 19426 26024 19432 26036
rect 19383 25996 19432 26024
rect 19383 25993 19395 25996
rect 19337 25987 19395 25993
rect 19426 25984 19432 25996
rect 19484 25984 19490 26036
rect 20073 26027 20131 26033
rect 20073 25993 20085 26027
rect 20119 26024 20131 26027
rect 20438 26024 20444 26036
rect 20119 25996 20444 26024
rect 20119 25993 20131 25996
rect 20073 25987 20131 25993
rect 20438 25984 20444 25996
rect 20496 25984 20502 26036
rect 23017 26027 23075 26033
rect 23017 26024 23029 26027
rect 20640 25996 23029 26024
rect 12713 25959 12771 25965
rect 12713 25925 12725 25959
rect 12759 25925 12771 25959
rect 12713 25919 12771 25925
rect 16301 25959 16359 25965
rect 16301 25925 16313 25959
rect 16347 25956 16359 25959
rect 16666 25956 16672 25968
rect 16347 25928 16672 25956
rect 16347 25925 16359 25928
rect 16301 25919 16359 25925
rect 16666 25916 16672 25928
rect 16724 25956 16730 25968
rect 17957 25959 18015 25965
rect 17957 25956 17969 25959
rect 16724 25928 17969 25956
rect 16724 25916 16730 25928
rect 17957 25925 17969 25928
rect 18003 25925 18015 25959
rect 19978 25956 19984 25968
rect 17957 25919 18015 25925
rect 18156 25928 19984 25956
rect 18156 25900 18184 25928
rect 19978 25916 19984 25928
rect 20036 25916 20042 25968
rect 20162 25916 20168 25968
rect 20220 25956 20226 25968
rect 20257 25959 20315 25965
rect 20257 25956 20269 25959
rect 20220 25928 20269 25956
rect 20220 25916 20226 25928
rect 20257 25925 20269 25928
rect 20303 25925 20315 25959
rect 20640 25956 20668 25996
rect 23017 25993 23029 25996
rect 23063 25993 23075 26027
rect 24213 26027 24271 26033
rect 24213 26024 24225 26027
rect 23017 25987 23075 25993
rect 23492 25996 24225 26024
rect 21085 25959 21143 25965
rect 20640 25928 20693 25956
rect 20257 25919 20315 25925
rect 11885 25891 11943 25897
rect 11624 25858 11836 25886
rect 11072 25820 11100 25848
rect 9416 25792 9628 25820
rect 9600 25764 9628 25792
rect 9968 25792 11100 25820
rect 11149 25823 11207 25829
rect 9048 25724 9536 25752
rect 9508 25696 9536 25724
rect 9582 25712 9588 25764
rect 9640 25752 9646 25764
rect 9968 25752 9996 25792
rect 11149 25789 11161 25823
rect 11195 25820 11207 25823
rect 11624 25820 11652 25858
rect 11808 25854 11836 25858
rect 11885 25857 11897 25891
rect 11931 25857 11943 25891
rect 11808 25829 11837 25854
rect 11885 25851 11943 25857
rect 12345 25891 12403 25897
rect 12345 25857 12357 25891
rect 12391 25857 12403 25891
rect 12345 25851 12403 25857
rect 12438 25891 12496 25897
rect 12438 25857 12450 25891
rect 12484 25857 12496 25891
rect 12438 25851 12496 25857
rect 11195 25792 11652 25820
rect 11702 25823 11760 25829
rect 11195 25789 11207 25792
rect 11149 25783 11207 25789
rect 11702 25789 11714 25823
rect 11748 25789 11760 25823
rect 11702 25783 11760 25789
rect 11793 25823 11851 25829
rect 11793 25789 11805 25823
rect 11839 25789 11851 25823
rect 11793 25783 11851 25789
rect 9640 25724 9996 25752
rect 11716 25752 11744 25783
rect 11974 25780 11980 25832
rect 12032 25780 12038 25832
rect 12360 25820 12388 25851
rect 12618 25848 12624 25900
rect 12676 25848 12682 25900
rect 12802 25848 12808 25900
rect 12860 25897 12866 25900
rect 12860 25888 12868 25897
rect 13817 25891 13875 25897
rect 13817 25888 13829 25891
rect 12860 25860 13829 25888
rect 12860 25851 12868 25860
rect 13817 25857 13829 25860
rect 13863 25857 13875 25891
rect 13817 25851 13875 25857
rect 12860 25848 12866 25851
rect 14458 25848 14464 25900
rect 14516 25848 14522 25900
rect 14826 25888 14832 25900
rect 14787 25860 14832 25888
rect 14826 25848 14832 25860
rect 14884 25848 14890 25900
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25857 14979 25891
rect 14921 25851 14979 25857
rect 12526 25820 12532 25832
rect 12360 25792 12532 25820
rect 12526 25780 12532 25792
rect 12584 25820 12590 25832
rect 14553 25823 14611 25829
rect 14553 25820 14565 25823
rect 12584 25792 14565 25820
rect 12584 25780 12590 25792
rect 14553 25789 14565 25792
rect 14599 25789 14611 25823
rect 14936 25820 14964 25851
rect 15010 25848 15016 25900
rect 15068 25848 15074 25900
rect 15194 25848 15200 25900
rect 15252 25848 15258 25900
rect 15930 25848 15936 25900
rect 15988 25848 15994 25900
rect 17589 25891 17647 25897
rect 17589 25857 17601 25891
rect 17635 25888 17647 25891
rect 17635 25860 18092 25888
rect 17635 25857 17647 25860
rect 17589 25851 17647 25857
rect 15102 25820 15108 25832
rect 14936 25792 15108 25820
rect 14553 25783 14611 25789
rect 15102 25780 15108 25792
rect 15160 25820 15166 25832
rect 15657 25823 15715 25829
rect 15657 25820 15669 25823
rect 15160 25792 15669 25820
rect 15160 25780 15166 25792
rect 15657 25789 15669 25792
rect 15703 25789 15715 25823
rect 15657 25783 15715 25789
rect 15838 25780 15844 25832
rect 15896 25820 15902 25832
rect 17405 25823 17463 25829
rect 17405 25820 17417 25823
rect 15896 25792 17417 25820
rect 15896 25780 15902 25792
rect 17405 25789 17417 25792
rect 17451 25789 17463 25823
rect 17405 25783 17463 25789
rect 17862 25780 17868 25832
rect 17920 25780 17926 25832
rect 18064 25820 18092 25860
rect 18138 25848 18144 25900
rect 18196 25848 18202 25900
rect 18414 25848 18420 25900
rect 18472 25848 18478 25900
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25857 18659 25891
rect 18601 25851 18659 25857
rect 18325 25823 18383 25829
rect 18325 25820 18337 25823
rect 18064 25792 18337 25820
rect 18325 25789 18337 25792
rect 18371 25820 18383 25823
rect 18509 25823 18567 25829
rect 18509 25820 18521 25823
rect 18371 25792 18521 25820
rect 18371 25789 18383 25792
rect 18325 25783 18383 25789
rect 18509 25789 18521 25792
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 11716 25724 12480 25752
rect 9640 25712 9646 25724
rect 12452 25696 12480 25724
rect 16482 25712 16488 25764
rect 16540 25752 16546 25764
rect 18616 25752 18644 25851
rect 18874 25848 18880 25900
rect 18932 25888 18938 25900
rect 20665 25897 20693 25928
rect 21085 25925 21097 25959
rect 21131 25956 21143 25959
rect 21358 25956 21364 25968
rect 21131 25928 21364 25956
rect 21131 25925 21143 25928
rect 21085 25919 21143 25925
rect 21358 25916 21364 25928
rect 21416 25916 21422 25968
rect 22741 25959 22799 25965
rect 22112 25928 22600 25956
rect 19061 25891 19119 25897
rect 19061 25888 19073 25891
rect 18932 25860 19073 25888
rect 18932 25848 18938 25860
rect 19061 25857 19073 25860
rect 19107 25857 19119 25891
rect 20625 25891 20693 25897
rect 19061 25851 19119 25857
rect 19260 25860 20576 25888
rect 18782 25780 18788 25832
rect 18840 25820 18846 25832
rect 19153 25823 19211 25829
rect 19153 25820 19165 25823
rect 18840 25792 19165 25820
rect 18840 25780 18846 25792
rect 19153 25789 19165 25792
rect 19199 25789 19211 25823
rect 19153 25783 19211 25789
rect 19260 25752 19288 25860
rect 19429 25823 19487 25829
rect 19429 25789 19441 25823
rect 19475 25789 19487 25823
rect 19429 25783 19487 25789
rect 16540 25724 19288 25752
rect 19444 25752 19472 25783
rect 19518 25780 19524 25832
rect 19576 25780 19582 25832
rect 19978 25780 19984 25832
rect 20036 25820 20042 25832
rect 20346 25820 20352 25832
rect 20036 25792 20352 25820
rect 20036 25780 20042 25792
rect 20346 25780 20352 25792
rect 20404 25780 20410 25832
rect 20548 25820 20576 25860
rect 20625 25857 20637 25891
rect 20671 25860 20693 25891
rect 20732 25860 21404 25888
rect 20671 25857 20683 25860
rect 20625 25851 20683 25857
rect 20732 25820 20760 25860
rect 20548 25792 20760 25820
rect 21174 25780 21180 25832
rect 21232 25780 21238 25832
rect 21376 25829 21404 25860
rect 22002 25848 22008 25900
rect 22060 25848 22066 25900
rect 22112 25897 22140 25928
rect 22572 25900 22600 25928
rect 22741 25925 22753 25959
rect 22787 25956 22799 25959
rect 22830 25956 22836 25968
rect 22787 25928 22836 25956
rect 22787 25925 22799 25928
rect 22741 25919 22799 25925
rect 22830 25916 22836 25928
rect 22888 25916 22894 25968
rect 23492 25965 23520 25996
rect 24213 25993 24225 25996
rect 24259 25993 24271 26027
rect 24213 25987 24271 25993
rect 29638 25984 29644 26036
rect 29696 26024 29702 26036
rect 29733 26027 29791 26033
rect 29733 26024 29745 26027
rect 29696 25996 29745 26024
rect 29696 25984 29702 25996
rect 29733 25993 29745 25996
rect 29779 25993 29791 26027
rect 29733 25987 29791 25993
rect 29901 26027 29959 26033
rect 29901 25993 29913 26027
rect 29947 26024 29959 26027
rect 30558 26024 30564 26036
rect 29947 25996 30564 26024
rect 29947 25993 29959 25996
rect 29901 25987 29959 25993
rect 30558 25984 30564 25996
rect 30616 25984 30622 26036
rect 32122 25984 32128 26036
rect 32180 25984 32186 26036
rect 32306 25984 32312 26036
rect 32364 26024 32370 26036
rect 32364 25996 32444 26024
rect 32364 25984 32370 25996
rect 23477 25959 23535 25965
rect 23477 25925 23489 25959
rect 23523 25925 23535 25959
rect 23477 25919 23535 25925
rect 24412 25928 24900 25956
rect 22097 25891 22155 25897
rect 22097 25857 22109 25891
rect 22143 25857 22155 25891
rect 22097 25851 22155 25857
rect 22281 25891 22339 25897
rect 22281 25857 22293 25891
rect 22327 25857 22339 25891
rect 22281 25851 22339 25857
rect 22373 25891 22431 25897
rect 22373 25857 22385 25891
rect 22419 25857 22431 25891
rect 22373 25851 22431 25857
rect 21361 25823 21419 25829
rect 21361 25789 21373 25823
rect 21407 25820 21419 25823
rect 21542 25820 21548 25832
rect 21407 25792 21548 25820
rect 21407 25789 21419 25792
rect 21361 25783 21419 25789
rect 21542 25780 21548 25792
rect 21600 25780 21606 25832
rect 20806 25752 20812 25764
rect 19444 25724 20812 25752
rect 16540 25712 16546 25724
rect 20806 25712 20812 25724
rect 20864 25712 20870 25764
rect 9306 25684 9312 25696
rect 8956 25656 9312 25684
rect 9306 25644 9312 25656
rect 9364 25644 9370 25696
rect 9398 25644 9404 25696
rect 9456 25644 9462 25696
rect 9490 25644 9496 25696
rect 9548 25684 9554 25696
rect 9766 25684 9772 25696
rect 9548 25656 9772 25684
rect 9548 25644 9554 25656
rect 9766 25644 9772 25656
rect 9824 25644 9830 25696
rect 10137 25687 10195 25693
rect 10137 25653 10149 25687
rect 10183 25684 10195 25687
rect 10686 25684 10692 25696
rect 10183 25656 10692 25684
rect 10183 25653 10195 25656
rect 10137 25647 10195 25653
rect 10686 25644 10692 25656
rect 10744 25644 10750 25696
rect 10962 25644 10968 25696
rect 11020 25684 11026 25696
rect 11517 25687 11575 25693
rect 11517 25684 11529 25687
rect 11020 25656 11529 25684
rect 11020 25644 11026 25656
rect 11517 25653 11529 25656
rect 11563 25653 11575 25687
rect 11517 25647 11575 25653
rect 12434 25644 12440 25696
rect 12492 25644 12498 25696
rect 12986 25644 12992 25696
rect 13044 25644 13050 25696
rect 14090 25644 14096 25696
rect 14148 25644 14154 25696
rect 17773 25687 17831 25693
rect 17773 25653 17785 25687
rect 17819 25684 17831 25687
rect 17862 25684 17868 25696
rect 17819 25656 17868 25684
rect 17819 25653 17831 25656
rect 17773 25647 17831 25653
rect 17862 25644 17868 25656
rect 17920 25644 17926 25696
rect 18874 25644 18880 25696
rect 18932 25684 18938 25696
rect 19610 25684 19616 25696
rect 18932 25656 19616 25684
rect 18932 25644 18938 25656
rect 19610 25644 19616 25656
rect 19668 25644 19674 25696
rect 19978 25644 19984 25696
rect 20036 25684 20042 25696
rect 20257 25687 20315 25693
rect 20257 25684 20269 25687
rect 20036 25656 20269 25684
rect 20036 25644 20042 25656
rect 20257 25653 20269 25656
rect 20303 25653 20315 25687
rect 20257 25647 20315 25653
rect 20346 25644 20352 25696
rect 20404 25684 20410 25696
rect 20717 25687 20775 25693
rect 20717 25684 20729 25687
rect 20404 25656 20729 25684
rect 20404 25644 20410 25656
rect 20717 25653 20729 25656
rect 20763 25653 20775 25687
rect 20717 25647 20775 25653
rect 21726 25644 21732 25696
rect 21784 25684 21790 25696
rect 21821 25687 21879 25693
rect 21821 25684 21833 25687
rect 21784 25656 21833 25684
rect 21784 25644 21790 25656
rect 21821 25653 21833 25656
rect 21867 25653 21879 25687
rect 22296 25684 22324 25851
rect 22388 25820 22416 25851
rect 22554 25848 22560 25900
rect 22612 25848 22618 25900
rect 23201 25891 23259 25897
rect 23201 25857 23213 25891
rect 23247 25857 23259 25891
rect 23201 25851 23259 25857
rect 23014 25820 23020 25832
rect 22388 25792 23020 25820
rect 23014 25780 23020 25792
rect 23072 25820 23078 25832
rect 23216 25820 23244 25851
rect 23566 25848 23572 25900
rect 23624 25848 23630 25900
rect 23658 25848 23664 25900
rect 23716 25888 23722 25900
rect 23716 25860 23761 25888
rect 23716 25848 23722 25860
rect 23842 25848 23848 25900
rect 23900 25848 23906 25900
rect 23934 25848 23940 25900
rect 23992 25848 23998 25900
rect 24075 25891 24133 25897
rect 24075 25857 24087 25891
rect 24121 25888 24133 25891
rect 24412 25888 24440 25928
rect 24872 25900 24900 25928
rect 24946 25916 24952 25968
rect 25004 25956 25010 25968
rect 25222 25956 25228 25968
rect 25004 25928 25228 25956
rect 25004 25916 25010 25928
rect 25222 25916 25228 25928
rect 25280 25956 25286 25968
rect 25280 25928 29592 25956
rect 25280 25916 25286 25928
rect 24121 25860 24440 25888
rect 24489 25891 24547 25897
rect 24121 25857 24133 25860
rect 24075 25851 24133 25857
rect 24489 25857 24501 25891
rect 24535 25857 24547 25891
rect 24489 25851 24547 25857
rect 23072 25792 23244 25820
rect 23385 25823 23443 25829
rect 23072 25780 23078 25792
rect 23385 25789 23397 25823
rect 23431 25820 23443 25823
rect 24305 25823 24363 25829
rect 24305 25820 24317 25823
rect 23431 25792 24317 25820
rect 23431 25789 23443 25792
rect 23385 25783 23443 25789
rect 24305 25789 24317 25792
rect 24351 25789 24363 25823
rect 24305 25783 24363 25789
rect 22925 25755 22983 25761
rect 22925 25721 22937 25755
rect 22971 25752 22983 25755
rect 24210 25752 24216 25764
rect 22971 25724 24216 25752
rect 22971 25721 22983 25724
rect 22925 25715 22983 25721
rect 24210 25712 24216 25724
rect 24268 25752 24274 25764
rect 24504 25752 24532 25851
rect 24578 25848 24584 25900
rect 24636 25848 24642 25900
rect 24854 25848 24860 25900
rect 24912 25848 24918 25900
rect 25314 25848 25320 25900
rect 25372 25848 25378 25900
rect 26050 25848 26056 25900
rect 26108 25848 26114 25900
rect 26602 25848 26608 25900
rect 26660 25888 26666 25900
rect 27525 25891 27583 25897
rect 27525 25888 27537 25891
rect 26660 25860 27537 25888
rect 26660 25848 26666 25860
rect 27525 25857 27537 25860
rect 27571 25857 27583 25891
rect 27525 25851 27583 25857
rect 27614 25848 27620 25900
rect 27672 25888 27678 25900
rect 27709 25891 27767 25897
rect 27709 25888 27721 25891
rect 27672 25860 27721 25888
rect 27672 25848 27678 25860
rect 27709 25857 27721 25860
rect 27755 25857 27767 25891
rect 27709 25851 27767 25857
rect 28905 25891 28963 25897
rect 28905 25857 28917 25891
rect 28951 25857 28963 25891
rect 28905 25851 28963 25857
rect 29089 25891 29147 25897
rect 29089 25857 29101 25891
rect 29135 25888 29147 25891
rect 29178 25888 29184 25900
rect 29135 25860 29184 25888
rect 29135 25857 29147 25860
rect 29089 25851 29147 25857
rect 28626 25820 28632 25832
rect 25976 25792 28632 25820
rect 25976 25761 26004 25792
rect 28626 25780 28632 25792
rect 28684 25820 28690 25832
rect 28920 25820 28948 25851
rect 29178 25848 29184 25860
rect 29236 25848 29242 25900
rect 29564 25897 29592 25928
rect 30006 25916 30012 25968
rect 30064 25956 30070 25968
rect 30101 25959 30159 25965
rect 30101 25956 30113 25959
rect 30064 25928 30113 25956
rect 30064 25916 30070 25928
rect 30101 25925 30113 25928
rect 30147 25925 30159 25959
rect 30101 25919 30159 25925
rect 29457 25891 29515 25897
rect 29457 25857 29469 25891
rect 29503 25857 29515 25891
rect 29457 25851 29515 25857
rect 29549 25891 29607 25897
rect 29549 25857 29561 25891
rect 29595 25857 29607 25891
rect 30576 25888 30604 25984
rect 32416 25965 32444 25996
rect 32582 25984 32588 26036
rect 32640 26024 32646 26036
rect 32640 25996 33456 26024
rect 32640 25984 32646 25996
rect 32401 25959 32459 25965
rect 32401 25925 32413 25959
rect 32447 25925 32459 25959
rect 32858 25956 32864 25968
rect 32401 25919 32459 25925
rect 32692 25928 32864 25956
rect 31018 25888 31024 25900
rect 30576 25860 31024 25888
rect 29549 25851 29607 25857
rect 28684 25792 28948 25820
rect 28997 25823 29055 25829
rect 28684 25780 28690 25792
rect 28997 25789 29009 25823
rect 29043 25820 29055 25823
rect 29362 25820 29368 25832
rect 29043 25792 29368 25820
rect 29043 25789 29055 25792
rect 28997 25783 29055 25789
rect 29362 25780 29368 25792
rect 29420 25780 29426 25832
rect 29472 25820 29500 25851
rect 31018 25848 31024 25860
rect 31076 25888 31082 25900
rect 32030 25888 32036 25900
rect 31076 25860 32036 25888
rect 31076 25848 31082 25860
rect 32030 25848 32036 25860
rect 32088 25888 32094 25900
rect 32277 25891 32335 25897
rect 32277 25888 32289 25891
rect 32088 25860 32289 25888
rect 32088 25848 32094 25860
rect 32277 25857 32289 25860
rect 32323 25857 32335 25891
rect 32277 25851 32335 25857
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25888 32551 25891
rect 32582 25888 32588 25900
rect 32539 25860 32588 25888
rect 32539 25857 32551 25860
rect 32493 25851 32551 25857
rect 32582 25848 32588 25860
rect 32640 25848 32646 25900
rect 32692 25897 32720 25928
rect 32858 25916 32864 25928
rect 32916 25916 32922 25968
rect 33428 25956 33456 25996
rect 33502 25984 33508 26036
rect 33560 26024 33566 26036
rect 34698 26024 34704 26036
rect 33560 25996 34704 26024
rect 33560 25984 33566 25996
rect 34698 25984 34704 25996
rect 34756 25984 34762 26036
rect 34422 25956 34428 25968
rect 33428 25928 33640 25956
rect 33612 25922 33640 25928
rect 33704 25928 34428 25956
rect 33704 25922 33732 25928
rect 32677 25891 32735 25897
rect 32677 25857 32689 25891
rect 32723 25857 32735 25891
rect 32677 25851 32735 25857
rect 32769 25891 32827 25897
rect 32769 25857 32781 25891
rect 32815 25857 32827 25891
rect 32769 25851 32827 25857
rect 32784 25820 32812 25851
rect 33318 25848 33324 25900
rect 33376 25888 33382 25900
rect 33505 25891 33563 25897
rect 33612 25894 33732 25922
rect 34422 25916 34428 25928
rect 34480 25956 34486 25968
rect 34480 25928 34822 25956
rect 34480 25916 34486 25928
rect 33781 25894 33839 25897
rect 33505 25888 33517 25891
rect 33376 25860 33517 25888
rect 33376 25848 33382 25860
rect 33505 25857 33517 25860
rect 33551 25857 33563 25891
rect 33505 25851 33563 25857
rect 33781 25891 33916 25894
rect 33781 25857 33793 25891
rect 33827 25888 33916 25891
rect 33962 25888 33968 25900
rect 33827 25866 33968 25888
rect 33827 25857 33839 25866
rect 33888 25860 33968 25866
rect 33781 25851 33839 25857
rect 33962 25848 33968 25860
rect 34020 25848 34026 25900
rect 34054 25848 34060 25900
rect 34112 25848 34118 25900
rect 29472 25792 29960 25820
rect 24268 25724 24532 25752
rect 25961 25755 26019 25761
rect 24268 25712 24274 25724
rect 25961 25721 25973 25755
rect 26007 25721 26019 25755
rect 25961 25715 26019 25721
rect 27709 25755 27767 25761
rect 27709 25721 27721 25755
rect 27755 25752 27767 25755
rect 29730 25752 29736 25764
rect 27755 25724 29736 25752
rect 27755 25721 27767 25724
rect 27709 25715 27767 25721
rect 29730 25712 29736 25724
rect 29788 25712 29794 25764
rect 29932 25696 29960 25792
rect 32416 25792 32812 25820
rect 33689 25823 33747 25829
rect 32416 25764 32444 25792
rect 33689 25789 33701 25823
rect 33735 25820 33747 25823
rect 33870 25820 33876 25832
rect 33735 25792 33876 25820
rect 33735 25789 33747 25792
rect 33689 25783 33747 25789
rect 33870 25780 33876 25792
rect 33928 25780 33934 25832
rect 34333 25823 34391 25829
rect 34333 25820 34345 25823
rect 33980 25792 34345 25820
rect 32122 25712 32128 25764
rect 32180 25752 32186 25764
rect 32398 25752 32404 25764
rect 32180 25724 32404 25752
rect 32180 25712 32186 25724
rect 32398 25712 32404 25724
rect 32456 25712 32462 25764
rect 33980 25761 34008 25792
rect 34333 25789 34345 25792
rect 34379 25789 34391 25823
rect 34333 25783 34391 25789
rect 36078 25780 36084 25832
rect 36136 25780 36142 25832
rect 33965 25755 34023 25761
rect 32508 25724 33640 25752
rect 23385 25687 23443 25693
rect 23385 25684 23397 25687
rect 22296 25656 23397 25684
rect 21821 25647 21879 25653
rect 23385 25653 23397 25656
rect 23431 25684 23443 25687
rect 23474 25684 23480 25696
rect 23431 25656 23480 25684
rect 23431 25653 23443 25656
rect 23385 25647 23443 25653
rect 23474 25644 23480 25656
rect 23532 25644 23538 25696
rect 23934 25644 23940 25696
rect 23992 25684 23998 25696
rect 24765 25687 24823 25693
rect 24765 25684 24777 25687
rect 23992 25656 24777 25684
rect 23992 25644 23998 25656
rect 24765 25653 24777 25656
rect 24811 25653 24823 25687
rect 24765 25647 24823 25653
rect 29273 25687 29331 25693
rect 29273 25653 29285 25687
rect 29319 25684 29331 25687
rect 29362 25684 29368 25696
rect 29319 25656 29368 25684
rect 29319 25653 29331 25656
rect 29273 25647 29331 25653
rect 29362 25644 29368 25656
rect 29420 25644 29426 25696
rect 29914 25644 29920 25696
rect 29972 25644 29978 25696
rect 30190 25644 30196 25696
rect 30248 25684 30254 25696
rect 32508 25684 32536 25724
rect 30248 25656 32536 25684
rect 30248 25644 30254 25656
rect 33502 25644 33508 25696
rect 33560 25644 33566 25696
rect 33612 25684 33640 25724
rect 33965 25721 33977 25755
rect 34011 25721 34023 25755
rect 33965 25715 34023 25721
rect 35434 25684 35440 25696
rect 33612 25656 35440 25684
rect 35434 25644 35440 25656
rect 35492 25644 35498 25696
rect 1104 25594 36432 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 36432 25594
rect 1104 25520 36432 25542
rect 3142 25440 3148 25492
rect 3200 25480 3206 25492
rect 4614 25480 4620 25492
rect 3200 25452 4620 25480
rect 3200 25440 3206 25452
rect 4614 25440 4620 25452
rect 4672 25440 4678 25492
rect 4706 25440 4712 25492
rect 4764 25480 4770 25492
rect 4801 25483 4859 25489
rect 4801 25480 4813 25483
rect 4764 25452 4813 25480
rect 4764 25440 4770 25452
rect 4801 25449 4813 25452
rect 4847 25449 4859 25483
rect 4801 25443 4859 25449
rect 6641 25483 6699 25489
rect 6641 25449 6653 25483
rect 6687 25480 6699 25483
rect 9398 25480 9404 25492
rect 6687 25452 9404 25480
rect 6687 25449 6699 25452
rect 6641 25443 6699 25449
rect 9398 25440 9404 25452
rect 9456 25440 9462 25492
rect 9766 25440 9772 25492
rect 9824 25440 9830 25492
rect 10134 25440 10140 25492
rect 10192 25480 10198 25492
rect 10410 25480 10416 25492
rect 10192 25452 10416 25480
rect 10192 25440 10198 25452
rect 10410 25440 10416 25452
rect 10468 25480 10474 25492
rect 10962 25480 10968 25492
rect 10468 25452 10968 25480
rect 10468 25440 10474 25452
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 18141 25483 18199 25489
rect 18141 25449 18153 25483
rect 18187 25480 18199 25483
rect 18414 25480 18420 25492
rect 18187 25452 18420 25480
rect 18187 25449 18199 25452
rect 18141 25443 18199 25449
rect 18414 25440 18420 25452
rect 18472 25440 18478 25492
rect 19613 25483 19671 25489
rect 19613 25449 19625 25483
rect 19659 25480 19671 25483
rect 19794 25480 19800 25492
rect 19659 25452 19800 25480
rect 19659 25449 19671 25452
rect 19613 25443 19671 25449
rect 19794 25440 19800 25452
rect 19852 25440 19858 25492
rect 21542 25480 21548 25492
rect 19904 25452 21548 25480
rect 7374 25372 7380 25424
rect 7432 25412 7438 25424
rect 8202 25412 8208 25424
rect 7432 25384 8208 25412
rect 7432 25372 7438 25384
rect 8202 25372 8208 25384
rect 8260 25372 8266 25424
rect 8478 25372 8484 25424
rect 8536 25412 8542 25424
rect 8846 25412 8852 25424
rect 8536 25384 8852 25412
rect 8536 25372 8542 25384
rect 8846 25372 8852 25384
rect 8904 25372 8910 25424
rect 9030 25372 9036 25424
rect 9088 25412 9094 25424
rect 11146 25412 11152 25424
rect 9088 25384 11152 25412
rect 9088 25372 9094 25384
rect 11146 25372 11152 25384
rect 11204 25412 11210 25424
rect 11974 25412 11980 25424
rect 11204 25384 11980 25412
rect 11204 25372 11210 25384
rect 11974 25372 11980 25384
rect 12032 25372 12038 25424
rect 15838 25412 15844 25424
rect 14660 25384 15844 25412
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2866 25344 2872 25356
rect 1443 25316 2872 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2866 25304 2872 25316
rect 2924 25344 2930 25356
rect 4525 25347 4583 25353
rect 4525 25344 4537 25347
rect 2924 25316 4537 25344
rect 2924 25304 2930 25316
rect 4525 25313 4537 25316
rect 4571 25313 4583 25347
rect 4525 25307 4583 25313
rect 5258 25304 5264 25356
rect 5316 25304 5322 25356
rect 5445 25347 5503 25353
rect 5445 25313 5457 25347
rect 5491 25344 5503 25347
rect 5534 25344 5540 25356
rect 5491 25316 5540 25344
rect 5491 25313 5503 25316
rect 5445 25307 5503 25313
rect 5534 25304 5540 25316
rect 5592 25304 5598 25356
rect 6914 25304 6920 25356
rect 6972 25344 6978 25356
rect 7285 25347 7343 25353
rect 6972 25316 7236 25344
rect 6972 25304 6978 25316
rect 7208 25288 7236 25316
rect 7285 25313 7297 25347
rect 7331 25344 7343 25347
rect 8113 25347 8171 25353
rect 8113 25344 8125 25347
rect 7331 25316 8125 25344
rect 7331 25313 7343 25316
rect 7285 25307 7343 25313
rect 8113 25313 8125 25316
rect 8159 25313 8171 25347
rect 8113 25307 8171 25313
rect 8297 25347 8355 25353
rect 8297 25313 8309 25347
rect 8343 25344 8355 25347
rect 9953 25347 10011 25353
rect 9953 25344 9965 25347
rect 8343 25316 9965 25344
rect 8343 25313 8355 25316
rect 8297 25307 8355 25313
rect 9953 25313 9965 25316
rect 9999 25313 10011 25347
rect 11882 25344 11888 25356
rect 9953 25307 10011 25313
rect 11716 25316 11888 25344
rect 2774 25236 2780 25288
rect 2832 25276 2838 25288
rect 3970 25276 3976 25288
rect 2832 25248 3976 25276
rect 2832 25236 2838 25248
rect 3970 25236 3976 25248
rect 4028 25236 4034 25288
rect 5902 25236 5908 25288
rect 5960 25236 5966 25288
rect 6549 25279 6607 25285
rect 6549 25245 6561 25279
rect 6595 25276 6607 25279
rect 6595 25248 7052 25276
rect 6595 25245 6607 25248
rect 6549 25239 6607 25245
rect 1670 25168 1676 25220
rect 1728 25168 1734 25220
rect 3789 25211 3847 25217
rect 3789 25177 3801 25211
rect 3835 25208 3847 25211
rect 4062 25208 4068 25220
rect 3835 25180 4068 25208
rect 3835 25177 3847 25180
rect 3789 25171 3847 25177
rect 4062 25168 4068 25180
rect 4120 25168 4126 25220
rect 6086 25168 6092 25220
rect 6144 25208 6150 25220
rect 6457 25211 6515 25217
rect 6457 25208 6469 25211
rect 6144 25180 6469 25208
rect 6144 25168 6150 25180
rect 6457 25177 6469 25180
rect 6503 25177 6515 25211
rect 6457 25171 6515 25177
rect 6822 25168 6828 25220
rect 6880 25168 6886 25220
rect 6914 25168 6920 25220
rect 6972 25168 6978 25220
rect 2314 25100 2320 25152
rect 2372 25140 2378 25152
rect 3142 25140 3148 25152
rect 2372 25112 3148 25140
rect 2372 25100 2378 25112
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 4614 25100 4620 25152
rect 4672 25140 4678 25152
rect 5169 25143 5227 25149
rect 5169 25140 5181 25143
rect 4672 25112 5181 25140
rect 4672 25100 4678 25112
rect 5169 25109 5181 25112
rect 5215 25140 5227 25143
rect 5442 25140 5448 25152
rect 5215 25112 5448 25140
rect 5215 25109 5227 25112
rect 5169 25103 5227 25109
rect 5442 25100 5448 25112
rect 5500 25100 5506 25152
rect 5718 25100 5724 25152
rect 5776 25100 5782 25152
rect 7024 25140 7052 25248
rect 7190 25236 7196 25288
rect 7248 25236 7254 25288
rect 7374 25236 7380 25288
rect 7432 25276 7438 25288
rect 7650 25276 7656 25288
rect 7432 25248 7656 25276
rect 7432 25236 7438 25248
rect 7650 25236 7656 25248
rect 7708 25236 7714 25288
rect 8018 25236 8024 25288
rect 8076 25236 8082 25288
rect 8202 25236 8208 25288
rect 8260 25236 8266 25288
rect 8478 25236 8484 25288
rect 8536 25276 8542 25288
rect 9217 25279 9275 25285
rect 9217 25276 9229 25279
rect 8536 25248 9229 25276
rect 8536 25236 8542 25248
rect 9217 25245 9229 25248
rect 9263 25245 9275 25279
rect 9217 25239 9275 25245
rect 9398 25236 9404 25288
rect 9456 25236 9462 25288
rect 9582 25236 9588 25288
rect 9640 25236 9646 25288
rect 9766 25236 9772 25288
rect 9824 25276 9830 25288
rect 9861 25279 9919 25285
rect 9861 25276 9873 25279
rect 9824 25248 9873 25276
rect 9824 25236 9830 25248
rect 9861 25245 9873 25248
rect 9907 25245 9919 25279
rect 9861 25239 9919 25245
rect 10042 25236 10048 25288
rect 10100 25236 10106 25288
rect 10962 25236 10968 25288
rect 11020 25276 11026 25288
rect 11517 25279 11575 25285
rect 11517 25276 11529 25279
rect 11020 25248 11529 25276
rect 11020 25236 11026 25248
rect 11517 25245 11529 25248
rect 11563 25245 11575 25279
rect 11517 25239 11575 25245
rect 11606 25236 11612 25288
rect 11664 25236 11670 25288
rect 11716 25285 11744 25316
rect 11882 25304 11888 25316
rect 11940 25304 11946 25356
rect 11701 25279 11759 25285
rect 11701 25245 11713 25279
rect 11747 25245 11759 25279
rect 11701 25239 11759 25245
rect 14458 25236 14464 25288
rect 14516 25236 14522 25288
rect 14660 25285 14688 25384
rect 15838 25372 15844 25384
rect 15896 25372 15902 25424
rect 16577 25415 16635 25421
rect 16577 25381 16589 25415
rect 16623 25381 16635 25415
rect 18874 25412 18880 25424
rect 16577 25375 16635 25381
rect 17604 25384 18880 25412
rect 14921 25347 14979 25353
rect 14921 25313 14933 25347
rect 14967 25344 14979 25347
rect 15010 25344 15016 25356
rect 14967 25316 15016 25344
rect 14967 25313 14979 25316
rect 14921 25307 14979 25313
rect 15010 25304 15016 25316
rect 15068 25304 15074 25356
rect 16393 25347 16451 25353
rect 16393 25344 16405 25347
rect 15304 25316 16405 25344
rect 15304 25288 15332 25316
rect 16393 25313 16405 25316
rect 16439 25344 16451 25347
rect 16592 25344 16620 25375
rect 16439 25316 16620 25344
rect 16439 25313 16451 25316
rect 16393 25307 16451 25313
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 14645 25279 14703 25285
rect 14645 25245 14657 25279
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 8036 25208 8064 25236
rect 9030 25208 9036 25220
rect 8036 25180 9036 25208
rect 9030 25168 9036 25180
rect 9088 25168 9094 25220
rect 9493 25211 9551 25217
rect 9493 25177 9505 25211
rect 9539 25208 9551 25211
rect 10870 25208 10876 25220
rect 9539 25180 10876 25208
rect 9539 25177 9551 25180
rect 9493 25171 9551 25177
rect 10870 25168 10876 25180
rect 10928 25168 10934 25220
rect 11330 25168 11336 25220
rect 11388 25208 11394 25220
rect 11425 25211 11483 25217
rect 11425 25208 11437 25211
rect 11388 25180 11437 25208
rect 11388 25168 11394 25180
rect 11425 25177 11437 25180
rect 11471 25177 11483 25211
rect 11425 25171 11483 25177
rect 11885 25211 11943 25217
rect 11885 25177 11897 25211
rect 11931 25208 11943 25211
rect 12158 25208 12164 25220
rect 11931 25180 12164 25208
rect 11931 25177 11943 25180
rect 11885 25171 11943 25177
rect 12158 25168 12164 25180
rect 12216 25208 12222 25220
rect 13078 25208 13084 25220
rect 12216 25180 13084 25208
rect 12216 25168 12222 25180
rect 13078 25168 13084 25180
rect 13136 25208 13142 25220
rect 13446 25208 13452 25220
rect 13136 25180 13452 25208
rect 13136 25168 13142 25180
rect 13446 25168 13452 25180
rect 13504 25168 13510 25220
rect 13814 25168 13820 25220
rect 13872 25208 13878 25220
rect 14274 25208 14280 25220
rect 13872 25180 14280 25208
rect 13872 25168 13878 25180
rect 14274 25168 14280 25180
rect 14332 25208 14338 25220
rect 14568 25208 14596 25239
rect 15102 25236 15108 25288
rect 15160 25236 15166 25288
rect 15286 25236 15292 25288
rect 15344 25236 15350 25288
rect 15381 25279 15439 25285
rect 15381 25245 15393 25279
rect 15427 25276 15439 25279
rect 16209 25279 16267 25285
rect 16209 25276 16221 25279
rect 15427 25248 16221 25276
rect 15427 25245 15439 25248
rect 15381 25239 15439 25245
rect 16209 25245 16221 25248
rect 16255 25276 16267 25279
rect 16298 25276 16304 25288
rect 16255 25248 16304 25276
rect 16255 25245 16267 25248
rect 16209 25239 16267 25245
rect 16298 25236 16304 25248
rect 16356 25236 16362 25288
rect 16758 25236 16764 25288
rect 16816 25236 16822 25288
rect 16942 25236 16948 25288
rect 17000 25276 17006 25288
rect 17604 25285 17632 25384
rect 18874 25372 18880 25384
rect 18932 25372 18938 25424
rect 18966 25372 18972 25424
rect 19024 25412 19030 25424
rect 19904 25412 19932 25452
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 21818 25440 21824 25492
rect 21876 25480 21882 25492
rect 22830 25480 22836 25492
rect 21876 25452 22836 25480
rect 21876 25440 21882 25452
rect 22830 25440 22836 25452
rect 22888 25440 22894 25492
rect 23290 25440 23296 25492
rect 23348 25440 23354 25492
rect 24854 25440 24860 25492
rect 24912 25440 24918 25492
rect 26418 25440 26424 25492
rect 26476 25480 26482 25492
rect 33042 25480 33048 25492
rect 26476 25452 33048 25480
rect 26476 25440 26482 25452
rect 33042 25440 33048 25452
rect 33100 25440 33106 25492
rect 33318 25440 33324 25492
rect 33376 25440 33382 25492
rect 33594 25440 33600 25492
rect 33652 25480 33658 25492
rect 33781 25483 33839 25489
rect 33781 25480 33793 25483
rect 33652 25452 33793 25480
rect 33652 25440 33658 25452
rect 33781 25449 33793 25452
rect 33827 25449 33839 25483
rect 33781 25443 33839 25449
rect 34422 25440 34428 25492
rect 34480 25480 34486 25492
rect 35897 25483 35955 25489
rect 35897 25480 35909 25483
rect 34480 25452 35909 25480
rect 34480 25440 34486 25452
rect 35897 25449 35909 25452
rect 35943 25449 35955 25483
rect 35897 25443 35955 25449
rect 19024 25384 19932 25412
rect 19024 25372 19030 25384
rect 20070 25372 20076 25424
rect 20128 25412 20134 25424
rect 20349 25415 20407 25421
rect 20349 25412 20361 25415
rect 20128 25384 20361 25412
rect 20128 25372 20134 25384
rect 20349 25381 20361 25384
rect 20395 25381 20407 25415
rect 20349 25375 20407 25381
rect 20548 25384 22416 25412
rect 20548 25344 20576 25384
rect 21082 25344 21088 25356
rect 17880 25316 20576 25344
rect 20640 25316 21088 25344
rect 17880 25285 17908 25316
rect 17589 25279 17647 25285
rect 17589 25276 17601 25279
rect 17000 25248 17601 25276
rect 17000 25236 17006 25248
rect 17589 25245 17601 25248
rect 17635 25245 17647 25279
rect 17589 25239 17647 25245
rect 17865 25279 17923 25285
rect 17865 25245 17877 25279
rect 17911 25245 17923 25279
rect 17865 25239 17923 25245
rect 17957 25279 18015 25285
rect 17957 25245 17969 25279
rect 18003 25276 18015 25279
rect 18874 25276 18880 25288
rect 18003 25248 18880 25276
rect 18003 25245 18015 25248
rect 17957 25239 18015 25245
rect 18874 25236 18880 25248
rect 18932 25236 18938 25288
rect 18969 25279 19027 25285
rect 18969 25245 18981 25279
rect 19015 25276 19027 25279
rect 20640 25276 20668 25316
rect 21082 25304 21088 25316
rect 21140 25304 21146 25356
rect 21634 25344 21640 25356
rect 21376 25316 21640 25344
rect 19015 25248 20668 25276
rect 19015 25245 19027 25248
rect 18969 25239 19027 25245
rect 20714 25236 20720 25288
rect 20772 25236 20778 25288
rect 20901 25279 20959 25285
rect 20901 25245 20913 25279
rect 20947 25276 20959 25279
rect 21376 25276 21404 25316
rect 21634 25304 21640 25316
rect 21692 25304 21698 25356
rect 22388 25344 22416 25384
rect 23014 25372 23020 25424
rect 23072 25412 23078 25424
rect 23477 25415 23535 25421
rect 23477 25412 23489 25415
rect 23072 25384 23489 25412
rect 23072 25372 23078 25384
rect 23477 25381 23489 25384
rect 23523 25412 23535 25415
rect 23658 25412 23664 25424
rect 23523 25384 23664 25412
rect 23523 25381 23535 25384
rect 23477 25375 23535 25381
rect 23658 25372 23664 25384
rect 23716 25372 23722 25424
rect 25038 25372 25044 25424
rect 25096 25372 25102 25424
rect 32122 25372 32128 25424
rect 32180 25372 32186 25424
rect 32769 25415 32827 25421
rect 32769 25381 32781 25415
rect 32815 25412 32827 25415
rect 33689 25415 33747 25421
rect 33689 25412 33701 25415
rect 32815 25384 33701 25412
rect 32815 25381 32827 25384
rect 32769 25375 32827 25381
rect 33689 25381 33701 25384
rect 33735 25381 33747 25415
rect 33689 25375 33747 25381
rect 23201 25347 23259 25353
rect 23201 25344 23213 25347
rect 22388 25316 23213 25344
rect 23201 25313 23213 25316
rect 23247 25344 23259 25347
rect 23382 25344 23388 25356
rect 23247 25316 23388 25344
rect 23247 25313 23259 25316
rect 23201 25307 23259 25313
rect 23382 25304 23388 25316
rect 23440 25304 23446 25356
rect 25314 25304 25320 25356
rect 25372 25344 25378 25356
rect 32030 25344 32036 25356
rect 25372 25316 32036 25344
rect 25372 25304 25378 25316
rect 32030 25304 32036 25316
rect 32088 25304 32094 25356
rect 32140 25295 32168 25372
rect 32125 25289 32183 25295
rect 20947 25248 21404 25276
rect 21453 25279 21511 25285
rect 20947 25245 20959 25248
rect 20901 25239 20959 25245
rect 21453 25245 21465 25279
rect 21499 25245 21511 25279
rect 21453 25239 21511 25245
rect 14332 25180 14596 25208
rect 14737 25211 14795 25217
rect 14332 25168 14338 25180
rect 14737 25177 14749 25211
rect 14783 25208 14795 25211
rect 15930 25208 15936 25220
rect 14783 25180 15936 25208
rect 14783 25177 14795 25180
rect 14737 25171 14795 25177
rect 15930 25168 15936 25180
rect 15988 25168 15994 25220
rect 16022 25168 16028 25220
rect 16080 25168 16086 25220
rect 16666 25208 16672 25220
rect 16500 25180 16672 25208
rect 13722 25140 13728 25152
rect 7024 25112 13728 25140
rect 13722 25100 13728 25112
rect 13780 25100 13786 25152
rect 14826 25100 14832 25152
rect 14884 25140 14890 25152
rect 15105 25143 15163 25149
rect 15105 25140 15117 25143
rect 14884 25112 15117 25140
rect 14884 25100 14890 25112
rect 15105 25109 15117 25112
rect 15151 25109 15163 25143
rect 15105 25103 15163 25109
rect 15838 25100 15844 25152
rect 15896 25100 15902 25152
rect 16117 25143 16175 25149
rect 16117 25109 16129 25143
rect 16163 25140 16175 25143
rect 16500 25140 16528 25180
rect 16666 25168 16672 25180
rect 16724 25168 16730 25220
rect 17773 25211 17831 25217
rect 17773 25177 17785 25211
rect 17819 25177 17831 25211
rect 17773 25171 17831 25177
rect 16163 25112 16528 25140
rect 16163 25109 16175 25112
rect 16117 25103 16175 25109
rect 16758 25100 16764 25152
rect 16816 25140 16822 25152
rect 17788 25140 17816 25171
rect 18598 25168 18604 25220
rect 18656 25168 18662 25220
rect 19797 25211 19855 25217
rect 19797 25177 19809 25211
rect 19843 25208 19855 25211
rect 20162 25208 20168 25220
rect 19843 25180 20168 25208
rect 19843 25177 19855 25180
rect 19797 25171 19855 25177
rect 20162 25168 20168 25180
rect 20220 25168 20226 25220
rect 20349 25211 20407 25217
rect 20349 25177 20361 25211
rect 20395 25208 20407 25211
rect 21468 25208 21496 25239
rect 21542 25236 21548 25288
rect 21600 25236 21606 25288
rect 21726 25236 21732 25288
rect 21784 25236 21790 25288
rect 21821 25279 21879 25285
rect 21821 25245 21833 25279
rect 21867 25276 21879 25279
rect 22738 25276 22744 25288
rect 21867 25248 22744 25276
rect 21867 25245 21879 25248
rect 21821 25239 21879 25245
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 23109 25279 23167 25285
rect 23109 25245 23121 25279
rect 23155 25276 23167 25279
rect 24210 25276 24216 25288
rect 23155 25248 24216 25276
rect 23155 25245 23167 25248
rect 23109 25239 23167 25245
rect 24210 25236 24216 25248
rect 24268 25236 24274 25288
rect 25406 25236 25412 25288
rect 25464 25276 25470 25288
rect 28994 25276 29000 25288
rect 25464 25248 29000 25276
rect 25464 25236 25470 25248
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 32125 25255 32137 25289
rect 32171 25255 32183 25289
rect 32263 25279 32321 25285
rect 32263 25276 32275 25279
rect 32248 25266 32275 25276
rect 32125 25249 32183 25255
rect 21913 25211 21971 25217
rect 21913 25208 21925 25211
rect 20395 25180 20852 25208
rect 21468 25180 21925 25208
rect 20395 25177 20407 25180
rect 20349 25171 20407 25177
rect 16816 25112 17816 25140
rect 19889 25143 19947 25149
rect 16816 25100 16822 25112
rect 19889 25109 19901 25143
rect 19935 25140 19947 25143
rect 20438 25140 20444 25152
rect 19935 25112 20444 25140
rect 19935 25109 19947 25112
rect 19889 25103 19947 25109
rect 20438 25100 20444 25112
rect 20496 25100 20502 25152
rect 20530 25100 20536 25152
rect 20588 25100 20594 25152
rect 20824 25140 20852 25180
rect 21913 25177 21925 25180
rect 21959 25177 21971 25211
rect 21913 25171 21971 25177
rect 22097 25211 22155 25217
rect 22097 25177 22109 25211
rect 22143 25208 22155 25211
rect 22186 25208 22192 25220
rect 22143 25180 22192 25208
rect 22143 25177 22155 25180
rect 22097 25171 22155 25177
rect 22186 25168 22192 25180
rect 22244 25168 22250 25220
rect 22281 25211 22339 25217
rect 22281 25177 22293 25211
rect 22327 25208 22339 25211
rect 23014 25208 23020 25220
rect 22327 25180 23020 25208
rect 22327 25177 22339 25180
rect 22281 25171 22339 25177
rect 23014 25168 23020 25180
rect 23072 25168 23078 25220
rect 25317 25211 25375 25217
rect 25317 25177 25329 25211
rect 25363 25208 25375 25211
rect 26050 25208 26056 25220
rect 25363 25180 26056 25208
rect 25363 25177 25375 25180
rect 25317 25171 25375 25177
rect 26050 25168 26056 25180
rect 26108 25208 26114 25220
rect 32122 25208 32128 25220
rect 26108 25180 32128 25208
rect 26108 25168 26114 25180
rect 32122 25168 32128 25180
rect 32180 25168 32186 25220
rect 32230 25214 32236 25266
rect 32309 25245 32321 25279
rect 32617 25279 32675 25285
rect 32288 25239 32321 25245
rect 32288 25214 32294 25239
rect 32401 25211 32459 25217
rect 32401 25177 32413 25211
rect 32447 25177 32459 25211
rect 32490 25202 32496 25254
rect 32548 25202 32554 25254
rect 32617 25245 32629 25279
rect 32663 25276 32675 25279
rect 32766 25276 32772 25288
rect 32663 25248 32772 25276
rect 32663 25245 32675 25248
rect 32617 25239 32675 25245
rect 32766 25236 32772 25248
rect 32824 25236 32830 25288
rect 33597 25279 33655 25285
rect 33597 25245 33609 25279
rect 33643 25276 33655 25279
rect 33686 25276 33692 25288
rect 33643 25248 33692 25276
rect 33643 25245 33655 25248
rect 33597 25239 33655 25245
rect 33686 25236 33692 25248
rect 33744 25236 33750 25288
rect 33778 25236 33784 25288
rect 33836 25276 33842 25288
rect 34057 25279 34115 25285
rect 34057 25276 34069 25279
rect 33836 25248 34069 25276
rect 33836 25236 33842 25248
rect 34057 25245 34069 25248
rect 34103 25245 34115 25279
rect 34057 25239 34115 25245
rect 35434 25236 35440 25288
rect 35492 25276 35498 25288
rect 35713 25279 35771 25285
rect 35713 25276 35725 25279
rect 35492 25248 35725 25276
rect 35492 25236 35498 25248
rect 35713 25245 35725 25248
rect 35759 25245 35771 25279
rect 35713 25239 35771 25245
rect 36078 25208 36084 25220
rect 32401 25171 32459 25177
rect 32784 25180 36084 25208
rect 21269 25143 21327 25149
rect 21269 25140 21281 25143
rect 20824 25112 21281 25140
rect 21269 25109 21281 25112
rect 21315 25109 21327 25143
rect 21269 25103 21327 25109
rect 22002 25100 22008 25152
rect 22060 25140 22066 25152
rect 24854 25140 24860 25152
rect 22060 25112 24860 25140
rect 22060 25100 22066 25112
rect 24854 25100 24860 25112
rect 24912 25100 24918 25152
rect 28258 25100 28264 25152
rect 28316 25140 28322 25152
rect 30006 25140 30012 25152
rect 28316 25112 30012 25140
rect 28316 25100 28322 25112
rect 30006 25100 30012 25112
rect 30064 25100 30070 25152
rect 32140 25140 32168 25168
rect 32416 25140 32444 25171
rect 32784 25140 32812 25180
rect 36078 25168 36084 25180
rect 36136 25168 36142 25220
rect 32140 25112 32812 25140
rect 33962 25100 33968 25152
rect 34020 25140 34026 25152
rect 34606 25140 34612 25152
rect 34020 25112 34612 25140
rect 34020 25100 34026 25112
rect 34606 25100 34612 25112
rect 34664 25100 34670 25152
rect 1104 25050 36432 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 36432 25050
rect 1104 24976 36432 24998
rect 3970 24896 3976 24948
rect 4028 24936 4034 24948
rect 4028 24908 5304 24936
rect 4028 24896 4034 24908
rect 2498 24828 2504 24880
rect 2556 24868 2562 24880
rect 2593 24871 2651 24877
rect 2593 24868 2605 24871
rect 2556 24840 2605 24868
rect 2556 24828 2562 24840
rect 2593 24837 2605 24840
rect 2639 24837 2651 24871
rect 2593 24831 2651 24837
rect 2685 24871 2743 24877
rect 2685 24837 2697 24871
rect 2731 24868 2743 24871
rect 3142 24868 3148 24880
rect 2731 24840 3148 24868
rect 2731 24837 2743 24840
rect 2685 24831 2743 24837
rect 3142 24828 3148 24840
rect 3200 24828 3206 24880
rect 5276 24868 5304 24908
rect 5902 24896 5908 24948
rect 5960 24936 5966 24948
rect 9214 24936 9220 24948
rect 5960 24908 9220 24936
rect 5960 24896 5966 24908
rect 9214 24896 9220 24908
rect 9272 24896 9278 24948
rect 11606 24896 11612 24948
rect 11664 24936 11670 24948
rect 12161 24939 12219 24945
rect 12161 24936 12173 24939
rect 11664 24908 12173 24936
rect 11664 24896 11670 24908
rect 12161 24905 12173 24908
rect 12207 24905 12219 24939
rect 12526 24936 12532 24948
rect 12161 24899 12219 24905
rect 12268 24908 12532 24936
rect 5718 24868 5724 24880
rect 5198 24840 5724 24868
rect 5718 24828 5724 24840
rect 5776 24828 5782 24880
rect 6086 24828 6092 24880
rect 6144 24868 6150 24880
rect 6365 24871 6423 24877
rect 6365 24868 6377 24871
rect 6144 24840 6377 24868
rect 6144 24828 6150 24840
rect 6365 24837 6377 24840
rect 6411 24868 6423 24871
rect 8018 24868 8024 24880
rect 6411 24840 8024 24868
rect 6411 24837 6423 24840
rect 6365 24831 6423 24837
rect 2866 24760 2872 24812
rect 2924 24800 2930 24812
rect 3697 24803 3755 24809
rect 3697 24800 3709 24803
rect 2924 24772 3709 24800
rect 2924 24760 2930 24772
rect 3697 24769 3709 24772
rect 3743 24769 3755 24803
rect 3697 24763 3755 24769
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24800 6607 24803
rect 6730 24800 6736 24812
rect 6595 24772 6736 24800
rect 6595 24769 6607 24772
rect 6549 24763 6607 24769
rect 6730 24760 6736 24772
rect 6788 24760 6794 24812
rect 6932 24809 6960 24840
rect 8018 24828 8024 24840
rect 8076 24828 8082 24880
rect 8389 24871 8447 24877
rect 8389 24837 8401 24871
rect 8435 24868 8447 24871
rect 9306 24868 9312 24880
rect 8435 24840 9312 24868
rect 8435 24837 8447 24840
rect 8389 24831 8447 24837
rect 6917 24803 6975 24809
rect 6917 24769 6929 24803
rect 6963 24769 6975 24803
rect 6917 24763 6975 24769
rect 7006 24760 7012 24812
rect 7064 24760 7070 24812
rect 7101 24803 7159 24809
rect 7101 24769 7113 24803
rect 7147 24800 7159 24803
rect 7282 24800 7288 24812
rect 7147 24772 7288 24800
rect 7147 24769 7159 24772
rect 7101 24763 7159 24769
rect 7282 24760 7288 24772
rect 7340 24760 7346 24812
rect 8573 24803 8631 24809
rect 8573 24769 8585 24803
rect 8619 24769 8631 24803
rect 8573 24763 8631 24769
rect 8665 24803 8723 24809
rect 8665 24769 8677 24803
rect 8711 24800 8723 24803
rect 9030 24800 9036 24812
rect 8711 24772 9036 24800
rect 8711 24769 8723 24772
rect 8665 24763 8723 24769
rect 2777 24735 2835 24741
rect 2777 24701 2789 24735
rect 2823 24732 2835 24735
rect 3050 24732 3056 24744
rect 2823 24704 3056 24732
rect 2823 24701 2835 24704
rect 2777 24695 2835 24701
rect 3050 24692 3056 24704
rect 3108 24692 3114 24744
rect 3970 24692 3976 24744
rect 4028 24692 4034 24744
rect 6181 24735 6239 24741
rect 6181 24701 6193 24735
rect 6227 24701 6239 24735
rect 8478 24732 8484 24744
rect 6181 24695 6239 24701
rect 7024 24704 8484 24732
rect 5445 24667 5503 24673
rect 5445 24633 5457 24667
rect 5491 24664 5503 24667
rect 6196 24664 6224 24695
rect 7024 24676 7052 24704
rect 8478 24692 8484 24704
rect 8536 24692 8542 24744
rect 8588 24676 8616 24763
rect 9030 24760 9036 24772
rect 9088 24760 9094 24812
rect 9140 24809 9168 24840
rect 9306 24828 9312 24840
rect 9364 24868 9370 24880
rect 10594 24868 10600 24880
rect 9364 24840 10600 24868
rect 9364 24828 9370 24840
rect 10594 24828 10600 24840
rect 10652 24868 10658 24880
rect 12268 24868 12296 24908
rect 12526 24896 12532 24908
rect 12584 24896 12590 24948
rect 16298 24896 16304 24948
rect 16356 24896 16362 24948
rect 21450 24896 21456 24948
rect 21508 24936 21514 24948
rect 21818 24936 21824 24948
rect 21508 24908 21824 24936
rect 21508 24896 21514 24908
rect 21818 24896 21824 24908
rect 21876 24896 21882 24948
rect 22738 24896 22744 24948
rect 22796 24896 22802 24948
rect 24026 24896 24032 24948
rect 24084 24936 24090 24948
rect 25682 24936 25688 24948
rect 24084 24908 25688 24936
rect 24084 24896 24090 24908
rect 25682 24896 25688 24908
rect 25740 24896 25746 24948
rect 25866 24896 25872 24948
rect 25924 24896 25930 24948
rect 27982 24896 27988 24948
rect 28040 24936 28046 24948
rect 28721 24939 28779 24945
rect 28721 24936 28733 24939
rect 28040 24908 28733 24936
rect 28040 24896 28046 24908
rect 28721 24905 28733 24908
rect 28767 24905 28779 24939
rect 29362 24936 29368 24948
rect 28721 24899 28779 24905
rect 28828 24908 29368 24936
rect 13354 24868 13360 24880
rect 10652 24840 12296 24868
rect 12452 24840 13360 24868
rect 10652 24828 10658 24840
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24769 9183 24803
rect 9125 24763 9183 24769
rect 9218 24803 9276 24809
rect 9218 24769 9230 24803
rect 9264 24769 9276 24803
rect 9218 24763 9276 24769
rect 8846 24692 8852 24744
rect 8904 24732 8910 24744
rect 9233 24732 9261 24763
rect 9398 24760 9404 24812
rect 9456 24760 9462 24812
rect 9493 24803 9551 24809
rect 9493 24769 9505 24803
rect 9539 24769 9551 24803
rect 9493 24763 9551 24769
rect 8904 24704 9261 24732
rect 9508 24732 9536 24763
rect 9582 24760 9588 24812
rect 9640 24809 9646 24812
rect 9640 24800 9648 24809
rect 9640 24772 9685 24800
rect 9640 24763 9648 24772
rect 9640 24760 9646 24763
rect 11146 24760 11152 24812
rect 11204 24760 11210 24812
rect 11330 24760 11336 24812
rect 11388 24760 11394 24812
rect 11532 24809 11560 24840
rect 11517 24803 11575 24809
rect 11517 24769 11529 24803
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 11610 24803 11668 24809
rect 11610 24769 11622 24803
rect 11656 24769 11668 24803
rect 11610 24763 11668 24769
rect 9950 24732 9956 24744
rect 9508 24704 9956 24732
rect 8904 24692 8910 24704
rect 9950 24692 9956 24704
rect 10008 24692 10014 24744
rect 11625 24732 11653 24763
rect 11790 24760 11796 24812
rect 11848 24760 11854 24812
rect 12066 24809 12072 24812
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24769 11943 24803
rect 11885 24763 11943 24769
rect 12023 24803 12072 24809
rect 12023 24769 12035 24803
rect 12069 24769 12072 24803
rect 12023 24763 12072 24769
rect 11164 24704 11653 24732
rect 11900 24732 11928 24763
rect 12066 24760 12072 24763
rect 12124 24760 12130 24812
rect 12250 24760 12256 24812
rect 12308 24760 12314 24812
rect 12452 24809 12480 24840
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 18506 24868 18512 24880
rect 16316 24840 18512 24868
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24769 12495 24803
rect 12437 24763 12495 24769
rect 12526 24760 12532 24812
rect 12584 24760 12590 24812
rect 12641 24803 12699 24809
rect 12641 24769 12653 24803
rect 12687 24800 12699 24803
rect 12687 24772 12757 24800
rect 12687 24769 12699 24772
rect 12641 24763 12699 24769
rect 12729 24732 12757 24772
rect 12802 24760 12808 24812
rect 12860 24760 12866 24812
rect 12894 24760 12900 24812
rect 12952 24800 12958 24812
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12952 24772 13001 24800
rect 12952 24760 12958 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13078 24760 13084 24812
rect 13136 24760 13142 24812
rect 14274 24760 14280 24812
rect 14332 24800 14338 24812
rect 16316 24809 16344 24840
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 14332 24772 16313 24800
rect 14332 24760 14338 24772
rect 16301 24769 16313 24772
rect 16347 24769 16359 24803
rect 16301 24763 16359 24769
rect 16485 24803 16543 24809
rect 16485 24769 16497 24803
rect 16531 24769 16543 24803
rect 16485 24763 16543 24769
rect 13170 24732 13176 24744
rect 11900 24704 12664 24732
rect 12729 24704 13176 24732
rect 7006 24664 7012 24676
rect 5491 24636 7012 24664
rect 5491 24633 5503 24636
rect 5445 24627 5503 24633
rect 7006 24624 7012 24636
rect 7064 24624 7070 24676
rect 8202 24624 8208 24676
rect 8260 24664 8266 24676
rect 8389 24667 8447 24673
rect 8389 24664 8401 24667
rect 8260 24636 8401 24664
rect 8260 24624 8266 24636
rect 8389 24633 8401 24636
rect 8435 24633 8447 24667
rect 8389 24627 8447 24633
rect 8570 24624 8576 24676
rect 8628 24664 8634 24676
rect 10870 24664 10876 24676
rect 8628 24636 10876 24664
rect 8628 24624 8634 24636
rect 10870 24624 10876 24636
rect 10928 24624 10934 24676
rect 11164 24608 11192 24704
rect 12253 24667 12311 24673
rect 12253 24633 12265 24667
rect 12299 24664 12311 24667
rect 12434 24664 12440 24676
rect 12299 24636 12440 24664
rect 12299 24633 12311 24636
rect 12253 24627 12311 24633
rect 12434 24624 12440 24636
rect 12492 24624 12498 24676
rect 12636 24664 12664 24704
rect 13170 24692 13176 24704
rect 13228 24732 13234 24744
rect 14826 24732 14832 24744
rect 13228 24704 14832 24732
rect 13228 24692 13234 24704
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 16500 24732 16528 24763
rect 16666 24760 16672 24812
rect 16724 24800 16730 24812
rect 17236 24809 17264 24840
rect 18506 24828 18512 24840
rect 18564 24828 18570 24880
rect 18598 24828 18604 24880
rect 18656 24868 18662 24880
rect 18656 24840 19288 24868
rect 18656 24828 18662 24840
rect 17129 24803 17187 24809
rect 17129 24800 17141 24803
rect 16724 24772 17141 24800
rect 16724 24760 16730 24772
rect 17129 24769 17141 24772
rect 17175 24769 17187 24803
rect 17129 24763 17187 24769
rect 17221 24803 17279 24809
rect 17221 24769 17233 24803
rect 17267 24769 17279 24803
rect 17221 24763 17279 24769
rect 17405 24803 17463 24809
rect 17405 24769 17417 24803
rect 17451 24769 17463 24803
rect 17405 24763 17463 24769
rect 17420 24732 17448 24763
rect 17954 24760 17960 24812
rect 18012 24760 18018 24812
rect 18782 24760 18788 24812
rect 18840 24760 18846 24812
rect 18966 24760 18972 24812
rect 19024 24760 19030 24812
rect 19260 24809 19288 24840
rect 20806 24828 20812 24880
rect 20864 24868 20870 24880
rect 22002 24868 22008 24880
rect 20864 24840 22008 24868
rect 20864 24828 20870 24840
rect 22002 24828 22008 24840
rect 22060 24828 22066 24880
rect 25884 24868 25912 24896
rect 25884 24840 26193 24868
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24769 19303 24803
rect 19245 24763 19303 24769
rect 19610 24760 19616 24812
rect 19668 24760 19674 24812
rect 22922 24760 22928 24812
rect 22980 24760 22986 24812
rect 23382 24760 23388 24812
rect 23440 24760 23446 24812
rect 23661 24803 23719 24809
rect 23661 24769 23673 24803
rect 23707 24800 23719 24803
rect 23842 24800 23848 24812
rect 23707 24772 23848 24800
rect 23707 24769 23719 24772
rect 23661 24763 23719 24769
rect 23842 24760 23848 24772
rect 23900 24800 23906 24812
rect 24946 24800 24952 24812
rect 23900 24772 24952 24800
rect 23900 24760 23906 24772
rect 24946 24760 24952 24772
rect 25004 24760 25010 24812
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 25685 24763 25743 24769
rect 25778 24803 25836 24809
rect 25778 24769 25790 24803
rect 25824 24800 25836 24803
rect 25866 24800 25872 24812
rect 25824 24772 25872 24800
rect 25824 24769 25836 24772
rect 25778 24763 25836 24769
rect 17586 24732 17592 24744
rect 16500 24704 17592 24732
rect 17586 24692 17592 24704
rect 17644 24692 17650 24744
rect 17972 24732 18000 24760
rect 18877 24735 18935 24741
rect 18877 24732 18889 24735
rect 17972 24704 18889 24732
rect 18877 24701 18889 24704
rect 18923 24701 18935 24735
rect 18877 24695 18935 24701
rect 23109 24735 23167 24741
rect 23109 24701 23121 24735
rect 23155 24732 23167 24735
rect 23477 24735 23535 24741
rect 23477 24732 23489 24735
rect 23155 24704 23489 24732
rect 23155 24701 23167 24704
rect 23109 24695 23167 24701
rect 23477 24701 23489 24704
rect 23523 24701 23535 24735
rect 23477 24695 23535 24701
rect 23750 24692 23756 24744
rect 23808 24732 23814 24744
rect 23937 24735 23995 24741
rect 23937 24732 23949 24735
rect 23808 24704 23949 24732
rect 23808 24692 23814 24704
rect 23937 24701 23949 24704
rect 23983 24732 23995 24735
rect 24670 24732 24676 24744
rect 23983 24704 24676 24732
rect 23983 24701 23995 24704
rect 23937 24695 23995 24701
rect 24670 24692 24676 24704
rect 24728 24732 24734 24744
rect 25700 24732 25728 24763
rect 25866 24760 25872 24772
rect 25924 24760 25930 24812
rect 25958 24760 25964 24812
rect 26016 24760 26022 24812
rect 26050 24760 26056 24812
rect 26108 24760 26114 24812
rect 26165 24809 26193 24840
rect 27172 24840 27384 24868
rect 26150 24803 26208 24809
rect 26150 24769 26162 24803
rect 26196 24800 26208 24803
rect 26418 24800 26424 24812
rect 26196 24772 26424 24800
rect 26196 24769 26208 24772
rect 26150 24763 26208 24769
rect 26418 24760 26424 24772
rect 26476 24760 26482 24812
rect 26602 24760 26608 24812
rect 26660 24800 26666 24812
rect 27172 24800 27200 24840
rect 26660 24772 27200 24800
rect 26660 24760 26666 24772
rect 27246 24760 27252 24812
rect 27304 24760 27310 24812
rect 27356 24800 27384 24840
rect 27433 24803 27491 24809
rect 27433 24800 27445 24803
rect 27356 24772 27445 24800
rect 27433 24769 27445 24772
rect 27479 24769 27491 24803
rect 27433 24763 27491 24769
rect 27522 24760 27528 24812
rect 27580 24760 27586 24812
rect 27982 24760 27988 24812
rect 28040 24800 28046 24812
rect 28040 24772 28120 24800
rect 28040 24760 28046 24772
rect 28092 24766 28120 24772
rect 28169 24769 28227 24775
rect 28169 24766 28181 24769
rect 26620 24732 26648 24760
rect 28092 24738 28181 24766
rect 28169 24735 28181 24738
rect 28215 24735 28227 24769
rect 28258 24760 28264 24812
rect 28316 24760 28322 24812
rect 28828 24800 28856 24908
rect 29362 24896 29368 24908
rect 29420 24936 29426 24948
rect 29546 24936 29552 24948
rect 29420 24908 29552 24936
rect 29420 24896 29426 24908
rect 29546 24896 29552 24908
rect 29604 24896 29610 24948
rect 32030 24896 32036 24948
rect 32088 24936 32094 24948
rect 32582 24936 32588 24948
rect 32088 24908 32588 24936
rect 32088 24896 32094 24908
rect 32582 24896 32588 24908
rect 32640 24896 32646 24948
rect 35897 24939 35955 24945
rect 35897 24905 35909 24939
rect 35943 24936 35955 24939
rect 35986 24936 35992 24948
rect 35943 24908 35992 24936
rect 35943 24905 35955 24908
rect 35897 24899 35955 24905
rect 35986 24896 35992 24908
rect 36044 24896 36050 24948
rect 28902 24828 28908 24880
rect 28960 24868 28966 24880
rect 29638 24868 29644 24880
rect 28960 24840 29644 24868
rect 28960 24828 28966 24840
rect 29638 24828 29644 24840
rect 29696 24828 29702 24880
rect 34146 24868 34152 24880
rect 30300 24840 34152 24868
rect 28997 24803 29055 24809
rect 28997 24800 29009 24803
rect 28828 24772 29009 24800
rect 28997 24769 29009 24772
rect 29043 24769 29055 24803
rect 28997 24763 29055 24769
rect 29135 24803 29193 24809
rect 29135 24769 29147 24803
rect 29181 24800 29193 24803
rect 30300 24800 30328 24840
rect 34146 24828 34152 24840
rect 34204 24828 34210 24880
rect 33873 24803 33931 24809
rect 33873 24800 33885 24803
rect 29181 24772 30328 24800
rect 30392 24772 33885 24800
rect 29181 24769 29193 24772
rect 29135 24763 29193 24769
rect 24728 24704 25176 24732
rect 25700 24704 26648 24732
rect 27264 24704 28028 24732
rect 28169 24729 28227 24735
rect 28353 24735 28411 24741
rect 24728 24692 24734 24704
rect 13262 24664 13268 24676
rect 12636 24636 13268 24664
rect 13262 24624 13268 24636
rect 13320 24624 13326 24676
rect 15194 24624 15200 24676
rect 15252 24664 15258 24676
rect 16669 24667 16727 24673
rect 16669 24664 16681 24667
rect 15252 24636 16681 24664
rect 15252 24624 15258 24636
rect 16669 24633 16681 24636
rect 16715 24633 16727 24667
rect 16669 24627 16727 24633
rect 17310 24624 17316 24676
rect 17368 24664 17374 24676
rect 18414 24664 18420 24676
rect 17368 24636 18420 24664
rect 17368 24624 17374 24636
rect 18414 24624 18420 24636
rect 18472 24664 18478 24676
rect 18782 24664 18788 24676
rect 18472 24636 18788 24664
rect 18472 24624 18478 24636
rect 18782 24624 18788 24636
rect 18840 24624 18846 24676
rect 20530 24664 20536 24676
rect 18892 24636 20536 24664
rect 1670 24556 1676 24608
rect 1728 24596 1734 24608
rect 2225 24599 2283 24605
rect 2225 24596 2237 24599
rect 1728 24568 2237 24596
rect 1728 24556 1734 24568
rect 2225 24565 2237 24568
rect 2271 24565 2283 24599
rect 2225 24559 2283 24565
rect 5258 24556 5264 24608
rect 5316 24596 5322 24608
rect 5537 24599 5595 24605
rect 5537 24596 5549 24599
rect 5316 24568 5549 24596
rect 5316 24556 5322 24568
rect 5537 24565 5549 24568
rect 5583 24565 5595 24599
rect 5537 24559 5595 24565
rect 6454 24556 6460 24608
rect 6512 24596 6518 24608
rect 6641 24599 6699 24605
rect 6641 24596 6653 24599
rect 6512 24568 6653 24596
rect 6512 24556 6518 24568
rect 6641 24565 6653 24568
rect 6687 24565 6699 24599
rect 6641 24559 6699 24565
rect 9030 24556 9036 24608
rect 9088 24596 9094 24608
rect 9674 24596 9680 24608
rect 9088 24568 9680 24596
rect 9088 24556 9094 24568
rect 9674 24556 9680 24568
rect 9732 24556 9738 24608
rect 9769 24599 9827 24605
rect 9769 24565 9781 24599
rect 9815 24596 9827 24599
rect 9950 24596 9956 24608
rect 9815 24568 9956 24596
rect 9815 24565 9827 24568
rect 9769 24559 9827 24565
rect 9950 24556 9956 24568
rect 10008 24556 10014 24608
rect 11146 24556 11152 24608
rect 11204 24556 11210 24608
rect 11330 24556 11336 24608
rect 11388 24556 11394 24608
rect 12342 24556 12348 24608
rect 12400 24596 12406 24608
rect 12805 24599 12863 24605
rect 12805 24596 12817 24599
rect 12400 24568 12817 24596
rect 12400 24556 12406 24568
rect 12805 24565 12817 24568
rect 12851 24565 12863 24599
rect 12805 24559 12863 24565
rect 16942 24556 16948 24608
rect 17000 24556 17006 24608
rect 17034 24556 17040 24608
rect 17092 24556 17098 24608
rect 17862 24556 17868 24608
rect 17920 24556 17926 24608
rect 17954 24556 17960 24608
rect 18012 24596 18018 24608
rect 18892 24596 18920 24636
rect 20530 24624 20536 24636
rect 20588 24624 20594 24676
rect 25038 24664 25044 24676
rect 22066 24636 25044 24664
rect 18012 24568 18920 24596
rect 18012 24556 18018 24568
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 20254 24596 20260 24608
rect 19484 24568 20260 24596
rect 19484 24556 19490 24568
rect 20254 24556 20260 24568
rect 20312 24596 20318 24608
rect 22066 24596 22094 24636
rect 25038 24624 25044 24636
rect 25096 24624 25102 24676
rect 25148 24664 25176 24704
rect 26234 24664 26240 24676
rect 25148 24636 26240 24664
rect 26234 24624 26240 24636
rect 26292 24624 26298 24676
rect 26329 24667 26387 24673
rect 26329 24633 26341 24667
rect 26375 24664 26387 24667
rect 27154 24664 27160 24676
rect 26375 24636 27160 24664
rect 26375 24633 26387 24636
rect 26329 24627 26387 24633
rect 27154 24624 27160 24636
rect 27212 24624 27218 24676
rect 20312 24568 22094 24596
rect 23293 24599 23351 24605
rect 20312 24556 20318 24568
rect 23293 24565 23305 24599
rect 23339 24596 23351 24599
rect 23566 24596 23572 24608
rect 23339 24568 23572 24596
rect 23339 24565 23351 24568
rect 23293 24559 23351 24565
rect 23566 24556 23572 24568
rect 23624 24596 23630 24608
rect 23750 24596 23756 24608
rect 23624 24568 23756 24596
rect 23624 24556 23630 24568
rect 23750 24556 23756 24568
rect 23808 24556 23814 24608
rect 23845 24599 23903 24605
rect 23845 24565 23857 24599
rect 23891 24596 23903 24599
rect 24210 24596 24216 24608
rect 23891 24568 24216 24596
rect 23891 24565 23903 24568
rect 23845 24559 23903 24565
rect 24210 24556 24216 24568
rect 24268 24556 24274 24608
rect 25130 24556 25136 24608
rect 25188 24596 25194 24608
rect 27264 24596 27292 24704
rect 27706 24624 27712 24676
rect 27764 24624 27770 24676
rect 28000 24664 28028 24704
rect 28353 24701 28365 24735
rect 28399 24701 28411 24735
rect 28353 24695 28411 24701
rect 28445 24735 28503 24741
rect 28445 24701 28457 24735
rect 28491 24701 28503 24735
rect 28445 24695 28503 24701
rect 28368 24664 28396 24695
rect 28000 24636 28396 24664
rect 25188 24568 27292 24596
rect 27525 24599 27583 24605
rect 25188 24556 25194 24568
rect 27525 24565 27537 24599
rect 27571 24596 27583 24599
rect 27890 24596 27896 24608
rect 27571 24568 27896 24596
rect 27571 24565 27583 24568
rect 27525 24559 27583 24565
rect 27890 24556 27896 24568
rect 27948 24556 27954 24608
rect 28258 24556 28264 24608
rect 28316 24596 28322 24608
rect 28460 24596 28488 24695
rect 28810 24692 28816 24744
rect 28868 24732 28874 24744
rect 28905 24735 28963 24741
rect 28905 24732 28917 24735
rect 28868 24704 28917 24732
rect 28868 24692 28874 24704
rect 28905 24701 28917 24704
rect 28951 24701 28963 24735
rect 28905 24695 28963 24701
rect 29270 24692 29276 24744
rect 29328 24692 29334 24744
rect 29365 24735 29423 24741
rect 29365 24701 29377 24735
rect 29411 24732 29423 24735
rect 29638 24732 29644 24744
rect 29411 24704 29644 24732
rect 29411 24701 29423 24704
rect 29365 24695 29423 24701
rect 29638 24692 29644 24704
rect 29696 24692 29702 24744
rect 29822 24692 29828 24744
rect 29880 24732 29886 24744
rect 30392 24732 30420 24772
rect 33873 24769 33885 24772
rect 33919 24769 33931 24803
rect 33873 24763 33931 24769
rect 34057 24803 34115 24809
rect 34057 24769 34069 24803
rect 34103 24800 34115 24803
rect 34330 24800 34336 24812
rect 34103 24772 34336 24800
rect 34103 24769 34115 24772
rect 34057 24763 34115 24769
rect 34330 24760 34336 24772
rect 34388 24760 34394 24812
rect 35161 24803 35219 24809
rect 35161 24769 35173 24803
rect 35207 24800 35219 24803
rect 35250 24800 35256 24812
rect 35207 24772 35256 24800
rect 35207 24769 35219 24772
rect 35161 24763 35219 24769
rect 35250 24760 35256 24772
rect 35308 24760 35314 24812
rect 35345 24803 35403 24809
rect 35345 24769 35357 24803
rect 35391 24769 35403 24803
rect 35345 24763 35403 24769
rect 29880 24704 30420 24732
rect 29880 24692 29886 24704
rect 30650 24692 30656 24744
rect 30708 24732 30714 24744
rect 31938 24732 31944 24744
rect 30708 24704 31944 24732
rect 30708 24692 30714 24704
rect 31938 24692 31944 24704
rect 31996 24692 32002 24744
rect 28629 24667 28687 24673
rect 28629 24633 28641 24667
rect 28675 24664 28687 24667
rect 28675 24636 30052 24664
rect 28675 24633 28687 24636
rect 28629 24627 28687 24633
rect 28316 24568 28488 24596
rect 28316 24556 28322 24568
rect 28718 24556 28724 24608
rect 28776 24596 28782 24608
rect 29822 24596 29828 24608
rect 28776 24568 29828 24596
rect 28776 24556 28782 24568
rect 29822 24556 29828 24568
rect 29880 24556 29886 24608
rect 30024 24596 30052 24636
rect 30282 24624 30288 24676
rect 30340 24664 30346 24676
rect 35360 24664 35388 24763
rect 35986 24760 35992 24812
rect 36044 24760 36050 24812
rect 30340 24636 35388 24664
rect 30340 24624 30346 24636
rect 33686 24596 33692 24608
rect 30024 24568 33692 24596
rect 33686 24556 33692 24568
rect 33744 24596 33750 24608
rect 33873 24599 33931 24605
rect 33873 24596 33885 24599
rect 33744 24568 33885 24596
rect 33744 24556 33750 24568
rect 33873 24565 33885 24568
rect 33919 24565 33931 24599
rect 33873 24559 33931 24565
rect 34146 24556 34152 24608
rect 34204 24596 34210 24608
rect 34241 24599 34299 24605
rect 34241 24596 34253 24599
rect 34204 24568 34253 24596
rect 34204 24556 34210 24568
rect 34241 24565 34253 24568
rect 34287 24565 34299 24599
rect 34241 24559 34299 24565
rect 34330 24556 34336 24608
rect 34388 24596 34394 24608
rect 35529 24599 35587 24605
rect 35529 24596 35541 24599
rect 34388 24568 35541 24596
rect 34388 24556 34394 24568
rect 35529 24565 35541 24568
rect 35575 24596 35587 24599
rect 35894 24596 35900 24608
rect 35575 24568 35900 24596
rect 35575 24565 35587 24568
rect 35529 24559 35587 24565
rect 35894 24556 35900 24568
rect 35952 24556 35958 24608
rect 1104 24506 36432 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 36432 24506
rect 1104 24432 36432 24454
rect 3142 24352 3148 24404
rect 3200 24392 3206 24404
rect 3602 24392 3608 24404
rect 3200 24364 3608 24392
rect 3200 24352 3206 24364
rect 3602 24352 3608 24364
rect 3660 24352 3666 24404
rect 3970 24352 3976 24404
rect 4028 24392 4034 24404
rect 4801 24395 4859 24401
rect 4801 24392 4813 24395
rect 4028 24364 4813 24392
rect 4028 24352 4034 24364
rect 4801 24361 4813 24364
rect 4847 24361 4859 24395
rect 5721 24395 5779 24401
rect 4801 24355 4859 24361
rect 5184 24364 5672 24392
rect 5184 24324 5212 24364
rect 4816 24296 5212 24324
rect 5644 24324 5672 24364
rect 5721 24361 5733 24395
rect 5767 24392 5779 24395
rect 5810 24392 5816 24404
rect 5767 24364 5816 24392
rect 5767 24361 5779 24364
rect 5721 24355 5779 24361
rect 5810 24352 5816 24364
rect 5868 24352 5874 24404
rect 6914 24392 6920 24404
rect 6104 24364 6920 24392
rect 6104 24324 6132 24364
rect 6914 24352 6920 24364
rect 6972 24352 6978 24404
rect 10962 24352 10968 24404
rect 11020 24392 11026 24404
rect 11609 24395 11667 24401
rect 11609 24392 11621 24395
rect 11020 24364 11621 24392
rect 11020 24352 11026 24364
rect 11609 24361 11621 24364
rect 11655 24361 11667 24395
rect 12618 24392 12624 24404
rect 11609 24355 11667 24361
rect 12360 24364 12624 24392
rect 5644 24296 6132 24324
rect 4816 24268 4844 24296
rect 6178 24284 6184 24336
rect 6236 24324 6242 24336
rect 6641 24327 6699 24333
rect 6641 24324 6653 24327
rect 6236 24296 6653 24324
rect 6236 24284 6242 24296
rect 6641 24293 6653 24296
rect 6687 24293 6699 24327
rect 6641 24287 6699 24293
rect 7282 24284 7288 24336
rect 7340 24284 7346 24336
rect 9309 24327 9367 24333
rect 9309 24324 9321 24327
rect 7391 24296 9321 24324
rect 1670 24216 1676 24268
rect 1728 24216 1734 24268
rect 4798 24216 4804 24268
rect 4856 24216 4862 24268
rect 5258 24216 5264 24268
rect 5316 24216 5322 24268
rect 5442 24216 5448 24268
rect 5500 24216 5506 24268
rect 7391 24256 7419 24296
rect 9309 24293 9321 24296
rect 9355 24293 9367 24327
rect 9309 24287 9367 24293
rect 10042 24284 10048 24336
rect 10100 24324 10106 24336
rect 10100 24296 11652 24324
rect 10100 24284 10106 24296
rect 7300 24228 7419 24256
rect 8205 24259 8263 24265
rect 1394 24148 1400 24200
rect 1452 24148 1458 24200
rect 2774 24148 2780 24200
rect 2832 24148 2838 24200
rect 6362 24148 6368 24200
rect 6420 24188 6426 24200
rect 6825 24191 6883 24197
rect 6825 24188 6837 24191
rect 6420 24160 6837 24188
rect 6420 24148 6426 24160
rect 6825 24157 6837 24160
rect 6871 24157 6883 24191
rect 6825 24151 6883 24157
rect 6917 24191 6975 24197
rect 6917 24157 6929 24191
rect 6963 24188 6975 24191
rect 7009 24191 7067 24197
rect 7009 24188 7021 24191
rect 6963 24160 7021 24188
rect 6963 24157 6975 24160
rect 6917 24151 6975 24157
rect 7009 24157 7021 24160
rect 7055 24188 7067 24191
rect 7190 24188 7196 24200
rect 7055 24160 7196 24188
rect 7055 24157 7067 24160
rect 7009 24151 7067 24157
rect 7190 24148 7196 24160
rect 7248 24148 7254 24200
rect 7300 24197 7328 24228
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8294 24256 8300 24268
rect 8251 24228 8300 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8294 24216 8300 24228
rect 8352 24216 8358 24268
rect 10239 24256 10267 24296
rect 10870 24256 10876 24268
rect 9600 24228 10267 24256
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 7374 24148 7380 24200
rect 7432 24148 7438 24200
rect 9488 24191 9546 24197
rect 9488 24157 9500 24191
rect 9534 24188 9546 24191
rect 9600 24188 9628 24228
rect 9534 24160 9628 24188
rect 9534 24157 9546 24160
rect 9488 24151 9546 24157
rect 9766 24148 9772 24200
rect 9824 24197 9830 24200
rect 9824 24191 9863 24197
rect 9851 24157 9863 24191
rect 9824 24151 9863 24157
rect 9824 24148 9830 24151
rect 9950 24148 9956 24200
rect 10008 24148 10014 24200
rect 10239 24197 10267 24228
rect 10336 24228 10876 24256
rect 10336 24197 10364 24228
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11514 24256 11520 24268
rect 11072 24228 11520 24256
rect 10224 24191 10282 24197
rect 10224 24157 10236 24191
rect 10270 24157 10282 24191
rect 10224 24151 10282 24157
rect 10321 24191 10379 24197
rect 10321 24157 10333 24191
rect 10367 24157 10379 24191
rect 10321 24151 10379 24157
rect 10502 24148 10508 24200
rect 10560 24197 10566 24200
rect 10560 24191 10599 24197
rect 10587 24157 10599 24191
rect 10560 24151 10599 24157
rect 10560 24148 10566 24151
rect 10686 24148 10692 24200
rect 10744 24148 10750 24200
rect 11072 24197 11100 24228
rect 11514 24216 11520 24228
rect 11572 24216 11578 24268
rect 11057 24191 11115 24197
rect 11057 24157 11069 24191
rect 11103 24157 11115 24191
rect 11057 24151 11115 24157
rect 11241 24191 11299 24197
rect 11241 24157 11253 24191
rect 11287 24157 11299 24191
rect 11241 24151 11299 24157
rect 11425 24191 11483 24197
rect 11425 24157 11437 24191
rect 11471 24188 11483 24191
rect 11624 24188 11652 24296
rect 11974 24284 11980 24336
rect 12032 24324 12038 24336
rect 12360 24333 12388 24364
rect 12618 24352 12624 24364
rect 12676 24352 12682 24404
rect 13262 24352 13268 24404
rect 13320 24392 13326 24404
rect 13320 24364 13584 24392
rect 13320 24352 13326 24364
rect 12161 24327 12219 24333
rect 12161 24324 12173 24327
rect 12032 24296 12173 24324
rect 12032 24284 12038 24296
rect 12161 24293 12173 24296
rect 12207 24293 12219 24327
rect 12161 24287 12219 24293
rect 12345 24327 12403 24333
rect 12345 24293 12357 24327
rect 12391 24293 12403 24327
rect 12345 24287 12403 24293
rect 13170 24284 13176 24336
rect 13228 24324 13234 24336
rect 13556 24324 13584 24364
rect 13722 24352 13728 24404
rect 13780 24392 13786 24404
rect 14277 24395 14335 24401
rect 14277 24392 14289 24395
rect 13780 24364 14289 24392
rect 13780 24352 13786 24364
rect 14277 24361 14289 24364
rect 14323 24361 14335 24395
rect 14277 24355 14335 24361
rect 14458 24352 14464 24404
rect 14516 24392 14522 24404
rect 14921 24395 14979 24401
rect 14921 24392 14933 24395
rect 14516 24364 14933 24392
rect 14516 24352 14522 24364
rect 14921 24361 14933 24364
rect 14967 24361 14979 24395
rect 14921 24355 14979 24361
rect 17129 24395 17187 24401
rect 17129 24361 17141 24395
rect 17175 24392 17187 24395
rect 17862 24392 17868 24404
rect 17175 24364 17868 24392
rect 17175 24361 17187 24364
rect 17129 24355 17187 24361
rect 17862 24352 17868 24364
rect 17920 24352 17926 24404
rect 18969 24395 19027 24401
rect 18969 24361 18981 24395
rect 19015 24392 19027 24395
rect 19150 24392 19156 24404
rect 19015 24364 19156 24392
rect 19015 24361 19027 24364
rect 18969 24355 19027 24361
rect 19150 24352 19156 24364
rect 19208 24352 19214 24404
rect 19794 24352 19800 24404
rect 19852 24392 19858 24404
rect 20073 24395 20131 24401
rect 20073 24392 20085 24395
rect 19852 24364 20085 24392
rect 19852 24352 19858 24364
rect 20073 24361 20085 24364
rect 20119 24361 20131 24395
rect 20073 24355 20131 24361
rect 20530 24352 20536 24404
rect 20588 24392 20594 24404
rect 20625 24395 20683 24401
rect 20625 24392 20637 24395
rect 20588 24364 20637 24392
rect 20588 24352 20594 24364
rect 20625 24361 20637 24364
rect 20671 24361 20683 24395
rect 20625 24355 20683 24361
rect 20990 24352 20996 24404
rect 21048 24392 21054 24404
rect 21085 24395 21143 24401
rect 21085 24392 21097 24395
rect 21048 24364 21097 24392
rect 21048 24352 21054 24364
rect 21085 24361 21097 24364
rect 21131 24361 21143 24395
rect 21085 24355 21143 24361
rect 21358 24352 21364 24404
rect 21416 24392 21422 24404
rect 24026 24392 24032 24404
rect 21416 24364 24032 24392
rect 21416 24352 21422 24364
rect 24026 24352 24032 24364
rect 24084 24352 24090 24404
rect 25317 24395 25375 24401
rect 25317 24361 25329 24395
rect 25363 24392 25375 24395
rect 26050 24392 26056 24404
rect 25363 24364 26056 24392
rect 25363 24361 25375 24364
rect 25317 24355 25375 24361
rect 26050 24352 26056 24364
rect 26108 24352 26114 24404
rect 26234 24352 26240 24404
rect 26292 24392 26298 24404
rect 26510 24392 26516 24404
rect 26292 24364 26516 24392
rect 26292 24352 26298 24364
rect 26510 24352 26516 24364
rect 26568 24352 26574 24404
rect 26602 24352 26608 24404
rect 26660 24352 26666 24404
rect 26970 24392 26976 24404
rect 26804 24364 26976 24392
rect 16022 24324 16028 24336
rect 13228 24296 13491 24324
rect 13556 24296 14504 24324
rect 13228 24284 13234 24296
rect 12268 24228 13308 24256
rect 11974 24188 11980 24200
rect 11471 24160 11980 24188
rect 11471 24157 11483 24160
rect 11425 24151 11483 24157
rect 5169 24123 5227 24129
rect 5169 24089 5181 24123
rect 5215 24120 5227 24123
rect 5350 24120 5356 24132
rect 5215 24092 5356 24120
rect 5215 24089 5227 24092
rect 5169 24083 5227 24089
rect 5350 24080 5356 24092
rect 5408 24120 5414 24132
rect 5534 24120 5540 24132
rect 5408 24092 5540 24120
rect 5408 24080 5414 24092
rect 5534 24080 5540 24092
rect 5592 24080 5598 24132
rect 5810 24080 5816 24132
rect 5868 24080 5874 24132
rect 5994 24080 6000 24132
rect 6052 24080 6058 24132
rect 6270 24080 6276 24132
rect 6328 24120 6334 24132
rect 6546 24120 6552 24132
rect 6328 24092 6552 24120
rect 6328 24080 6334 24092
rect 6546 24080 6552 24092
rect 6604 24080 6610 24132
rect 6641 24123 6699 24129
rect 6641 24089 6653 24123
rect 6687 24120 6699 24123
rect 6687 24092 7420 24120
rect 6687 24089 6699 24092
rect 6641 24083 6699 24089
rect 6914 24012 6920 24064
rect 6972 24052 6978 24064
rect 7101 24055 7159 24061
rect 7101 24052 7113 24055
rect 6972 24024 7113 24052
rect 6972 24012 6978 24024
rect 7101 24021 7113 24024
rect 7147 24021 7159 24055
rect 7392 24052 7420 24092
rect 8220 24092 9444 24120
rect 8220 24052 8248 24092
rect 7392 24024 8248 24052
rect 9416 24052 9444 24092
rect 9582 24080 9588 24132
rect 9640 24080 9646 24132
rect 9674 24080 9680 24132
rect 9732 24120 9738 24132
rect 10413 24123 10471 24129
rect 10413 24120 10425 24123
rect 9732 24092 10425 24120
rect 9732 24080 9738 24092
rect 10413 24089 10425 24092
rect 10459 24120 10471 24123
rect 11256 24120 11284 24151
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 10459 24092 11284 24120
rect 10459 24089 10471 24092
rect 10413 24083 10471 24089
rect 10045 24055 10103 24061
rect 10045 24052 10057 24055
rect 9416 24024 10057 24052
rect 7101 24015 7159 24021
rect 10045 24021 10057 24024
rect 10091 24021 10103 24055
rect 11256 24052 11284 24092
rect 11330 24080 11336 24132
rect 11388 24080 11394 24132
rect 12268 24120 12296 24228
rect 13280 24200 13308 24228
rect 12986 24148 12992 24200
rect 13044 24148 13050 24200
rect 13078 24148 13084 24200
rect 13136 24188 13142 24200
rect 13136 24160 13181 24188
rect 13136 24148 13142 24160
rect 13262 24148 13268 24200
rect 13320 24148 13326 24200
rect 13463 24197 13491 24296
rect 14476 24256 14504 24296
rect 15028 24296 16028 24324
rect 15028 24265 15056 24296
rect 16022 24284 16028 24296
rect 16080 24324 16086 24336
rect 16080 24296 17356 24324
rect 16080 24284 16086 24296
rect 15013 24259 15071 24265
rect 14476 24228 14964 24256
rect 14476 24197 14504 24228
rect 13454 24191 13512 24197
rect 13454 24157 13466 24191
rect 13500 24157 13512 24191
rect 13454 24151 13512 24157
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24188 14611 24191
rect 14734 24188 14740 24200
rect 14599 24160 14740 24188
rect 14599 24157 14611 24160
rect 14553 24151 14611 24157
rect 14734 24148 14740 24160
rect 14792 24148 14798 24200
rect 14826 24148 14832 24200
rect 14884 24148 14890 24200
rect 14936 24188 14964 24228
rect 15013 24225 15025 24259
rect 15059 24225 15071 24259
rect 15013 24219 15071 24225
rect 15105 24259 15163 24265
rect 15105 24225 15117 24259
rect 15151 24256 15163 24259
rect 16482 24256 16488 24268
rect 15151 24228 16488 24256
rect 15151 24225 15163 24228
rect 15105 24219 15163 24225
rect 16482 24216 16488 24228
rect 16540 24256 16546 24268
rect 17328 24265 17356 24296
rect 17586 24284 17592 24336
rect 17644 24284 17650 24336
rect 17770 24284 17776 24336
rect 17828 24324 17834 24336
rect 20898 24324 20904 24336
rect 17828 24296 19748 24324
rect 17828 24284 17834 24296
rect 17221 24259 17279 24265
rect 17221 24256 17233 24259
rect 16540 24228 17233 24256
rect 16540 24216 16546 24228
rect 17221 24225 17233 24228
rect 17267 24225 17279 24259
rect 17221 24219 17279 24225
rect 17313 24259 17371 24265
rect 17313 24225 17325 24259
rect 17359 24256 17371 24259
rect 17954 24256 17960 24268
rect 17359 24228 17960 24256
rect 17359 24225 17371 24228
rect 17313 24219 17371 24225
rect 17954 24216 17960 24228
rect 18012 24216 18018 24268
rect 18046 24216 18052 24268
rect 18104 24256 18110 24268
rect 18104 24228 19012 24256
rect 18104 24216 18110 24228
rect 18984 24200 19012 24228
rect 15838 24188 15844 24200
rect 14936 24160 15844 24188
rect 15838 24148 15844 24160
rect 15896 24148 15902 24200
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 16899 24160 18644 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 11440 24092 12296 24120
rect 11440 24052 11468 24092
rect 12618 24080 12624 24132
rect 12676 24080 12682 24132
rect 13377 24123 13435 24129
rect 13377 24089 13389 24123
rect 13423 24120 13435 24123
rect 13722 24120 13728 24132
rect 13423 24092 13728 24120
rect 13423 24089 13435 24092
rect 13377 24083 13435 24089
rect 13722 24080 13728 24092
rect 13780 24080 13786 24132
rect 14642 24080 14648 24132
rect 14700 24080 14706 24132
rect 15010 24080 15016 24132
rect 15068 24120 15074 24132
rect 15381 24123 15439 24129
rect 15381 24120 15393 24123
rect 15068 24092 15393 24120
rect 15068 24080 15074 24092
rect 15381 24089 15393 24092
rect 15427 24120 15439 24123
rect 16868 24120 16896 24151
rect 15427 24092 16896 24120
rect 15427 24089 15439 24092
rect 15381 24083 15439 24089
rect 17218 24080 17224 24132
rect 17276 24120 17282 24132
rect 17770 24120 17776 24132
rect 17276 24092 17776 24120
rect 17276 24080 17282 24092
rect 17770 24080 17776 24092
rect 17828 24080 17834 24132
rect 18616 24120 18644 24160
rect 18782 24148 18788 24200
rect 18840 24148 18846 24200
rect 18966 24148 18972 24200
rect 19024 24148 19030 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19444 24120 19472 24151
rect 19518 24148 19524 24200
rect 19576 24148 19582 24200
rect 19720 24188 19748 24296
rect 19812 24296 20904 24324
rect 19812 24265 19840 24296
rect 20898 24284 20904 24296
rect 20956 24284 20962 24336
rect 21177 24327 21235 24333
rect 21177 24293 21189 24327
rect 21223 24324 21235 24327
rect 21818 24324 21824 24336
rect 21223 24296 21824 24324
rect 21223 24293 21235 24296
rect 21177 24287 21235 24293
rect 19797 24259 19855 24265
rect 19797 24225 19809 24259
rect 19843 24225 19855 24259
rect 19797 24219 19855 24225
rect 19886 24216 19892 24268
rect 19944 24216 19950 24268
rect 21192 24256 21220 24287
rect 21818 24284 21824 24296
rect 21876 24284 21882 24336
rect 20364 24228 21220 24256
rect 20364 24197 20392 24228
rect 23382 24216 23388 24268
rect 23440 24256 23446 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 23440 24228 24593 24256
rect 23440 24216 23446 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 26068 24256 26096 24352
rect 26602 24256 26608 24268
rect 24581 24219 24639 24225
rect 24964 24228 26096 24256
rect 26344 24228 26608 24256
rect 20257 24191 20315 24197
rect 20257 24188 20269 24191
rect 19720 24160 20269 24188
rect 20257 24157 20269 24160
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 20349 24191 20407 24197
rect 20349 24157 20361 24191
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 20806 24148 20812 24200
rect 20864 24148 20870 24200
rect 20898 24148 20904 24200
rect 20956 24188 20962 24200
rect 21634 24188 21640 24200
rect 20956 24160 21640 24188
rect 20956 24148 20962 24160
rect 21634 24148 21640 24160
rect 21692 24188 21698 24200
rect 23198 24188 23204 24200
rect 21692 24160 23204 24188
rect 21692 24148 21698 24160
rect 23198 24148 23204 24160
rect 23256 24148 23262 24200
rect 24302 24148 24308 24200
rect 24360 24188 24366 24200
rect 24453 24191 24511 24197
rect 24453 24188 24465 24191
rect 24360 24160 24465 24188
rect 24360 24148 24366 24160
rect 24453 24157 24465 24160
rect 24499 24157 24511 24191
rect 24964 24188 24992 24228
rect 24453 24151 24511 24157
rect 24596 24160 24992 24188
rect 25041 24191 25099 24197
rect 19794 24120 19800 24132
rect 18616 24092 19800 24120
rect 19794 24080 19800 24092
rect 19852 24080 19858 24132
rect 20073 24123 20131 24129
rect 20073 24089 20085 24123
rect 20119 24120 20131 24123
rect 20622 24120 20628 24132
rect 20119 24092 20628 24120
rect 20119 24089 20131 24092
rect 20073 24083 20131 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 21082 24080 21088 24132
rect 21140 24120 21146 24132
rect 21545 24123 21603 24129
rect 21545 24120 21557 24123
rect 21140 24092 21557 24120
rect 21140 24080 21146 24092
rect 21545 24089 21557 24092
rect 21591 24120 21603 24123
rect 23658 24120 23664 24132
rect 21591 24092 23664 24120
rect 21591 24089 21603 24092
rect 21545 24083 21603 24089
rect 23658 24080 23664 24092
rect 23716 24080 23722 24132
rect 24596 24129 24624 24160
rect 25041 24157 25053 24191
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 24581 24123 24639 24129
rect 24581 24089 24593 24123
rect 24627 24089 24639 24123
rect 24581 24083 24639 24089
rect 24673 24123 24731 24129
rect 24673 24089 24685 24123
rect 24719 24089 24731 24123
rect 24673 24083 24731 24089
rect 11256 24024 11468 24052
rect 10045 24015 10103 24021
rect 12250 24012 12256 24064
rect 12308 24052 12314 24064
rect 13633 24055 13691 24061
rect 13633 24052 13645 24055
rect 12308 24024 13645 24052
rect 12308 24012 12314 24024
rect 13633 24021 13645 24024
rect 13679 24021 13691 24055
rect 13633 24015 13691 24021
rect 14090 24012 14096 24064
rect 14148 24052 14154 24064
rect 15289 24055 15347 24061
rect 15289 24052 15301 24055
rect 14148 24024 15301 24052
rect 14148 24012 14154 24024
rect 15289 24021 15301 24024
rect 15335 24052 15347 24055
rect 16945 24055 17003 24061
rect 16945 24052 16957 24055
rect 15335 24024 16957 24052
rect 15335 24021 15347 24024
rect 15289 24015 15347 24021
rect 16945 24021 16957 24024
rect 16991 24021 17003 24055
rect 16945 24015 17003 24021
rect 17586 24012 17592 24064
rect 17644 24052 17650 24064
rect 19150 24052 19156 24064
rect 17644 24024 19156 24052
rect 17644 24012 17650 24024
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 19242 24012 19248 24064
rect 19300 24012 19306 24064
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 20346 24052 20352 24064
rect 19944 24024 20352 24052
rect 19944 24012 19950 24024
rect 20346 24012 20352 24024
rect 20404 24012 20410 24064
rect 20530 24012 20536 24064
rect 20588 24012 20594 24064
rect 21345 24055 21403 24061
rect 21345 24021 21357 24055
rect 21391 24052 21403 24055
rect 21910 24052 21916 24064
rect 21391 24024 21916 24052
rect 21391 24021 21403 24024
rect 21345 24015 21403 24021
rect 21910 24012 21916 24024
rect 21968 24012 21974 24064
rect 24210 24012 24216 24064
rect 24268 24052 24274 24064
rect 24688 24052 24716 24083
rect 24854 24080 24860 24132
rect 24912 24080 24918 24132
rect 25056 24120 25084 24151
rect 25130 24148 25136 24200
rect 25188 24148 25194 24200
rect 25774 24148 25780 24200
rect 25832 24188 25838 24200
rect 25958 24188 25964 24200
rect 25832 24160 25964 24188
rect 25832 24148 25838 24160
rect 25958 24148 25964 24160
rect 26016 24188 26022 24200
rect 26344 24197 26372 24228
rect 26602 24216 26608 24228
rect 26660 24216 26666 24268
rect 26804 24256 26832 24364
rect 26970 24352 26976 24364
rect 27028 24392 27034 24404
rect 27798 24392 27804 24404
rect 27028 24364 27804 24392
rect 27028 24352 27034 24364
rect 27798 24352 27804 24364
rect 27856 24352 27862 24404
rect 27890 24352 27896 24404
rect 27948 24392 27954 24404
rect 28810 24392 28816 24404
rect 27948 24364 28816 24392
rect 27948 24352 27954 24364
rect 28810 24352 28816 24364
rect 28868 24352 28874 24404
rect 31573 24395 31631 24401
rect 31573 24361 31585 24395
rect 31619 24361 31631 24395
rect 31573 24355 31631 24361
rect 27249 24327 27307 24333
rect 27249 24293 27261 24327
rect 27295 24324 27307 24327
rect 27522 24324 27528 24336
rect 27295 24296 27528 24324
rect 27295 24293 27307 24296
rect 27249 24287 27307 24293
rect 27522 24284 27528 24296
rect 27580 24324 27586 24336
rect 30282 24324 30288 24336
rect 27580 24296 30288 24324
rect 27580 24284 27586 24296
rect 30282 24284 30288 24296
rect 30340 24284 30346 24336
rect 30926 24324 30932 24336
rect 30760 24296 30932 24324
rect 26712 24228 26832 24256
rect 27080 24228 27752 24256
rect 26053 24191 26111 24197
rect 26053 24188 26065 24191
rect 26016 24160 26065 24188
rect 26016 24148 26022 24160
rect 26053 24157 26065 24160
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26329 24191 26387 24197
rect 26329 24157 26341 24191
rect 26375 24157 26387 24191
rect 26329 24151 26387 24157
rect 26418 24148 26424 24200
rect 26476 24148 26482 24200
rect 26712 24197 26740 24228
rect 27080 24197 27108 24228
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24157 26755 24191
rect 26973 24191 27031 24197
rect 26973 24188 26985 24191
rect 26697 24151 26755 24157
rect 26804 24160 26985 24188
rect 25222 24120 25228 24132
rect 25056 24092 25228 24120
rect 25222 24080 25228 24092
rect 25280 24080 25286 24132
rect 26234 24080 26240 24132
rect 26292 24080 26298 24132
rect 26804 24120 26832 24160
rect 26973 24157 26985 24160
rect 27019 24157 27031 24191
rect 26973 24151 27031 24157
rect 27065 24191 27123 24197
rect 27065 24157 27077 24191
rect 27111 24157 27123 24191
rect 27065 24151 27123 24157
rect 26436 24092 26832 24120
rect 26436 24064 26464 24092
rect 26878 24080 26884 24132
rect 26936 24080 26942 24132
rect 24268 24024 24716 24052
rect 24268 24012 24274 24024
rect 26418 24012 26424 24064
rect 26476 24012 26482 24064
rect 26510 24012 26516 24064
rect 26568 24052 26574 24064
rect 27080 24052 27108 24151
rect 27154 24148 27160 24200
rect 27212 24188 27218 24200
rect 27341 24191 27399 24197
rect 27341 24188 27353 24191
rect 27212 24160 27353 24188
rect 27212 24148 27218 24160
rect 27341 24157 27353 24160
rect 27387 24157 27399 24191
rect 27341 24151 27399 24157
rect 26568 24024 27108 24052
rect 27356 24052 27384 24151
rect 27522 24148 27528 24200
rect 27580 24148 27586 24200
rect 27724 24197 27752 24228
rect 27798 24216 27804 24268
rect 27856 24256 27862 24268
rect 30006 24256 30012 24268
rect 27856 24228 30012 24256
rect 27856 24216 27862 24228
rect 30006 24216 30012 24228
rect 30064 24216 30070 24268
rect 27709 24191 27767 24197
rect 27709 24157 27721 24191
rect 27755 24188 27767 24191
rect 28258 24188 28264 24200
rect 27755 24160 28264 24188
rect 27755 24157 27767 24160
rect 27709 24151 27767 24157
rect 28258 24148 28264 24160
rect 28316 24148 28322 24200
rect 29270 24148 29276 24200
rect 29328 24188 29334 24200
rect 30650 24188 30656 24200
rect 29328 24160 30656 24188
rect 29328 24148 29334 24160
rect 30650 24148 30656 24160
rect 30708 24148 30714 24200
rect 27614 24080 27620 24132
rect 27672 24080 27678 24132
rect 28166 24080 28172 24132
rect 28224 24120 28230 24132
rect 30760 24120 30788 24296
rect 30926 24284 30932 24296
rect 30984 24284 30990 24336
rect 31588 24324 31616 24355
rect 31754 24352 31760 24404
rect 31812 24352 31818 24404
rect 35897 24395 35955 24401
rect 35897 24361 35909 24395
rect 35943 24392 35955 24395
rect 36170 24392 36176 24404
rect 35943 24364 36176 24392
rect 35943 24361 35955 24364
rect 35897 24355 35955 24361
rect 36170 24352 36176 24364
rect 36228 24352 36234 24404
rect 31846 24324 31852 24336
rect 31588 24296 31852 24324
rect 31846 24284 31852 24296
rect 31904 24284 31910 24336
rect 31481 24259 31539 24265
rect 30852 24228 31432 24256
rect 30852 24197 30880 24228
rect 30837 24191 30895 24197
rect 30837 24157 30849 24191
rect 30883 24157 30895 24191
rect 30837 24151 30895 24157
rect 31018 24148 31024 24200
rect 31076 24148 31082 24200
rect 28224 24092 30788 24120
rect 28224 24080 28230 24092
rect 30926 24080 30932 24132
rect 30984 24080 30990 24132
rect 31294 24080 31300 24132
rect 31352 24080 31358 24132
rect 31404 24120 31432 24228
rect 31481 24225 31493 24259
rect 31527 24256 31539 24259
rect 31754 24256 31760 24268
rect 31527 24228 31760 24256
rect 31527 24225 31539 24228
rect 31481 24219 31539 24225
rect 31754 24216 31760 24228
rect 31812 24216 31818 24268
rect 31570 24148 31576 24200
rect 31628 24148 31634 24200
rect 36078 24148 36084 24200
rect 36136 24148 36142 24200
rect 33410 24120 33416 24132
rect 31404 24092 33416 24120
rect 33410 24080 33416 24092
rect 33468 24080 33474 24132
rect 29270 24052 29276 24064
rect 27356 24024 29276 24052
rect 26568 24012 26574 24024
rect 29270 24012 29276 24024
rect 29328 24012 29334 24064
rect 30834 24012 30840 24064
rect 30892 24052 30898 24064
rect 31205 24055 31263 24061
rect 31205 24052 31217 24055
rect 30892 24024 31217 24052
rect 30892 24012 30898 24024
rect 31205 24021 31217 24024
rect 31251 24052 31263 24055
rect 31570 24052 31576 24064
rect 31251 24024 31576 24052
rect 31251 24021 31263 24024
rect 31205 24015 31263 24021
rect 31570 24012 31576 24024
rect 31628 24012 31634 24064
rect 1104 23962 36432 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 36432 23962
rect 1104 23888 36432 23910
rect 6086 23808 6092 23860
rect 6144 23848 6150 23860
rect 7009 23851 7067 23857
rect 7009 23848 7021 23851
rect 6144 23820 7021 23848
rect 6144 23808 6150 23820
rect 7009 23817 7021 23820
rect 7055 23817 7067 23851
rect 7009 23811 7067 23817
rect 8849 23851 8907 23857
rect 8849 23817 8861 23851
rect 8895 23848 8907 23851
rect 8938 23848 8944 23860
rect 8895 23820 8944 23848
rect 8895 23817 8907 23820
rect 8849 23811 8907 23817
rect 8938 23808 8944 23820
rect 8996 23808 9002 23860
rect 12250 23848 12256 23860
rect 9048 23820 12256 23848
rect 4062 23740 4068 23792
rect 4120 23780 4126 23792
rect 4341 23783 4399 23789
rect 4341 23780 4353 23783
rect 4120 23752 4353 23780
rect 4120 23740 4126 23752
rect 4341 23749 4353 23752
rect 4387 23749 4399 23783
rect 4341 23743 4399 23749
rect 5350 23740 5356 23792
rect 5408 23740 5414 23792
rect 2958 23672 2964 23724
rect 3016 23672 3022 23724
rect 4798 23672 4804 23724
rect 4856 23712 4862 23724
rect 5169 23715 5227 23721
rect 5169 23712 5181 23715
rect 4856 23684 5181 23712
rect 4856 23672 4862 23684
rect 5169 23681 5181 23684
rect 5215 23681 5227 23715
rect 5169 23675 5227 23681
rect 5445 23715 5503 23721
rect 5445 23681 5457 23715
rect 5491 23681 5503 23715
rect 5445 23675 5503 23681
rect 5537 23715 5595 23721
rect 5537 23681 5549 23715
rect 5583 23681 5595 23715
rect 5537 23675 5595 23681
rect 1394 23604 1400 23656
rect 1452 23644 1458 23656
rect 1581 23647 1639 23653
rect 1581 23644 1593 23647
rect 1452 23616 1593 23644
rect 1452 23604 1458 23616
rect 1581 23613 1593 23616
rect 1627 23613 1639 23647
rect 1581 23607 1639 23613
rect 1854 23604 1860 23656
rect 1912 23604 1918 23656
rect 2406 23604 2412 23656
rect 2464 23644 2470 23656
rect 3513 23647 3571 23653
rect 3513 23644 3525 23647
rect 2464 23616 3525 23644
rect 2464 23604 2470 23616
rect 3513 23613 3525 23616
rect 3559 23613 3571 23647
rect 3513 23607 3571 23613
rect 5077 23647 5135 23653
rect 5077 23613 5089 23647
rect 5123 23644 5135 23647
rect 5460 23644 5488 23675
rect 5123 23616 5488 23644
rect 5123 23613 5135 23616
rect 5077 23607 5135 23613
rect 3329 23579 3387 23585
rect 3329 23545 3341 23579
rect 3375 23576 3387 23579
rect 5092 23576 5120 23607
rect 5368 23588 5396 23616
rect 3375 23548 5120 23576
rect 3375 23545 3387 23548
rect 3329 23539 3387 23545
rect 5350 23536 5356 23588
rect 5408 23536 5414 23588
rect 2038 23468 2044 23520
rect 2096 23508 2102 23520
rect 2866 23508 2872 23520
rect 2096 23480 2872 23508
rect 2096 23468 2102 23480
rect 2866 23468 2872 23480
rect 2924 23468 2930 23520
rect 4433 23511 4491 23517
rect 4433 23477 4445 23511
rect 4479 23508 4491 23511
rect 4706 23508 4712 23520
rect 4479 23480 4712 23508
rect 4479 23477 4491 23480
rect 4433 23471 4491 23477
rect 4706 23468 4712 23480
rect 4764 23468 4770 23520
rect 5258 23468 5264 23520
rect 5316 23508 5322 23520
rect 5552 23508 5580 23675
rect 5810 23672 5816 23724
rect 5868 23712 5874 23724
rect 5997 23715 6055 23721
rect 5997 23712 6009 23715
rect 5868 23684 6009 23712
rect 5868 23672 5874 23684
rect 5997 23681 6009 23684
rect 6043 23681 6055 23715
rect 6104 23718 6132 23808
rect 9048 23789 9076 23820
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 12802 23808 12808 23860
rect 12860 23848 12866 23860
rect 12989 23851 13047 23857
rect 12989 23848 13001 23851
rect 12860 23820 13001 23848
rect 12860 23808 12866 23820
rect 12989 23817 13001 23820
rect 13035 23817 13047 23851
rect 12989 23811 13047 23817
rect 14826 23808 14832 23860
rect 14884 23848 14890 23860
rect 15010 23848 15016 23860
rect 14884 23820 15016 23848
rect 14884 23808 14890 23820
rect 15010 23808 15016 23820
rect 15068 23808 15074 23860
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 16390 23848 16396 23860
rect 15712 23820 16396 23848
rect 15712 23808 15718 23820
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 17678 23808 17684 23860
rect 17736 23848 17742 23860
rect 17736 23820 18092 23848
rect 17736 23808 17742 23820
rect 6733 23783 6791 23789
rect 6733 23749 6745 23783
rect 6779 23780 6791 23783
rect 9033 23783 9091 23789
rect 6779 23752 8984 23780
rect 6779 23749 6791 23752
rect 6733 23743 6791 23749
rect 6181 23718 6239 23721
rect 6104 23715 6239 23718
rect 6104 23690 6193 23715
rect 5997 23675 6055 23681
rect 6181 23681 6193 23690
rect 6227 23681 6239 23715
rect 6181 23675 6239 23681
rect 6365 23715 6423 23721
rect 6365 23681 6377 23715
rect 6411 23681 6423 23715
rect 6365 23675 6423 23681
rect 5626 23604 5632 23656
rect 5684 23604 5690 23656
rect 5718 23604 5724 23656
rect 5776 23644 5782 23656
rect 6380 23644 6408 23675
rect 6454 23672 6460 23724
rect 6512 23712 6518 23724
rect 6914 23721 6920 23724
rect 6641 23715 6699 23721
rect 6512 23684 6557 23712
rect 6512 23672 6518 23684
rect 6641 23681 6653 23715
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 6871 23715 6920 23721
rect 6871 23681 6883 23715
rect 6917 23681 6920 23715
rect 6871 23675 6920 23681
rect 5776 23616 6408 23644
rect 6656 23644 6684 23675
rect 6914 23672 6920 23675
rect 6972 23672 6978 23724
rect 7374 23712 7380 23724
rect 7024 23684 7380 23712
rect 7024 23644 7052 23684
rect 7374 23672 7380 23684
rect 7432 23672 7438 23724
rect 7926 23672 7932 23724
rect 7984 23672 7990 23724
rect 8294 23672 8300 23724
rect 8352 23672 8358 23724
rect 8757 23715 8815 23721
rect 8757 23681 8769 23715
rect 8803 23681 8815 23715
rect 8956 23712 8984 23752
rect 9033 23749 9045 23783
rect 9079 23749 9091 23783
rect 9033 23743 9091 23749
rect 9122 23740 9128 23792
rect 9180 23780 9186 23792
rect 9306 23780 9312 23792
rect 9180 23752 9312 23780
rect 9180 23740 9186 23752
rect 9306 23740 9312 23752
rect 9364 23780 9370 23792
rect 11685 23783 11743 23789
rect 9364 23752 11652 23780
rect 9364 23740 9370 23752
rect 10502 23712 10508 23724
rect 8956 23684 10508 23712
rect 8757 23675 8815 23681
rect 6656 23616 7052 23644
rect 5776 23604 5782 23616
rect 7190 23604 7196 23656
rect 7248 23644 7254 23656
rect 8772 23644 8800 23675
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 11054 23644 11060 23656
rect 7248 23616 11060 23644
rect 7248 23604 7254 23616
rect 11054 23604 11060 23616
rect 11112 23604 11118 23656
rect 11624 23644 11652 23752
rect 11685 23749 11697 23783
rect 11731 23749 11743 23783
rect 11685 23743 11743 23749
rect 11700 23712 11728 23743
rect 11882 23740 11888 23792
rect 11940 23740 11946 23792
rect 11974 23740 11980 23792
rect 12032 23780 12038 23792
rect 15930 23780 15936 23792
rect 12032 23752 13211 23780
rect 12032 23740 12038 23752
rect 13183 23724 13211 23752
rect 15764 23752 15936 23780
rect 12802 23712 12808 23724
rect 11700 23684 12808 23712
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 13170 23721 13176 23724
rect 13168 23712 13176 23721
rect 13131 23684 13176 23712
rect 13168 23675 13176 23684
rect 13170 23672 13176 23675
rect 13228 23672 13234 23724
rect 13262 23672 13268 23724
rect 13320 23672 13326 23724
rect 13354 23672 13360 23724
rect 13412 23672 13418 23724
rect 13538 23712 13544 23724
rect 13499 23684 13544 23712
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 13630 23672 13636 23724
rect 13688 23672 13694 23724
rect 15470 23672 15476 23724
rect 15528 23672 15534 23724
rect 15764 23721 15792 23752
rect 15930 23740 15936 23752
rect 15988 23780 15994 23792
rect 17696 23780 17724 23808
rect 15988 23752 17724 23780
rect 15988 23740 15994 23752
rect 17862 23740 17868 23792
rect 17920 23740 17926 23792
rect 18064 23789 18092 23820
rect 18138 23808 18144 23860
rect 18196 23848 18202 23860
rect 20165 23851 20223 23857
rect 20165 23848 20177 23851
rect 18196 23820 20177 23848
rect 18196 23808 18202 23820
rect 20165 23817 20177 23820
rect 20211 23848 20223 23851
rect 20211 23820 20300 23848
rect 20211 23817 20223 23820
rect 20165 23811 20223 23817
rect 18049 23783 18107 23789
rect 18049 23749 18061 23783
rect 18095 23749 18107 23783
rect 19242 23780 19248 23792
rect 18049 23743 18107 23749
rect 18616 23752 19248 23780
rect 15749 23715 15807 23721
rect 15749 23681 15761 23715
rect 15795 23681 15807 23715
rect 15749 23675 15807 23681
rect 15838 23672 15844 23724
rect 15896 23712 15902 23724
rect 18616 23721 18644 23752
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 19610 23740 19616 23792
rect 19668 23780 19674 23792
rect 19797 23783 19855 23789
rect 19797 23780 19809 23783
rect 19668 23752 19809 23780
rect 19668 23740 19674 23752
rect 19797 23749 19809 23752
rect 19843 23749 19855 23783
rect 19797 23743 19855 23749
rect 19886 23740 19892 23792
rect 19944 23780 19950 23792
rect 20272 23789 20300 23820
rect 20622 23808 20628 23860
rect 20680 23848 20686 23860
rect 20809 23851 20867 23857
rect 20809 23848 20821 23851
rect 20680 23820 20821 23848
rect 20680 23808 20686 23820
rect 20809 23817 20821 23820
rect 20855 23817 20867 23851
rect 24854 23848 24860 23860
rect 20809 23811 20867 23817
rect 22204 23820 24860 23848
rect 19997 23783 20055 23789
rect 19997 23780 20009 23783
rect 19944 23752 20009 23780
rect 19944 23740 19950 23752
rect 19997 23749 20009 23752
rect 20043 23749 20055 23783
rect 19997 23743 20055 23749
rect 20257 23783 20315 23789
rect 20257 23749 20269 23783
rect 20303 23749 20315 23783
rect 22204 23780 22232 23820
rect 24854 23808 24860 23820
rect 24912 23848 24918 23860
rect 26237 23851 26295 23857
rect 24912 23820 26004 23848
rect 24912 23808 24918 23820
rect 20257 23743 20315 23749
rect 20640 23752 22232 23780
rect 22281 23783 22339 23789
rect 20640 23724 20668 23752
rect 22281 23749 22293 23783
rect 22327 23780 22339 23783
rect 23934 23780 23940 23792
rect 22327 23752 23940 23780
rect 22327 23749 22339 23752
rect 22281 23743 22339 23749
rect 23934 23740 23940 23752
rect 23992 23740 23998 23792
rect 25130 23740 25136 23792
rect 25188 23780 25194 23792
rect 25976 23789 26004 23820
rect 26237 23817 26249 23851
rect 26283 23848 26295 23851
rect 27246 23848 27252 23860
rect 26283 23820 27252 23848
rect 26283 23817 26295 23820
rect 26237 23811 26295 23817
rect 27246 23808 27252 23820
rect 27304 23848 27310 23860
rect 29089 23851 29147 23857
rect 27304 23820 28856 23848
rect 27304 23808 27310 23820
rect 25961 23783 26019 23789
rect 25188 23752 25360 23780
rect 25188 23740 25194 23752
rect 18601 23715 18659 23721
rect 15896 23684 18460 23712
rect 15896 23672 15902 23684
rect 12342 23644 12348 23656
rect 11624 23616 12348 23644
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 5644 23576 5672 23604
rect 5644 23548 6408 23576
rect 5316 23480 5580 23508
rect 5316 23468 5322 23480
rect 5626 23468 5632 23520
rect 5684 23508 5690 23520
rect 5721 23511 5779 23517
rect 5721 23508 5733 23511
rect 5684 23480 5733 23508
rect 5684 23468 5690 23480
rect 5721 23477 5733 23480
rect 5767 23477 5779 23511
rect 5721 23471 5779 23477
rect 5902 23468 5908 23520
rect 5960 23508 5966 23520
rect 6270 23508 6276 23520
rect 5960 23480 6276 23508
rect 5960 23468 5966 23480
rect 6270 23468 6276 23480
rect 6328 23468 6334 23520
rect 6380 23508 6408 23548
rect 6454 23536 6460 23588
rect 6512 23576 6518 23588
rect 6638 23576 6644 23588
rect 6512 23548 6644 23576
rect 6512 23536 6518 23548
rect 6638 23536 6644 23548
rect 6696 23536 6702 23588
rect 7374 23536 7380 23588
rect 7432 23576 7438 23588
rect 14734 23576 14740 23588
rect 7432 23548 14740 23576
rect 7432 23536 7438 23548
rect 14734 23536 14740 23548
rect 14792 23536 14798 23588
rect 17034 23536 17040 23588
rect 17092 23576 17098 23588
rect 17770 23576 17776 23588
rect 17092 23548 17776 23576
rect 17092 23536 17098 23548
rect 17770 23536 17776 23548
rect 17828 23576 17834 23588
rect 18432 23576 18460 23684
rect 18601 23681 18613 23715
rect 18647 23681 18659 23715
rect 18601 23675 18659 23681
rect 18690 23672 18696 23724
rect 18748 23712 18754 23724
rect 18877 23715 18935 23721
rect 18877 23712 18889 23715
rect 18748 23684 18889 23712
rect 18748 23672 18754 23684
rect 18877 23681 18889 23684
rect 18923 23681 18935 23715
rect 18877 23675 18935 23681
rect 19153 23715 19211 23721
rect 19153 23681 19165 23715
rect 19199 23712 19211 23715
rect 19334 23712 19340 23724
rect 19199 23684 19340 23712
rect 19199 23681 19211 23684
rect 19153 23675 19211 23681
rect 19334 23672 19340 23684
rect 19392 23672 19398 23724
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23681 20499 23715
rect 20441 23675 20499 23681
rect 20533 23715 20591 23721
rect 20533 23681 20545 23715
rect 20579 23712 20591 23715
rect 20622 23712 20628 23724
rect 20579 23684 20628 23712
rect 20579 23681 20591 23684
rect 20533 23675 20591 23681
rect 18509 23647 18567 23653
rect 18509 23613 18521 23647
rect 18555 23644 18567 23647
rect 18555 23616 18741 23644
rect 18555 23613 18567 23616
rect 18509 23607 18567 23613
rect 18713 23576 18741 23616
rect 18966 23604 18972 23656
rect 19024 23604 19030 23656
rect 19242 23604 19248 23656
rect 19300 23644 19306 23656
rect 20456 23644 20484 23675
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 22094 23712 22100 23724
rect 20772 23684 22100 23712
rect 20772 23672 20778 23684
rect 22094 23672 22100 23684
rect 22152 23672 22158 23724
rect 22370 23672 22376 23724
rect 22428 23712 22434 23724
rect 25332 23721 25360 23752
rect 25961 23749 25973 23783
rect 26007 23749 26019 23783
rect 25961 23743 26019 23749
rect 28350 23740 28356 23792
rect 28408 23780 28414 23792
rect 28721 23783 28779 23789
rect 28721 23780 28733 23783
rect 28408 23752 28733 23780
rect 28408 23740 28414 23752
rect 28721 23749 28733 23752
rect 28767 23749 28779 23783
rect 28828 23780 28856 23820
rect 29089 23817 29101 23851
rect 29135 23848 29147 23851
rect 31846 23848 31852 23860
rect 29135 23820 31852 23848
rect 29135 23817 29147 23820
rect 29089 23811 29147 23817
rect 31846 23808 31852 23820
rect 31904 23808 31910 23860
rect 32122 23808 32128 23860
rect 32180 23848 32186 23860
rect 32398 23848 32404 23860
rect 32180 23820 32404 23848
rect 32180 23808 32186 23820
rect 32398 23808 32404 23820
rect 32456 23808 32462 23860
rect 28828 23752 29316 23780
rect 28721 23743 28779 23749
rect 22465 23715 22523 23721
rect 22465 23712 22477 23715
rect 22428 23684 22477 23712
rect 22428 23672 22434 23684
rect 22465 23681 22477 23684
rect 22511 23681 22523 23715
rect 22465 23675 22523 23681
rect 25317 23715 25375 23721
rect 25317 23681 25329 23715
rect 25363 23681 25375 23715
rect 25317 23675 25375 23681
rect 19300 23616 20484 23644
rect 19300 23604 19306 23616
rect 20990 23604 20996 23656
rect 21048 23604 21054 23656
rect 21082 23604 21088 23656
rect 21140 23644 21146 23656
rect 21358 23644 21364 23656
rect 21140 23616 21364 23644
rect 21140 23604 21146 23616
rect 21358 23604 21364 23616
rect 21416 23604 21422 23656
rect 21453 23647 21511 23653
rect 21453 23613 21465 23647
rect 21499 23613 21511 23647
rect 21453 23607 21511 23613
rect 17828 23548 18368 23576
rect 18432 23548 18552 23576
rect 18713 23548 18816 23576
rect 17828 23536 17834 23548
rect 7190 23508 7196 23520
rect 6380 23480 7196 23508
rect 7190 23468 7196 23480
rect 7248 23468 7254 23520
rect 7558 23468 7564 23520
rect 7616 23508 7622 23520
rect 8110 23508 8116 23520
rect 7616 23480 8116 23508
rect 7616 23468 7622 23480
rect 8110 23468 8116 23480
rect 8168 23508 8174 23520
rect 9033 23511 9091 23517
rect 9033 23508 9045 23511
rect 8168 23480 9045 23508
rect 8168 23468 8174 23480
rect 9033 23477 9045 23480
rect 9079 23477 9091 23511
rect 9033 23471 9091 23477
rect 11330 23468 11336 23520
rect 11388 23508 11394 23520
rect 11517 23511 11575 23517
rect 11517 23508 11529 23511
rect 11388 23480 11529 23508
rect 11388 23468 11394 23480
rect 11517 23477 11529 23480
rect 11563 23477 11575 23511
rect 11517 23471 11575 23477
rect 11698 23468 11704 23520
rect 11756 23508 11762 23520
rect 12250 23508 12256 23520
rect 11756 23480 12256 23508
rect 11756 23468 11762 23480
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 13078 23468 13084 23520
rect 13136 23508 13142 23520
rect 13538 23508 13544 23520
rect 13136 23480 13544 23508
rect 13136 23468 13142 23480
rect 13538 23468 13544 23480
rect 13596 23468 13602 23520
rect 17402 23468 17408 23520
rect 17460 23508 17466 23520
rect 17681 23511 17739 23517
rect 17681 23508 17693 23511
rect 17460 23480 17693 23508
rect 17460 23468 17466 23480
rect 17681 23477 17693 23480
rect 17727 23477 17739 23511
rect 17681 23471 17739 23477
rect 17862 23468 17868 23520
rect 17920 23468 17926 23520
rect 18138 23468 18144 23520
rect 18196 23508 18202 23520
rect 18233 23511 18291 23517
rect 18233 23508 18245 23511
rect 18196 23480 18245 23508
rect 18196 23468 18202 23480
rect 18233 23477 18245 23480
rect 18279 23477 18291 23511
rect 18340 23508 18368 23548
rect 18417 23511 18475 23517
rect 18417 23508 18429 23511
rect 18340 23480 18429 23508
rect 18233 23471 18291 23477
rect 18417 23477 18429 23480
rect 18463 23477 18475 23511
rect 18524 23508 18552 23548
rect 18693 23511 18751 23517
rect 18693 23508 18705 23511
rect 18524 23480 18705 23508
rect 18417 23471 18475 23477
rect 18693 23477 18705 23480
rect 18739 23477 18751 23511
rect 18788 23508 18816 23548
rect 19150 23536 19156 23588
rect 19208 23576 19214 23588
rect 20257 23579 20315 23585
rect 19208 23548 19334 23576
rect 19208 23536 19214 23548
rect 18966 23508 18972 23520
rect 18788 23480 18972 23508
rect 18693 23471 18751 23477
rect 18966 23468 18972 23480
rect 19024 23468 19030 23520
rect 19306 23508 19334 23548
rect 20257 23545 20269 23579
rect 20303 23576 20315 23579
rect 21468 23576 21496 23607
rect 25038 23604 25044 23656
rect 25096 23644 25102 23656
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 25096 23616 25145 23644
rect 25096 23604 25102 23616
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25332 23644 25360 23675
rect 25590 23672 25596 23724
rect 25648 23712 25654 23724
rect 25685 23715 25743 23721
rect 25685 23712 25697 23715
rect 25648 23684 25697 23712
rect 25648 23672 25654 23684
rect 25685 23681 25697 23684
rect 25731 23681 25743 23715
rect 25685 23675 25743 23681
rect 25869 23715 25927 23721
rect 25869 23681 25881 23715
rect 25915 23681 25927 23715
rect 25869 23675 25927 23681
rect 26053 23715 26111 23721
rect 26053 23681 26065 23715
rect 26099 23712 26111 23715
rect 26510 23712 26516 23724
rect 26099 23684 26516 23712
rect 26099 23681 26111 23684
rect 26053 23675 26111 23681
rect 25774 23644 25780 23656
rect 25332 23616 25780 23644
rect 25133 23607 25191 23613
rect 22094 23576 22100 23588
rect 20303 23548 22100 23576
rect 20303 23545 20315 23548
rect 20257 23539 20315 23545
rect 22094 23536 22100 23548
rect 22152 23536 22158 23588
rect 19981 23511 20039 23517
rect 19981 23508 19993 23511
rect 19306 23480 19993 23508
rect 19981 23477 19993 23480
rect 20027 23508 20039 23511
rect 20714 23508 20720 23520
rect 20027 23480 20720 23508
rect 20027 23477 20039 23480
rect 19981 23471 20039 23477
rect 20714 23468 20720 23480
rect 20772 23468 20778 23520
rect 21634 23468 21640 23520
rect 21692 23508 21698 23520
rect 22649 23511 22707 23517
rect 22649 23508 22661 23511
rect 21692 23480 22661 23508
rect 21692 23468 21698 23480
rect 22649 23477 22661 23480
rect 22695 23477 22707 23511
rect 25148 23508 25176 23607
rect 25774 23604 25780 23616
rect 25832 23604 25838 23656
rect 25884 23644 25912 23675
rect 26510 23672 26516 23684
rect 26568 23672 26574 23724
rect 28534 23672 28540 23724
rect 28592 23672 28598 23724
rect 28810 23672 28816 23724
rect 28868 23672 28874 23724
rect 28905 23715 28963 23721
rect 28905 23681 28917 23715
rect 28951 23681 28963 23715
rect 28905 23675 28963 23681
rect 25884 23616 26924 23644
rect 26896 23588 26924 23616
rect 28258 23604 28264 23656
rect 28316 23644 28322 23656
rect 28920 23644 28948 23675
rect 29178 23672 29184 23724
rect 29236 23672 29242 23724
rect 29288 23721 29316 23752
rect 30558 23740 30564 23792
rect 30616 23780 30622 23792
rect 30837 23783 30895 23789
rect 30837 23780 30849 23783
rect 30616 23752 30849 23780
rect 30616 23740 30622 23752
rect 30837 23749 30849 23752
rect 30883 23749 30895 23783
rect 30837 23743 30895 23749
rect 32600 23752 33364 23780
rect 29273 23715 29331 23721
rect 29273 23681 29285 23715
rect 29319 23681 29331 23715
rect 30699 23715 30757 23721
rect 30699 23712 30711 23715
rect 29273 23675 29331 23681
rect 29380 23684 30711 23712
rect 28316 23616 28948 23644
rect 28316 23604 28322 23616
rect 25501 23579 25559 23585
rect 25501 23545 25513 23579
rect 25547 23576 25559 23579
rect 26602 23576 26608 23588
rect 25547 23548 26608 23576
rect 25547 23545 25559 23548
rect 25501 23539 25559 23545
rect 26602 23536 26608 23548
rect 26660 23536 26666 23588
rect 26878 23536 26884 23588
rect 26936 23576 26942 23588
rect 29380 23576 29408 23684
rect 30699 23681 30711 23684
rect 30745 23681 30757 23715
rect 30699 23675 30757 23681
rect 30929 23715 30987 23721
rect 30929 23681 30941 23715
rect 30975 23681 30987 23715
rect 30929 23675 30987 23681
rect 29638 23604 29644 23656
rect 29696 23644 29702 23656
rect 30561 23647 30619 23653
rect 30561 23644 30573 23647
rect 29696 23616 30573 23644
rect 29696 23604 29702 23616
rect 30561 23613 30573 23616
rect 30607 23613 30619 23647
rect 30944 23644 30972 23675
rect 31018 23672 31024 23724
rect 31076 23672 31082 23724
rect 31110 23672 31116 23724
rect 31168 23712 31174 23724
rect 31168 23684 31432 23712
rect 31168 23672 31174 23684
rect 31294 23644 31300 23656
rect 30944 23616 31300 23644
rect 30561 23607 30619 23613
rect 31294 23604 31300 23616
rect 31352 23604 31358 23656
rect 31404 23644 31432 23684
rect 31478 23672 31484 23724
rect 31536 23712 31542 23724
rect 32600 23712 32628 23752
rect 33336 23721 33364 23752
rect 34146 23740 34152 23792
rect 34204 23780 34210 23792
rect 34204 23752 34744 23780
rect 34204 23740 34210 23752
rect 33321 23715 33379 23721
rect 31536 23684 32628 23712
rect 32784 23684 33180 23712
rect 31536 23672 31542 23684
rect 32784 23644 32812 23684
rect 31404 23616 32812 23644
rect 32858 23604 32864 23656
rect 32916 23644 32922 23656
rect 33042 23644 33048 23656
rect 32916 23616 33048 23644
rect 32916 23604 32922 23616
rect 33042 23604 33048 23616
rect 33100 23604 33106 23656
rect 33152 23644 33180 23684
rect 33321 23681 33333 23715
rect 33367 23681 33379 23715
rect 33321 23675 33379 23681
rect 34422 23672 34428 23724
rect 34480 23672 34486 23724
rect 34606 23672 34612 23724
rect 34664 23672 34670 23724
rect 34716 23721 34744 23752
rect 34701 23715 34759 23721
rect 34701 23681 34713 23715
rect 34747 23681 34759 23715
rect 34701 23675 34759 23681
rect 34790 23644 34796 23656
rect 33152 23616 34796 23644
rect 34790 23604 34796 23616
rect 34848 23604 34854 23656
rect 26936 23548 29408 23576
rect 29549 23579 29607 23585
rect 26936 23536 26942 23548
rect 29549 23545 29561 23579
rect 29595 23576 29607 23579
rect 33505 23579 33563 23585
rect 29595 23548 33456 23576
rect 29595 23545 29607 23548
rect 29549 23539 29607 23545
rect 26050 23508 26056 23520
rect 25148 23480 26056 23508
rect 22649 23471 22707 23477
rect 26050 23468 26056 23480
rect 26108 23468 26114 23520
rect 26234 23468 26240 23520
rect 26292 23508 26298 23520
rect 28902 23508 28908 23520
rect 26292 23480 28908 23508
rect 26292 23468 26298 23480
rect 28902 23468 28908 23480
rect 28960 23468 28966 23520
rect 29270 23468 29276 23520
rect 29328 23508 29334 23520
rect 29365 23511 29423 23517
rect 29365 23508 29377 23511
rect 29328 23480 29377 23508
rect 29328 23468 29334 23480
rect 29365 23477 29377 23480
rect 29411 23508 29423 23511
rect 31110 23508 31116 23520
rect 29411 23480 31116 23508
rect 29411 23477 29423 23480
rect 29365 23471 29423 23477
rect 31110 23468 31116 23480
rect 31168 23468 31174 23520
rect 31205 23511 31263 23517
rect 31205 23477 31217 23511
rect 31251 23508 31263 23511
rect 31754 23508 31760 23520
rect 31251 23480 31760 23508
rect 31251 23477 31263 23480
rect 31205 23471 31263 23477
rect 31754 23468 31760 23480
rect 31812 23508 31818 23520
rect 32766 23508 32772 23520
rect 31812 23480 32772 23508
rect 31812 23468 31818 23480
rect 32766 23468 32772 23480
rect 32824 23468 32830 23520
rect 33134 23468 33140 23520
rect 33192 23468 33198 23520
rect 33428 23508 33456 23548
rect 33505 23545 33517 23579
rect 33551 23576 33563 23579
rect 34606 23576 34612 23588
rect 33551 23548 34612 23576
rect 33551 23545 33563 23548
rect 33505 23539 33563 23545
rect 34606 23536 34612 23548
rect 34664 23536 34670 23588
rect 34517 23511 34575 23517
rect 34517 23508 34529 23511
rect 33428 23480 34529 23508
rect 34517 23477 34529 23480
rect 34563 23508 34575 23511
rect 34790 23508 34796 23520
rect 34563 23480 34796 23508
rect 34563 23477 34575 23480
rect 34517 23471 34575 23477
rect 34790 23468 34796 23480
rect 34848 23468 34854 23520
rect 34885 23511 34943 23517
rect 34885 23477 34897 23511
rect 34931 23508 34943 23511
rect 35434 23508 35440 23520
rect 34931 23480 35440 23508
rect 34931 23477 34943 23480
rect 34885 23471 34943 23477
rect 35434 23468 35440 23480
rect 35492 23468 35498 23520
rect 1104 23418 36432 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 36432 23418
rect 1104 23344 36432 23366
rect 4246 23264 4252 23316
rect 4304 23304 4310 23316
rect 5902 23304 5908 23316
rect 4304 23276 5908 23304
rect 4304 23264 4310 23276
rect 5902 23264 5908 23276
rect 5960 23264 5966 23316
rect 5994 23264 6000 23316
rect 6052 23304 6058 23316
rect 6273 23307 6331 23313
rect 6273 23304 6285 23307
rect 6052 23276 6285 23304
rect 6052 23264 6058 23276
rect 6273 23273 6285 23276
rect 6319 23273 6331 23307
rect 6273 23267 6331 23273
rect 6362 23264 6368 23316
rect 6420 23304 6426 23316
rect 6733 23307 6791 23313
rect 6733 23304 6745 23307
rect 6420 23276 6745 23304
rect 6420 23264 6426 23276
rect 6733 23273 6745 23276
rect 6779 23304 6791 23307
rect 7190 23304 7196 23316
rect 6779 23276 7196 23304
rect 6779 23273 6791 23276
rect 6733 23267 6791 23273
rect 7190 23264 7196 23276
rect 7248 23264 7254 23316
rect 9122 23264 9128 23316
rect 9180 23304 9186 23316
rect 11974 23304 11980 23316
rect 9180 23276 11980 23304
rect 9180 23264 9186 23276
rect 11974 23264 11980 23276
rect 12032 23264 12038 23316
rect 13081 23307 13139 23313
rect 13081 23304 13093 23307
rect 12192 23276 13093 23304
rect 3878 23196 3884 23248
rect 3936 23236 3942 23248
rect 3936 23208 5792 23236
rect 3936 23196 3942 23208
rect 2406 23168 2412 23180
rect 1412 23140 2412 23168
rect 1412 23112 1440 23140
rect 2406 23128 2412 23140
rect 2464 23168 2470 23180
rect 2464 23140 3280 23168
rect 2464 23128 2470 23140
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 3252 23109 3280 23140
rect 3326 23128 3332 23180
rect 3384 23168 3390 23180
rect 4246 23168 4252 23180
rect 3384 23140 4252 23168
rect 3384 23128 3390 23140
rect 4246 23128 4252 23140
rect 4304 23168 4310 23180
rect 4341 23171 4399 23177
rect 4341 23168 4353 23171
rect 4304 23140 4353 23168
rect 4304 23128 4310 23140
rect 4341 23137 4353 23140
rect 4387 23137 4399 23171
rect 4341 23131 4399 23137
rect 4448 23140 5028 23168
rect 3237 23103 3295 23109
rect 3237 23069 3249 23103
rect 3283 23069 3295 23103
rect 3237 23063 3295 23069
rect 3970 23060 3976 23112
rect 4028 23100 4034 23112
rect 4448 23100 4476 23140
rect 4028 23072 4476 23100
rect 4028 23060 4034 23072
rect 4522 23060 4528 23112
rect 4580 23100 4586 23112
rect 5000 23109 5028 23140
rect 4893 23103 4951 23109
rect 4893 23100 4905 23103
rect 4580 23072 4905 23100
rect 4580 23060 4586 23072
rect 4893 23069 4905 23072
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 4986 23103 5044 23109
rect 4986 23069 4998 23103
rect 5032 23069 5044 23103
rect 4986 23063 5044 23069
rect 5166 23060 5172 23112
rect 5224 23060 5230 23112
rect 5399 23103 5457 23109
rect 5399 23069 5411 23103
rect 5445 23069 5457 23103
rect 5626 23102 5632 23114
rect 5589 23074 5632 23102
rect 5399 23063 5457 23069
rect 1670 22992 1676 23044
rect 1728 22992 1734 23044
rect 2958 23032 2964 23044
rect 2898 23004 2964 23032
rect 2958 22992 2964 23004
rect 3016 22992 3022 23044
rect 4157 23035 4215 23041
rect 4157 23001 4169 23035
rect 4203 23032 4215 23035
rect 4614 23032 4620 23044
rect 4203 23004 4620 23032
rect 4203 23001 4215 23004
rect 4157 22995 4215 23001
rect 4614 22992 4620 23004
rect 4672 22992 4678 23044
rect 4798 22992 4804 23044
rect 4856 23032 4862 23044
rect 5184 23032 5212 23060
rect 4856 23004 5212 23032
rect 5261 23035 5319 23041
rect 4856 22992 4862 23004
rect 5261 23001 5273 23035
rect 5307 23001 5319 23035
rect 5414 23032 5442 23063
rect 5626 23062 5632 23074
rect 5684 23062 5690 23114
rect 5764 23109 5792 23208
rect 6914 23196 6920 23248
rect 6972 23196 6978 23248
rect 10318 23196 10324 23248
rect 10376 23236 10382 23248
rect 10962 23236 10968 23248
rect 10376 23208 10968 23236
rect 10376 23196 10382 23208
rect 10962 23196 10968 23208
rect 11020 23196 11026 23248
rect 12192 23236 12220 23276
rect 13081 23273 13093 23276
rect 13127 23304 13139 23307
rect 13170 23304 13176 23316
rect 13127 23276 13176 23304
rect 13127 23273 13139 23276
rect 13081 23267 13139 23273
rect 13170 23264 13176 23276
rect 13228 23264 13234 23316
rect 17034 23264 17040 23316
rect 17092 23264 17098 23316
rect 17221 23307 17279 23313
rect 17221 23273 17233 23307
rect 17267 23304 17279 23307
rect 17267 23276 17540 23304
rect 17267 23273 17279 23276
rect 17221 23267 17279 23273
rect 11072 23208 12220 23236
rect 6638 23168 6644 23180
rect 5917 23140 6644 23168
rect 5917 23109 5945 23140
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 6932 23168 6960 23196
rect 8202 23168 8208 23180
rect 6840 23140 8208 23168
rect 5764 23103 5825 23109
rect 5764 23072 5779 23103
rect 5767 23069 5779 23072
rect 5813 23069 5825 23103
rect 5767 23063 5825 23069
rect 5905 23103 5963 23109
rect 5905 23069 5917 23103
rect 5951 23069 5963 23103
rect 5905 23063 5963 23069
rect 6094 23103 6152 23109
rect 6094 23069 6106 23103
rect 6140 23100 6152 23103
rect 6840 23100 6868 23140
rect 6140 23072 6868 23100
rect 6140 23069 6152 23072
rect 6094 23063 6152 23069
rect 5414 23004 5856 23032
rect 5261 22995 5319 23001
rect 3145 22967 3203 22973
rect 3145 22933 3157 22967
rect 3191 22964 3203 22967
rect 3694 22964 3700 22976
rect 3191 22936 3700 22964
rect 3191 22933 3203 22936
rect 3145 22927 3203 22933
rect 3694 22924 3700 22936
rect 3752 22924 3758 22976
rect 3789 22967 3847 22973
rect 3789 22933 3801 22967
rect 3835 22964 3847 22967
rect 4062 22964 4068 22976
rect 3835 22936 4068 22964
rect 3835 22933 3847 22936
rect 3789 22927 3847 22933
rect 4062 22924 4068 22936
rect 4120 22924 4126 22976
rect 4246 22924 4252 22976
rect 4304 22924 4310 22976
rect 5074 22924 5080 22976
rect 5132 22964 5138 22976
rect 5276 22964 5304 22995
rect 5132 22936 5304 22964
rect 5537 22967 5595 22973
rect 5132 22924 5138 22936
rect 5537 22933 5549 22967
rect 5583 22964 5595 22967
rect 5626 22964 5632 22976
rect 5583 22936 5632 22964
rect 5583 22933 5595 22936
rect 5537 22927 5595 22933
rect 5626 22924 5632 22936
rect 5684 22924 5690 22976
rect 5828 22964 5856 23004
rect 5994 22992 6000 23044
rect 6052 22992 6058 23044
rect 6104 22964 6132 23063
rect 6914 23060 6920 23112
rect 6972 23100 6978 23112
rect 7101 23103 7159 23109
rect 7101 23100 7113 23103
rect 6972 23072 7113 23100
rect 6972 23060 6978 23072
rect 7101 23069 7113 23072
rect 7147 23069 7159 23103
rect 7101 23063 7159 23069
rect 7190 23060 7196 23112
rect 7248 23060 7254 23112
rect 7576 23109 7604 23140
rect 8202 23128 8208 23140
rect 8260 23168 8266 23180
rect 8260 23140 8892 23168
rect 8260 23128 8266 23140
rect 7566 23103 7624 23109
rect 7566 23069 7578 23103
rect 7612 23069 7624 23103
rect 7566 23063 7624 23069
rect 8386 23060 8392 23112
rect 8444 23060 8450 23112
rect 8573 23103 8631 23109
rect 8573 23069 8585 23103
rect 8619 23069 8631 23103
rect 8573 23063 8631 23069
rect 6638 22992 6644 23044
rect 6696 23032 6702 23044
rect 6825 23035 6883 23041
rect 6825 23032 6837 23035
rect 6696 23004 6837 23032
rect 6696 22992 6702 23004
rect 6825 23001 6837 23004
rect 6871 23001 6883 23035
rect 6825 22995 6883 23001
rect 7009 23035 7067 23041
rect 7009 23001 7021 23035
rect 7055 23001 7067 23035
rect 7009 22995 7067 23001
rect 5828 22936 6132 22964
rect 7024 22964 7052 22995
rect 7374 22992 7380 23044
rect 7432 22992 7438 23044
rect 7469 23035 7527 23041
rect 7469 23001 7481 23035
rect 7515 23032 7527 23035
rect 7515 23004 8432 23032
rect 7515 23001 7527 23004
rect 7469 22995 7527 23001
rect 7745 22967 7803 22973
rect 7745 22964 7757 22967
rect 7024 22936 7757 22964
rect 7745 22933 7757 22936
rect 7791 22933 7803 22967
rect 7745 22927 7803 22933
rect 7834 22924 7840 22976
rect 7892 22964 7898 22976
rect 8205 22967 8263 22973
rect 8205 22964 8217 22967
rect 7892 22936 8217 22964
rect 7892 22924 7898 22936
rect 8205 22933 8217 22936
rect 8251 22933 8263 22967
rect 8404 22964 8432 23004
rect 8478 22992 8484 23044
rect 8536 22992 8542 23044
rect 8588 23032 8616 23063
rect 8754 23060 8760 23112
rect 8812 23060 8818 23112
rect 8864 23100 8892 23140
rect 9582 23128 9588 23180
rect 9640 23168 9646 23180
rect 11072 23168 11100 23208
rect 9640 23140 11100 23168
rect 9640 23128 9646 23140
rect 11146 23128 11152 23180
rect 11204 23128 11210 23180
rect 11054 23100 11060 23112
rect 8864 23072 11060 23100
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 11330 23100 11336 23112
rect 11388 23109 11394 23112
rect 11514 23109 11520 23112
rect 11298 23072 11336 23100
rect 11330 23060 11336 23072
rect 11388 23063 11398 23109
rect 11481 23103 11520 23109
rect 11481 23069 11493 23103
rect 11481 23063 11520 23069
rect 11388 23060 11394 23063
rect 11514 23060 11520 23063
rect 11572 23060 11578 23112
rect 11798 23103 11856 23109
rect 11798 23069 11810 23103
rect 11844 23100 11856 23103
rect 11900 23100 11928 23208
rect 12250 23196 12256 23248
rect 12308 23236 12314 23248
rect 13357 23239 13415 23245
rect 13357 23236 13369 23239
rect 12308 23208 13369 23236
rect 12308 23196 12314 23208
rect 13357 23205 13369 23208
rect 13403 23205 13415 23239
rect 13357 23199 13415 23205
rect 14274 23196 14280 23248
rect 14332 23236 14338 23248
rect 14369 23239 14427 23245
rect 14369 23236 14381 23239
rect 14332 23208 14381 23236
rect 14332 23196 14338 23208
rect 14369 23205 14381 23208
rect 14415 23236 14427 23239
rect 14550 23236 14556 23248
rect 14415 23208 14556 23236
rect 14415 23205 14427 23208
rect 14369 23199 14427 23205
rect 14550 23196 14556 23208
rect 14608 23196 14614 23248
rect 16482 23196 16488 23248
rect 16540 23236 16546 23248
rect 17405 23239 17463 23245
rect 17405 23236 17417 23239
rect 16540 23208 17417 23236
rect 16540 23196 16546 23208
rect 17405 23205 17417 23208
rect 17451 23205 17463 23239
rect 17512 23236 17540 23276
rect 17586 23264 17592 23316
rect 17644 23264 17650 23316
rect 17678 23264 17684 23316
rect 17736 23304 17742 23316
rect 17736 23276 18552 23304
rect 17736 23264 17742 23276
rect 18230 23236 18236 23248
rect 17512 23208 18236 23236
rect 17405 23199 17463 23205
rect 18230 23196 18236 23208
rect 18288 23196 18294 23248
rect 13446 23128 13452 23180
rect 13504 23168 13510 23180
rect 13725 23171 13783 23177
rect 13725 23168 13737 23171
rect 13504 23140 13737 23168
rect 13504 23128 13510 23140
rect 13725 23137 13737 23140
rect 13771 23168 13783 23171
rect 14734 23168 14740 23180
rect 13771 23140 14740 23168
rect 13771 23137 13783 23140
rect 13725 23131 13783 23137
rect 14734 23128 14740 23140
rect 14792 23128 14798 23180
rect 15838 23168 15844 23180
rect 14936 23140 15844 23168
rect 11844 23072 11928 23100
rect 11844 23069 11856 23072
rect 11798 23063 11856 23069
rect 11974 23060 11980 23112
rect 12032 23100 12038 23112
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 12032 23072 12081 23100
rect 12032 23060 12038 23072
rect 12069 23069 12081 23072
rect 12115 23069 12127 23103
rect 12069 23063 12127 23069
rect 12253 23103 12311 23109
rect 12253 23069 12265 23103
rect 12299 23100 12311 23103
rect 12342 23100 12348 23112
rect 12299 23072 12348 23100
rect 12299 23069 12311 23072
rect 12253 23063 12311 23069
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 12618 23060 12624 23112
rect 12676 23060 12682 23112
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23100 12771 23103
rect 13081 23103 13139 23109
rect 13081 23100 13093 23103
rect 12759 23072 13093 23100
rect 12759 23069 12771 23072
rect 12713 23063 12771 23069
rect 13081 23069 13093 23072
rect 13127 23069 13139 23103
rect 13081 23063 13139 23069
rect 13265 23103 13323 23109
rect 13265 23069 13277 23103
rect 13311 23069 13323 23103
rect 13265 23063 13323 23069
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23100 13599 23103
rect 13587 23072 14320 23100
rect 13587 23069 13599 23072
rect 13541 23063 13599 23069
rect 8588 23004 8800 23032
rect 8772 22976 8800 23004
rect 11606 22992 11612 23044
rect 11664 22992 11670 23044
rect 11701 23035 11759 23041
rect 11701 23001 11713 23035
rect 11747 23001 11759 23035
rect 11701 22995 11759 23001
rect 8570 22964 8576 22976
rect 8404 22936 8576 22964
rect 8205 22927 8263 22933
rect 8570 22924 8576 22936
rect 8628 22924 8634 22976
rect 8754 22924 8760 22976
rect 8812 22924 8818 22976
rect 9398 22924 9404 22976
rect 9456 22964 9462 22976
rect 9950 22964 9956 22976
rect 9456 22936 9956 22964
rect 9456 22924 9462 22936
rect 9950 22924 9956 22936
rect 10008 22924 10014 22976
rect 10318 22924 10324 22976
rect 10376 22964 10382 22976
rect 10597 22967 10655 22973
rect 10597 22964 10609 22967
rect 10376 22936 10609 22964
rect 10376 22924 10382 22936
rect 10597 22933 10609 22936
rect 10643 22933 10655 22967
rect 10597 22927 10655 22933
rect 11054 22924 11060 22976
rect 11112 22964 11118 22976
rect 11716 22964 11744 22995
rect 11882 22992 11888 23044
rect 11940 23032 11946 23044
rect 12437 23035 12495 23041
rect 12437 23032 12449 23035
rect 11940 23004 12449 23032
rect 11940 22992 11946 23004
rect 12084 22976 12112 23004
rect 12437 23001 12449 23004
rect 12483 23001 12495 23035
rect 12437 22995 12495 23001
rect 12526 22992 12532 23044
rect 12584 23032 12590 23044
rect 12728 23032 12756 23063
rect 12584 23004 12756 23032
rect 12584 22992 12590 23004
rect 12802 22992 12808 23044
rect 12860 23032 12866 23044
rect 13280 23032 13308 23063
rect 13814 23032 13820 23044
rect 12860 23004 13820 23032
rect 12860 22992 12866 23004
rect 13814 22992 13820 23004
rect 13872 22992 13878 23044
rect 14292 23032 14320 23072
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 14550 23100 14556 23112
rect 14424 23072 14556 23100
rect 14424 23060 14430 23072
rect 14550 23060 14556 23072
rect 14608 23100 14614 23112
rect 14645 23103 14703 23109
rect 14645 23100 14657 23103
rect 14608 23072 14657 23100
rect 14608 23060 14614 23072
rect 14645 23069 14657 23072
rect 14691 23069 14703 23103
rect 14645 23063 14703 23069
rect 14936 23032 14964 23140
rect 15838 23128 15844 23140
rect 15896 23128 15902 23180
rect 17954 23128 17960 23180
rect 18012 23168 18018 23180
rect 18524 23177 18552 23276
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 20530 23304 20536 23316
rect 19392 23276 20536 23304
rect 19392 23264 19398 23276
rect 20530 23264 20536 23276
rect 20588 23264 20594 23316
rect 20990 23264 20996 23316
rect 21048 23304 21054 23316
rect 21634 23304 21640 23316
rect 21048 23276 21640 23304
rect 21048 23264 21054 23276
rect 21634 23264 21640 23276
rect 21692 23264 21698 23316
rect 22281 23307 22339 23313
rect 22281 23273 22293 23307
rect 22327 23304 22339 23307
rect 23382 23304 23388 23316
rect 22327 23276 23388 23304
rect 22327 23273 22339 23276
rect 22281 23267 22339 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 25222 23264 25228 23316
rect 25280 23304 25286 23316
rect 25593 23307 25651 23313
rect 25593 23304 25605 23307
rect 25280 23276 25605 23304
rect 25280 23264 25286 23276
rect 25593 23273 25605 23276
rect 25639 23304 25651 23307
rect 27614 23304 27620 23316
rect 25639 23276 27620 23304
rect 25639 23273 25651 23276
rect 25593 23267 25651 23273
rect 27614 23264 27620 23276
rect 27672 23264 27678 23316
rect 28445 23307 28503 23313
rect 28445 23273 28457 23307
rect 28491 23304 28503 23307
rect 29178 23304 29184 23316
rect 28491 23276 29184 23304
rect 28491 23273 28503 23276
rect 28445 23267 28503 23273
rect 29178 23264 29184 23276
rect 29236 23264 29242 23316
rect 32582 23264 32588 23316
rect 32640 23304 32646 23316
rect 33962 23304 33968 23316
rect 32640 23276 33968 23304
rect 32640 23264 32646 23276
rect 33962 23264 33968 23276
rect 34020 23264 34026 23316
rect 25314 23236 25320 23248
rect 18616 23208 25320 23236
rect 18616 23177 18644 23208
rect 25314 23196 25320 23208
rect 25372 23196 25378 23248
rect 25866 23196 25872 23248
rect 25924 23236 25930 23248
rect 26510 23236 26516 23248
rect 25924 23208 26516 23236
rect 25924 23196 25930 23208
rect 26510 23196 26516 23208
rect 26568 23196 26574 23248
rect 18325 23171 18383 23177
rect 18325 23168 18337 23171
rect 18012 23140 18337 23168
rect 18012 23128 18018 23140
rect 18325 23137 18337 23140
rect 18371 23137 18383 23171
rect 18325 23131 18383 23137
rect 18509 23171 18567 23177
rect 18509 23137 18521 23171
rect 18555 23137 18567 23171
rect 18509 23131 18567 23137
rect 18601 23171 18659 23177
rect 18601 23137 18613 23171
rect 18647 23137 18659 23171
rect 18601 23131 18659 23137
rect 18874 23128 18880 23180
rect 18932 23168 18938 23180
rect 19242 23168 19248 23180
rect 18932 23140 19248 23168
rect 18932 23128 18938 23140
rect 19242 23128 19248 23140
rect 19300 23128 19306 23180
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 20622 23168 20628 23180
rect 19392 23140 20628 23168
rect 19392 23128 19398 23140
rect 20622 23128 20628 23140
rect 20680 23168 20686 23180
rect 21545 23171 21603 23177
rect 21545 23168 21557 23171
rect 20680 23140 21557 23168
rect 20680 23128 20686 23140
rect 21545 23137 21557 23140
rect 21591 23137 21603 23171
rect 21545 23131 21603 23137
rect 21634 23128 21640 23180
rect 21692 23168 21698 23180
rect 21692 23140 23060 23168
rect 21692 23128 21698 23140
rect 15010 23060 15016 23112
rect 15068 23060 15074 23112
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23100 15531 23103
rect 15654 23100 15660 23112
rect 15519 23072 15660 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 15749 23103 15807 23109
rect 15749 23069 15761 23103
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 14292 23004 14964 23032
rect 15194 22992 15200 23044
rect 15252 23032 15258 23044
rect 15764 23032 15792 23063
rect 15930 23060 15936 23112
rect 15988 23060 15994 23112
rect 16117 23103 16175 23109
rect 16117 23069 16129 23103
rect 16163 23100 16175 23103
rect 16298 23100 16304 23112
rect 16163 23072 16304 23100
rect 16163 23069 16175 23072
rect 16117 23063 16175 23069
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 16850 23060 16856 23112
rect 16908 23060 16914 23112
rect 16942 23060 16948 23112
rect 17000 23060 17006 23112
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23100 18475 23103
rect 18690 23100 18696 23112
rect 18463 23072 18696 23100
rect 18463 23069 18475 23072
rect 18417 23063 18475 23069
rect 18690 23060 18696 23072
rect 18748 23060 18754 23112
rect 19610 23060 19616 23112
rect 19668 23100 19674 23112
rect 21821 23103 21879 23109
rect 21821 23100 21833 23103
rect 19668 23072 21833 23100
rect 19668 23060 19674 23072
rect 21821 23069 21833 23072
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 17034 23032 17040 23044
rect 15252 23004 17040 23032
rect 15252 22992 15258 23004
rect 17034 22992 17040 23004
rect 17092 22992 17098 23044
rect 17770 22992 17776 23044
rect 17828 23032 17834 23044
rect 18598 23032 18604 23044
rect 17828 23004 18604 23032
rect 17828 22992 17834 23004
rect 18598 22992 18604 23004
rect 18656 22992 18662 23044
rect 11112 22936 11744 22964
rect 11112 22924 11118 22936
rect 11974 22924 11980 22976
rect 12032 22924 12038 22976
rect 12066 22924 12072 22976
rect 12124 22924 12130 22976
rect 12158 22924 12164 22976
rect 12216 22924 12222 22976
rect 12894 22924 12900 22976
rect 12952 22964 12958 22976
rect 13722 22964 13728 22976
rect 12952 22936 13728 22964
rect 12952 22924 12958 22936
rect 13722 22924 13728 22936
rect 13780 22924 13786 22976
rect 15746 22924 15752 22976
rect 15804 22964 15810 22976
rect 16025 22967 16083 22973
rect 16025 22964 16037 22967
rect 15804 22936 16037 22964
rect 15804 22924 15810 22936
rect 16025 22933 16037 22936
rect 16071 22933 16083 22967
rect 16025 22927 16083 22933
rect 17573 22967 17631 22973
rect 17573 22933 17585 22967
rect 17619 22964 17631 22967
rect 17678 22964 17684 22976
rect 17619 22936 17684 22964
rect 17619 22933 17631 22936
rect 17573 22927 17631 22933
rect 17678 22924 17684 22936
rect 17736 22924 17742 22976
rect 18138 22924 18144 22976
rect 18196 22924 18202 22976
rect 21836 22964 21864 23063
rect 21910 23060 21916 23112
rect 21968 23100 21974 23112
rect 21968 23072 22232 23100
rect 21968 23060 21974 23072
rect 22002 22992 22008 23044
rect 22060 22992 22066 23044
rect 22094 22992 22100 23044
rect 22152 22992 22158 23044
rect 22204 23032 22232 23072
rect 22554 23060 22560 23112
rect 22612 23060 22618 23112
rect 22830 23060 22836 23112
rect 22888 23060 22894 23112
rect 23032 23109 23060 23140
rect 23017 23103 23075 23109
rect 23017 23069 23029 23103
rect 23063 23069 23075 23103
rect 23017 23063 23075 23069
rect 23109 23103 23167 23109
rect 23109 23069 23121 23103
rect 23155 23100 23167 23103
rect 24210 23100 24216 23112
rect 23155 23072 24216 23100
rect 23155 23069 23167 23072
rect 23109 23063 23167 23069
rect 24210 23060 24216 23072
rect 24268 23060 24274 23112
rect 25774 23060 25780 23112
rect 25832 23060 25838 23112
rect 25866 23060 25872 23112
rect 25924 23060 25930 23112
rect 27614 23060 27620 23112
rect 27672 23100 27678 23112
rect 27893 23103 27951 23109
rect 27893 23100 27905 23103
rect 27672 23072 27905 23100
rect 27672 23060 27678 23072
rect 27893 23069 27905 23072
rect 27939 23069 27951 23103
rect 27893 23063 27951 23069
rect 28258 23060 28264 23112
rect 28316 23060 28322 23112
rect 22297 23035 22355 23041
rect 22297 23032 22309 23035
rect 22204 23004 22309 23032
rect 22297 23001 22309 23004
rect 22343 23001 22355 23035
rect 22572 23032 22600 23060
rect 24118 23032 24124 23044
rect 22297 22995 22355 23001
rect 22388 23004 24124 23032
rect 22388 22964 22416 23004
rect 24118 22992 24124 23004
rect 24176 22992 24182 23044
rect 25590 22992 25596 23044
rect 25648 23032 25654 23044
rect 27062 23032 27068 23044
rect 25648 23004 27068 23032
rect 25648 22992 25654 23004
rect 27062 22992 27068 23004
rect 27120 23032 27126 23044
rect 28077 23035 28135 23041
rect 28077 23032 28089 23035
rect 27120 23004 28089 23032
rect 27120 22992 27126 23004
rect 28077 23001 28089 23004
rect 28123 23001 28135 23035
rect 28077 22995 28135 23001
rect 28166 22992 28172 23044
rect 28224 22992 28230 23044
rect 21836 22936 22416 22964
rect 22465 22967 22523 22973
rect 22465 22933 22477 22967
rect 22511 22964 22523 22967
rect 22554 22964 22560 22976
rect 22511 22936 22560 22964
rect 22511 22933 22523 22936
rect 22465 22927 22523 22933
rect 22554 22924 22560 22936
rect 22612 22924 22618 22976
rect 22646 22924 22652 22976
rect 22704 22924 22710 22976
rect 30558 22924 30564 22976
rect 30616 22964 30622 22976
rect 31018 22964 31024 22976
rect 30616 22936 31024 22964
rect 30616 22924 30622 22936
rect 31018 22924 31024 22936
rect 31076 22924 31082 22976
rect 1104 22874 36432 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 36432 22874
rect 1104 22800 36432 22822
rect 1765 22763 1823 22769
rect 1765 22729 1777 22763
rect 1811 22760 1823 22763
rect 1854 22760 1860 22772
rect 1811 22732 1860 22760
rect 1811 22729 1823 22732
rect 1765 22723 1823 22729
rect 1854 22720 1860 22732
rect 1912 22720 1918 22772
rect 2133 22763 2191 22769
rect 2133 22729 2145 22763
rect 2179 22760 2191 22763
rect 4706 22760 4712 22772
rect 2179 22732 4712 22760
rect 2179 22729 2191 22732
rect 2133 22723 2191 22729
rect 4706 22720 4712 22732
rect 4764 22720 4770 22772
rect 4890 22720 4896 22772
rect 4948 22760 4954 22772
rect 5169 22763 5227 22769
rect 5169 22760 5181 22763
rect 4948 22732 5181 22760
rect 4948 22720 4954 22732
rect 5169 22729 5181 22732
rect 5215 22729 5227 22763
rect 6822 22760 6828 22772
rect 5169 22723 5227 22729
rect 5764 22732 6828 22760
rect 4062 22652 4068 22704
rect 4120 22652 4126 22704
rect 4154 22652 4160 22704
rect 4212 22692 4218 22704
rect 5445 22695 5503 22701
rect 5445 22692 5457 22695
rect 4212 22664 5457 22692
rect 4212 22652 4218 22664
rect 5445 22661 5457 22664
rect 5491 22661 5503 22695
rect 5764 22692 5792 22732
rect 6822 22720 6828 22732
rect 6880 22720 6886 22772
rect 6914 22720 6920 22772
rect 6972 22720 6978 22772
rect 8202 22720 8208 22772
rect 8260 22760 8266 22772
rect 8481 22763 8539 22769
rect 8260 22732 8340 22760
rect 8260 22720 8266 22732
rect 6546 22692 6552 22704
rect 5445 22655 5503 22661
rect 5736 22664 5792 22692
rect 5920 22664 6552 22692
rect 2225 22627 2283 22633
rect 2225 22593 2237 22627
rect 2271 22624 2283 22627
rect 2498 22624 2504 22636
rect 2271 22596 2504 22624
rect 2271 22593 2283 22596
rect 2225 22587 2283 22593
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 2958 22584 2964 22636
rect 3016 22584 3022 22636
rect 4338 22584 4344 22636
rect 4396 22584 4402 22636
rect 5258 22584 5264 22636
rect 5316 22624 5322 22636
rect 5736 22633 5764 22664
rect 5353 22627 5411 22633
rect 5353 22624 5365 22627
rect 5316 22596 5365 22624
rect 5316 22584 5322 22596
rect 5353 22593 5365 22596
rect 5399 22593 5411 22627
rect 5353 22587 5411 22593
rect 5537 22627 5595 22633
rect 5537 22593 5549 22627
rect 5583 22593 5595 22627
rect 5537 22587 5595 22593
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22593 5779 22627
rect 5721 22587 5779 22593
rect 2409 22559 2467 22565
rect 2409 22525 2421 22559
rect 2455 22556 2467 22559
rect 3326 22556 3332 22568
rect 2455 22528 3332 22556
rect 2455 22525 2467 22528
rect 2409 22519 2467 22525
rect 3326 22516 3332 22528
rect 3384 22516 3390 22568
rect 3694 22516 3700 22568
rect 3752 22556 3758 22568
rect 5074 22556 5080 22568
rect 3752 22528 5080 22556
rect 3752 22516 3758 22528
rect 5074 22516 5080 22528
rect 5132 22516 5138 22568
rect 5552 22556 5580 22587
rect 5810 22584 5816 22636
rect 5868 22584 5874 22636
rect 5920 22556 5948 22664
rect 6546 22652 6552 22664
rect 6604 22652 6610 22704
rect 6641 22695 6699 22701
rect 6641 22661 6653 22695
rect 6687 22692 6699 22695
rect 6687 22664 7237 22692
rect 6687 22661 6699 22664
rect 6641 22655 6699 22661
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6086 22584 6092 22636
rect 6144 22624 6150 22636
rect 6365 22627 6423 22633
rect 6365 22624 6377 22627
rect 6144 22596 6377 22624
rect 6144 22584 6150 22596
rect 6365 22593 6377 22596
rect 6411 22593 6423 22627
rect 6733 22627 6791 22633
rect 6733 22624 6745 22627
rect 6365 22587 6423 22593
rect 6656 22596 6745 22624
rect 6656 22556 6684 22596
rect 6733 22593 6745 22596
rect 6779 22593 6791 22627
rect 6733 22587 6791 22593
rect 5552 22528 5948 22556
rect 6012 22528 6684 22556
rect 4338 22448 4344 22500
rect 4396 22488 4402 22500
rect 5810 22488 5816 22500
rect 4396 22460 5816 22488
rect 4396 22448 4402 22460
rect 5810 22448 5816 22460
rect 5868 22448 5874 22500
rect 2593 22423 2651 22429
rect 2593 22389 2605 22423
rect 2639 22420 2651 22423
rect 4062 22420 4068 22432
rect 2639 22392 4068 22420
rect 2639 22389 2651 22392
rect 2593 22383 2651 22389
rect 4062 22380 4068 22392
rect 4120 22380 4126 22432
rect 4433 22423 4491 22429
rect 4433 22389 4445 22423
rect 4479 22420 4491 22423
rect 4706 22420 4712 22432
rect 4479 22392 4712 22420
rect 4479 22389 4491 22392
rect 4433 22383 4491 22389
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 5258 22380 5264 22432
rect 5316 22420 5322 22432
rect 6012 22420 6040 22528
rect 7098 22516 7104 22568
rect 7156 22516 7162 22568
rect 7209 22556 7237 22664
rect 7374 22652 7380 22704
rect 7432 22692 7438 22704
rect 8110 22692 8116 22704
rect 7432 22664 8116 22692
rect 7432 22652 7438 22664
rect 8110 22652 8116 22664
rect 8168 22652 8174 22704
rect 7834 22584 7840 22636
rect 7892 22584 7898 22636
rect 7985 22627 8043 22633
rect 7985 22593 7997 22627
rect 8031 22624 8043 22627
rect 8031 22596 8156 22624
rect 8031 22593 8043 22596
rect 7985 22587 8043 22593
rect 8128 22568 8156 22596
rect 8202 22584 8208 22636
rect 8260 22584 8266 22636
rect 8312 22633 8340 22732
rect 8481 22729 8493 22763
rect 8527 22760 8539 22763
rect 9861 22763 9919 22769
rect 8527 22732 9444 22760
rect 8527 22729 8539 22732
rect 8481 22723 8539 22729
rect 8941 22695 8999 22701
rect 8496 22664 8709 22692
rect 8302 22627 8360 22633
rect 8302 22593 8314 22627
rect 8348 22593 8360 22627
rect 8302 22587 8360 22593
rect 7650 22556 7656 22568
rect 7209 22528 7656 22556
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 8110 22516 8116 22568
rect 8168 22516 8174 22568
rect 6822 22448 6828 22500
rect 6880 22488 6886 22500
rect 8496 22488 8524 22664
rect 8681 22633 8709 22664
rect 8941 22661 8953 22695
rect 8987 22692 8999 22695
rect 9122 22692 9128 22704
rect 8987 22664 9128 22692
rect 8987 22661 8999 22664
rect 8941 22655 8999 22661
rect 9122 22652 9128 22664
rect 9180 22652 9186 22704
rect 9416 22701 9444 22732
rect 9861 22729 9873 22763
rect 9907 22760 9919 22763
rect 10042 22760 10048 22772
rect 9907 22732 10048 22760
rect 9907 22729 9919 22732
rect 9861 22723 9919 22729
rect 10042 22720 10048 22732
rect 10100 22720 10106 22772
rect 10226 22720 10232 22772
rect 10284 22720 10290 22772
rect 10318 22720 10324 22772
rect 10376 22720 10382 22772
rect 11330 22760 11336 22772
rect 11072 22732 11336 22760
rect 9401 22695 9459 22701
rect 9401 22661 9413 22695
rect 9447 22661 9459 22695
rect 9401 22655 9459 22661
rect 9766 22652 9772 22704
rect 9824 22652 9830 22704
rect 10962 22652 10968 22704
rect 11020 22652 11026 22704
rect 11072 22701 11100 22732
rect 11330 22720 11336 22732
rect 11388 22760 11394 22772
rect 11698 22760 11704 22772
rect 11388 22732 11704 22760
rect 11388 22720 11394 22732
rect 11698 22720 11704 22732
rect 11756 22720 11762 22772
rect 12158 22760 12164 22772
rect 12084 22732 12164 22760
rect 11057 22695 11115 22701
rect 11057 22661 11069 22695
rect 11103 22661 11115 22695
rect 11057 22655 11115 22661
rect 11882 22652 11888 22704
rect 11940 22652 11946 22704
rect 11977 22695 12035 22701
rect 11977 22661 11989 22695
rect 12023 22692 12035 22695
rect 12084 22692 12112 22732
rect 12158 22720 12164 22732
rect 12216 22720 12222 22772
rect 14001 22763 14059 22769
rect 14001 22760 14013 22763
rect 12268 22732 14013 22760
rect 12268 22692 12296 22732
rect 14001 22729 14013 22732
rect 14047 22729 14059 22763
rect 14001 22723 14059 22729
rect 14642 22720 14648 22772
rect 14700 22760 14706 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 14700 22732 14933 22760
rect 14700 22720 14706 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 14921 22723 14979 22729
rect 15286 22720 15292 22772
rect 15344 22760 15350 22772
rect 15930 22760 15936 22772
rect 15344 22732 15936 22760
rect 15344 22720 15350 22732
rect 15930 22720 15936 22732
rect 15988 22720 15994 22772
rect 16942 22720 16948 22772
rect 17000 22760 17006 22772
rect 17494 22760 17500 22772
rect 17000 22732 17500 22760
rect 17000 22720 17006 22732
rect 17494 22720 17500 22732
rect 17552 22720 17558 22772
rect 19702 22720 19708 22772
rect 19760 22760 19766 22772
rect 19889 22763 19947 22769
rect 19889 22760 19901 22763
rect 19760 22732 19901 22760
rect 19760 22720 19766 22732
rect 19889 22729 19901 22732
rect 19935 22729 19947 22763
rect 20625 22763 20683 22769
rect 20625 22760 20637 22763
rect 19889 22723 19947 22729
rect 20088 22732 20637 22760
rect 12023 22664 12112 22692
rect 12175 22664 12296 22692
rect 12023 22661 12035 22664
rect 11977 22655 12035 22661
rect 12175 22636 12203 22664
rect 12618 22652 12624 22704
rect 12676 22692 12682 22704
rect 12802 22692 12808 22704
rect 12676 22664 12808 22692
rect 12676 22652 12682 22664
rect 12802 22652 12808 22664
rect 12860 22692 12866 22704
rect 12897 22695 12955 22701
rect 12897 22692 12909 22695
rect 12860 22664 12909 22692
rect 12860 22652 12866 22664
rect 12897 22661 12909 22664
rect 12943 22661 12955 22695
rect 12897 22655 12955 22661
rect 13170 22652 13176 22704
rect 13228 22652 13234 22704
rect 13354 22652 13360 22704
rect 13412 22692 13418 22704
rect 14369 22695 14427 22701
rect 14369 22692 14381 22695
rect 13412 22664 13676 22692
rect 13412 22652 13418 22664
rect 8573 22627 8631 22633
rect 8573 22593 8585 22627
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 8666 22627 8724 22633
rect 8666 22593 8678 22627
rect 8712 22593 8724 22627
rect 8666 22587 8724 22593
rect 8849 22627 8907 22633
rect 8849 22593 8861 22627
rect 8895 22593 8907 22627
rect 8849 22587 8907 22593
rect 8576 22586 8616 22587
rect 8576 22500 8604 22586
rect 8864 22556 8892 22587
rect 9030 22584 9036 22636
rect 9088 22633 9094 22636
rect 9088 22624 9096 22633
rect 9585 22627 9643 22633
rect 9585 22624 9597 22627
rect 9088 22596 9597 22624
rect 9088 22587 9096 22596
rect 9585 22593 9597 22596
rect 9631 22593 9643 22627
rect 9585 22587 9643 22593
rect 9088 22584 9094 22587
rect 9398 22556 9404 22568
rect 8864 22528 9404 22556
rect 9398 22516 9404 22528
rect 9456 22516 9462 22568
rect 6880 22460 8524 22488
rect 6880 22448 6886 22460
rect 8570 22448 8576 22500
rect 8628 22448 8634 22500
rect 9122 22448 9128 22500
rect 9180 22488 9186 22500
rect 9217 22491 9275 22497
rect 9217 22488 9229 22491
rect 9180 22460 9229 22488
rect 9180 22448 9186 22460
rect 9217 22457 9229 22460
rect 9263 22457 9275 22491
rect 9600 22488 9628 22587
rect 9674 22584 9680 22636
rect 9732 22624 9738 22636
rect 10827 22627 10885 22633
rect 10827 22624 10839 22627
rect 9732 22596 10839 22624
rect 9732 22584 9738 22596
rect 10827 22593 10839 22596
rect 10873 22593 10885 22627
rect 11149 22627 11207 22633
rect 11149 22624 11161 22627
rect 10827 22587 10885 22593
rect 10980 22596 11161 22624
rect 10980 22568 11008 22596
rect 11149 22593 11161 22596
rect 11195 22593 11207 22627
rect 11149 22587 11207 22593
rect 11698 22584 11704 22636
rect 11756 22633 11762 22636
rect 11756 22627 11805 22633
rect 11756 22593 11759 22627
rect 11793 22593 11805 22627
rect 11756 22587 11805 22593
rect 11756 22584 11762 22587
rect 12158 22584 12164 22636
rect 12216 22584 12222 22636
rect 12253 22627 12311 22633
rect 12253 22593 12265 22627
rect 12299 22593 12311 22627
rect 13446 22624 13452 22636
rect 13407 22596 13452 22624
rect 12253 22587 12311 22593
rect 10410 22516 10416 22568
rect 10468 22516 10474 22568
rect 10686 22516 10692 22568
rect 10744 22516 10750 22568
rect 10962 22516 10968 22568
rect 11020 22516 11026 22568
rect 11974 22516 11980 22568
rect 12032 22556 12038 22568
rect 12268 22556 12296 22587
rect 13446 22584 13452 22596
rect 13504 22584 13510 22636
rect 13538 22584 13544 22636
rect 13596 22584 13602 22636
rect 13648 22633 13676 22664
rect 13832 22664 14381 22692
rect 13832 22633 13860 22664
rect 14369 22661 14381 22664
rect 14415 22661 14427 22695
rect 14369 22655 14427 22661
rect 14553 22695 14611 22701
rect 14553 22661 14565 22695
rect 14599 22692 14611 22695
rect 14734 22692 14740 22704
rect 14599 22664 14740 22692
rect 14599 22661 14611 22664
rect 14553 22655 14611 22661
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 13817 22627 13875 22633
rect 13817 22593 13829 22627
rect 13863 22593 13875 22627
rect 13817 22587 13875 22593
rect 14001 22627 14059 22633
rect 14001 22593 14013 22627
rect 14047 22593 14059 22627
rect 14001 22587 14059 22593
rect 12032 22528 12296 22556
rect 12032 22516 12038 22528
rect 13722 22516 13728 22568
rect 13780 22556 13786 22568
rect 14016 22556 14044 22587
rect 14274 22584 14280 22636
rect 14332 22584 14338 22636
rect 13780 22528 14044 22556
rect 14384 22556 14412 22655
rect 14734 22652 14740 22664
rect 14792 22652 14798 22704
rect 15120 22664 16160 22692
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 15120 22633 15148 22664
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 15565 22627 15623 22633
rect 15565 22593 15577 22627
rect 15611 22624 15623 22627
rect 15746 22624 15752 22636
rect 15611 22596 15752 22624
rect 15611 22593 15623 22596
rect 15565 22587 15623 22593
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 16132 22633 16160 22664
rect 17862 22652 17868 22704
rect 17920 22692 17926 22704
rect 19334 22692 19340 22704
rect 17920 22664 19340 22692
rect 17920 22652 17926 22664
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22624 15991 22627
rect 16117 22627 16175 22633
rect 15979 22596 16068 22624
rect 15979 22593 15991 22596
rect 15933 22587 15991 22593
rect 14826 22556 14832 22568
rect 14384 22528 14832 22556
rect 13780 22516 13786 22528
rect 14826 22516 14832 22528
rect 14884 22516 14890 22568
rect 15197 22559 15255 22565
rect 15197 22525 15209 22559
rect 15243 22556 15255 22559
rect 15286 22556 15292 22568
rect 15243 22528 15292 22556
rect 15243 22525 15255 22528
rect 15197 22519 15255 22525
rect 15286 22516 15292 22528
rect 15344 22516 15350 22568
rect 15473 22559 15531 22565
rect 15473 22525 15485 22559
rect 15519 22525 15531 22559
rect 16040 22556 16068 22596
rect 16117 22593 16129 22627
rect 16163 22624 16175 22627
rect 17954 22624 17960 22636
rect 16163 22596 17960 22624
rect 16163 22593 16175 22596
rect 16117 22587 16175 22593
rect 17954 22584 17960 22596
rect 18012 22584 18018 22636
rect 18230 22584 18236 22636
rect 18288 22584 18294 22636
rect 18414 22584 18420 22636
rect 18472 22584 18478 22636
rect 18509 22627 18567 22633
rect 18509 22593 18521 22627
rect 18555 22624 18567 22627
rect 19426 22624 19432 22636
rect 18555 22596 19432 22624
rect 18555 22593 18567 22596
rect 18509 22587 18567 22593
rect 19426 22584 19432 22596
rect 19484 22584 19490 22636
rect 20088 22633 20116 22732
rect 20625 22729 20637 22732
rect 20671 22729 20683 22763
rect 20625 22723 20683 22729
rect 22830 22720 22836 22772
rect 22888 22760 22894 22772
rect 23385 22763 23443 22769
rect 23385 22760 23397 22763
rect 22888 22732 23397 22760
rect 22888 22720 22894 22732
rect 23385 22729 23397 22732
rect 23431 22729 23443 22763
rect 23385 22723 23443 22729
rect 25406 22720 25412 22772
rect 25464 22720 25470 22772
rect 25590 22720 25596 22772
rect 25648 22720 25654 22772
rect 32582 22760 32588 22772
rect 32416 22732 32588 22760
rect 20898 22692 20904 22704
rect 20272 22664 20904 22692
rect 20073 22627 20131 22633
rect 20073 22593 20085 22627
rect 20119 22593 20131 22627
rect 20073 22587 20131 22593
rect 16482 22556 16488 22568
rect 16040 22528 16488 22556
rect 15473 22519 15531 22525
rect 10502 22488 10508 22500
rect 9600 22460 10508 22488
rect 9217 22451 9275 22457
rect 10502 22448 10508 22460
rect 10560 22448 10566 22500
rect 11256 22460 11744 22488
rect 5316 22392 6040 22420
rect 5316 22380 5322 22392
rect 6086 22380 6092 22432
rect 6144 22420 6150 22432
rect 6362 22420 6368 22432
rect 6144 22392 6368 22420
rect 6144 22380 6150 22392
rect 6362 22380 6368 22392
rect 6420 22380 6426 22432
rect 8202 22380 8208 22432
rect 8260 22420 8266 22432
rect 11256 22420 11284 22460
rect 8260 22392 11284 22420
rect 11333 22423 11391 22429
rect 8260 22380 8266 22392
rect 11333 22389 11345 22423
rect 11379 22420 11391 22423
rect 11514 22420 11520 22432
rect 11379 22392 11520 22420
rect 11379 22389 11391 22392
rect 11333 22383 11391 22389
rect 11514 22380 11520 22392
rect 11572 22380 11578 22432
rect 11606 22380 11612 22432
rect 11664 22380 11670 22432
rect 11716 22420 11744 22460
rect 12342 22448 12348 22500
rect 12400 22488 12406 22500
rect 12437 22491 12495 22497
rect 12437 22488 12449 22491
rect 12400 22460 12449 22488
rect 12400 22448 12406 22460
rect 12437 22457 12449 22460
rect 12483 22457 12495 22491
rect 12437 22451 12495 22457
rect 12526 22448 12532 22500
rect 12584 22488 12590 22500
rect 14369 22491 14427 22497
rect 14369 22488 14381 22491
rect 12584 22460 14381 22488
rect 12584 22448 12590 22460
rect 14369 22457 14381 22460
rect 14415 22457 14427 22491
rect 14369 22451 14427 22457
rect 15010 22448 15016 22500
rect 15068 22488 15074 22500
rect 15488 22488 15516 22519
rect 16482 22516 16488 22528
rect 16540 22516 16546 22568
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22556 18107 22559
rect 18322 22556 18328 22568
rect 18095 22528 18328 22556
rect 18095 22525 18107 22528
rect 18049 22519 18107 22525
rect 18322 22516 18328 22528
rect 18380 22516 18386 22568
rect 18598 22516 18604 22568
rect 18656 22556 18662 22568
rect 20088 22556 20116 22587
rect 18656 22528 20116 22556
rect 18656 22516 18662 22528
rect 15068 22460 15516 22488
rect 15068 22448 15074 22460
rect 18230 22448 18236 22500
rect 18288 22488 18294 22500
rect 20272 22488 20300 22664
rect 20898 22652 20904 22664
rect 20956 22652 20962 22704
rect 22554 22652 22560 22704
rect 22612 22652 22618 22704
rect 23198 22652 23204 22704
rect 23256 22692 23262 22704
rect 25608 22692 25636 22720
rect 32416 22701 32444 22732
rect 32582 22720 32588 22732
rect 32640 22720 32646 22772
rect 32674 22720 32680 22772
rect 32732 22720 32738 22772
rect 32769 22763 32827 22769
rect 32769 22729 32781 22763
rect 32815 22729 32827 22763
rect 32769 22723 32827 22729
rect 35897 22763 35955 22769
rect 35897 22729 35909 22763
rect 35943 22760 35955 22763
rect 36262 22760 36268 22772
rect 35943 22732 36268 22760
rect 35943 22729 35955 22732
rect 35897 22723 35955 22729
rect 23256 22664 24532 22692
rect 23256 22652 23262 22664
rect 20530 22584 20536 22636
rect 20588 22584 20594 22636
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 22281 22627 22339 22633
rect 22281 22593 22293 22627
rect 22327 22624 22339 22627
rect 22646 22624 22652 22636
rect 22327 22596 22652 22624
rect 22327 22593 22339 22596
rect 22281 22587 22339 22593
rect 22646 22584 22652 22596
rect 22704 22584 22710 22636
rect 23474 22584 23480 22636
rect 23532 22624 23538 22636
rect 23569 22627 23627 22633
rect 23569 22624 23581 22627
rect 23532 22596 23581 22624
rect 23532 22584 23538 22596
rect 23569 22593 23581 22596
rect 23615 22593 23627 22627
rect 23569 22587 23627 22593
rect 23750 22584 23756 22636
rect 23808 22584 23814 22636
rect 23934 22584 23940 22636
rect 23992 22633 23998 22636
rect 23992 22627 24041 22633
rect 23992 22593 23995 22627
rect 24029 22593 24041 22627
rect 23992 22587 24041 22593
rect 23992 22584 23998 22587
rect 24118 22584 24124 22636
rect 24176 22584 24182 22636
rect 24210 22584 24216 22636
rect 24268 22584 24274 22636
rect 24394 22584 24400 22636
rect 24452 22584 24458 22636
rect 24504 22633 24532 22664
rect 25332 22664 25636 22692
rect 32401 22695 32459 22701
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22593 24547 22627
rect 24489 22587 24547 22593
rect 20349 22559 20407 22565
rect 20349 22525 20361 22559
rect 20395 22525 20407 22559
rect 23768 22556 23796 22584
rect 24302 22556 24308 22568
rect 23768 22528 24308 22556
rect 20349 22519 20407 22525
rect 18288 22460 20300 22488
rect 20364 22488 20392 22519
rect 24302 22516 24308 22528
rect 24360 22516 24366 22568
rect 21913 22491 21971 22497
rect 21913 22488 21925 22491
rect 20364 22460 21925 22488
rect 18288 22448 18294 22460
rect 21913 22457 21925 22460
rect 21959 22457 21971 22491
rect 25332 22488 25360 22664
rect 32401 22661 32413 22695
rect 32447 22661 32459 22695
rect 32401 22655 32459 22661
rect 32493 22695 32551 22701
rect 32493 22661 32505 22695
rect 32539 22692 32551 22695
rect 32692 22692 32720 22720
rect 32539 22664 32720 22692
rect 32784 22692 32812 22723
rect 36262 22720 36268 22732
rect 36320 22720 36326 22772
rect 33042 22692 33048 22704
rect 32784 22664 33048 22692
rect 32539 22661 32551 22664
rect 32493 22655 32551 22661
rect 33042 22652 33048 22664
rect 33100 22692 33106 22704
rect 33100 22664 33456 22692
rect 33100 22652 33106 22664
rect 25590 22584 25596 22636
rect 25648 22584 25654 22636
rect 25682 22584 25688 22636
rect 25740 22624 25746 22636
rect 27525 22627 27583 22633
rect 27525 22624 27537 22627
rect 25740 22596 27537 22624
rect 25740 22584 25746 22596
rect 27525 22593 27537 22596
rect 27571 22593 27583 22627
rect 27525 22587 27583 22593
rect 28074 22584 28080 22636
rect 28132 22624 28138 22636
rect 28445 22627 28503 22633
rect 28445 22624 28457 22627
rect 28132 22596 28457 22624
rect 28132 22584 28138 22596
rect 28445 22593 28457 22596
rect 28491 22593 28503 22627
rect 28445 22587 28503 22593
rect 28629 22627 28687 22633
rect 28629 22593 28641 22627
rect 28675 22624 28687 22627
rect 28718 22624 28724 22636
rect 28675 22596 28724 22624
rect 28675 22593 28687 22596
rect 28629 22587 28687 22593
rect 28718 22584 28724 22596
rect 28776 22584 28782 22636
rect 31846 22584 31852 22636
rect 31904 22624 31910 22636
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 31904 22596 32137 22624
rect 31904 22584 31910 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 32218 22627 32276 22633
rect 32218 22593 32230 22627
rect 32264 22593 32276 22627
rect 32629 22627 32687 22633
rect 32629 22624 32641 22627
rect 32218 22587 32276 22593
rect 32560 22596 32641 22624
rect 25406 22516 25412 22568
rect 25464 22556 25470 22568
rect 25777 22559 25835 22565
rect 25777 22556 25789 22559
rect 25464 22528 25789 22556
rect 25464 22516 25470 22528
rect 25777 22525 25789 22528
rect 25823 22556 25835 22559
rect 25866 22556 25872 22568
rect 25823 22528 25872 22556
rect 25823 22525 25835 22528
rect 25777 22519 25835 22525
rect 25866 22516 25872 22528
rect 25924 22516 25930 22568
rect 27798 22516 27804 22568
rect 27856 22516 27862 22568
rect 30834 22516 30840 22568
rect 30892 22556 30898 22568
rect 32232 22556 32260 22587
rect 30892 22528 32260 22556
rect 30892 22516 30898 22528
rect 25682 22488 25688 22500
rect 25332 22460 25688 22488
rect 21913 22451 21971 22457
rect 25682 22448 25688 22460
rect 25740 22448 25746 22500
rect 30742 22448 30748 22500
rect 30800 22488 30806 22500
rect 32560 22488 32588 22596
rect 32629 22593 32641 22596
rect 32675 22593 32687 22627
rect 32629 22587 32687 22593
rect 32766 22584 32772 22636
rect 32824 22624 32830 22636
rect 33428 22633 33456 22664
rect 33321 22627 33379 22633
rect 33321 22624 33333 22627
rect 32824 22596 33333 22624
rect 32824 22584 32830 22596
rect 33321 22593 33333 22596
rect 33367 22593 33379 22627
rect 33321 22587 33379 22593
rect 33413 22627 33471 22633
rect 33413 22593 33425 22627
rect 33459 22593 33471 22627
rect 33413 22587 33471 22593
rect 34517 22627 34575 22633
rect 34517 22593 34529 22627
rect 34563 22624 34575 22627
rect 34698 22624 34704 22636
rect 34563 22596 34704 22624
rect 34563 22593 34575 22596
rect 34517 22587 34575 22593
rect 34698 22584 34704 22596
rect 34756 22584 34762 22636
rect 34790 22584 34796 22636
rect 34848 22584 34854 22636
rect 36078 22584 36084 22636
rect 36136 22584 36142 22636
rect 34606 22516 34612 22568
rect 34664 22516 34670 22568
rect 30800 22460 32588 22488
rect 32692 22460 34560 22488
rect 30800 22448 30806 22460
rect 13078 22420 13084 22432
rect 11716 22392 13084 22420
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 15562 22380 15568 22432
rect 15620 22420 15626 22432
rect 15749 22423 15807 22429
rect 15749 22420 15761 22423
rect 15620 22392 15761 22420
rect 15620 22380 15626 22392
rect 15749 22389 15761 22392
rect 15795 22389 15807 22423
rect 15749 22383 15807 22389
rect 16482 22380 16488 22432
rect 16540 22420 16546 22432
rect 19886 22420 19892 22432
rect 16540 22392 19892 22420
rect 16540 22380 16546 22392
rect 19886 22380 19892 22392
rect 19944 22380 19950 22432
rect 20257 22423 20315 22429
rect 20257 22389 20269 22423
rect 20303 22420 20315 22423
rect 20346 22420 20352 22432
rect 20303 22392 20352 22420
rect 20303 22389 20315 22392
rect 20257 22383 20315 22389
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 22462 22380 22468 22432
rect 22520 22380 22526 22432
rect 23750 22380 23756 22432
rect 23808 22380 23814 22432
rect 23845 22423 23903 22429
rect 23845 22389 23857 22423
rect 23891 22420 23903 22423
rect 23934 22420 23940 22432
rect 23891 22392 23940 22420
rect 23891 22389 23903 22392
rect 23845 22383 23903 22389
rect 23934 22380 23940 22392
rect 23992 22380 23998 22432
rect 27614 22380 27620 22432
rect 27672 22420 27678 22432
rect 28445 22423 28503 22429
rect 28445 22420 28457 22423
rect 27672 22392 28457 22420
rect 27672 22380 27678 22392
rect 28445 22389 28457 22392
rect 28491 22389 28503 22423
rect 28445 22383 28503 22389
rect 30282 22380 30288 22432
rect 30340 22420 30346 22432
rect 32692 22420 32720 22460
rect 33520 22429 33548 22460
rect 30340 22392 32720 22420
rect 33505 22423 33563 22429
rect 30340 22380 30346 22392
rect 33505 22389 33517 22423
rect 33551 22389 33563 22423
rect 33505 22383 33563 22389
rect 33686 22380 33692 22432
rect 33744 22380 33750 22432
rect 34532 22429 34560 22460
rect 34517 22423 34575 22429
rect 34517 22389 34529 22423
rect 34563 22389 34575 22423
rect 34517 22383 34575 22389
rect 34790 22380 34796 22432
rect 34848 22420 34854 22432
rect 34977 22423 35035 22429
rect 34977 22420 34989 22423
rect 34848 22392 34989 22420
rect 34848 22380 34854 22392
rect 34977 22389 34989 22392
rect 35023 22389 35035 22423
rect 34977 22383 35035 22389
rect 1104 22330 36432 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 36432 22330
rect 1104 22256 36432 22278
rect 1670 22176 1676 22228
rect 1728 22216 1734 22228
rect 2317 22219 2375 22225
rect 2317 22216 2329 22219
rect 1728 22188 2329 22216
rect 1728 22176 1734 22188
rect 2317 22185 2329 22188
rect 2363 22185 2375 22219
rect 2317 22179 2375 22185
rect 4433 22219 4491 22225
rect 4433 22185 4445 22219
rect 4479 22216 4491 22219
rect 4614 22216 4620 22228
rect 4479 22188 4620 22216
rect 4479 22185 4491 22188
rect 4433 22179 4491 22185
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 5445 22219 5503 22225
rect 5445 22185 5457 22219
rect 5491 22216 5503 22219
rect 5718 22216 5724 22228
rect 5491 22188 5724 22216
rect 5491 22185 5503 22188
rect 5445 22179 5503 22185
rect 5718 22176 5724 22188
rect 5776 22176 5782 22228
rect 6546 22176 6552 22228
rect 6604 22216 6610 22228
rect 9296 22219 9354 22225
rect 6604 22188 8800 22216
rect 6604 22176 6610 22188
rect 8772 22160 8800 22188
rect 9296 22185 9308 22219
rect 9342 22216 9354 22219
rect 9674 22216 9680 22228
rect 9342 22188 9680 22216
rect 9342 22185 9354 22188
rect 9296 22179 9354 22185
rect 9674 22176 9680 22188
rect 9732 22176 9738 22228
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 11790 22216 11796 22228
rect 10008 22188 11796 22216
rect 10008 22176 10014 22188
rect 11790 22176 11796 22188
rect 11848 22216 11854 22228
rect 12342 22216 12348 22228
rect 11848 22188 12348 22216
rect 11848 22176 11854 22188
rect 12342 22176 12348 22188
rect 12400 22176 12406 22228
rect 13357 22219 13415 22225
rect 13357 22185 13369 22219
rect 13403 22216 13415 22219
rect 13538 22216 13544 22228
rect 13403 22188 13544 22216
rect 13403 22185 13415 22188
rect 13357 22179 13415 22185
rect 13538 22176 13544 22188
rect 13596 22216 13602 22228
rect 13596 22188 13676 22216
rect 13596 22176 13602 22188
rect 2682 22108 2688 22160
rect 2740 22148 2746 22160
rect 2740 22120 3004 22148
rect 2740 22108 2746 22120
rect 2774 22040 2780 22092
rect 2832 22040 2838 22092
rect 2976 22089 3004 22120
rect 5074 22108 5080 22160
rect 5132 22148 5138 22160
rect 5534 22148 5540 22160
rect 5132 22120 5540 22148
rect 5132 22108 5138 22120
rect 5534 22108 5540 22120
rect 5592 22108 5598 22160
rect 7926 22108 7932 22160
rect 7984 22148 7990 22160
rect 7984 22120 8248 22148
rect 7984 22108 7990 22120
rect 8220 22092 8248 22120
rect 8754 22108 8760 22160
rect 8812 22148 8818 22160
rect 11057 22151 11115 22157
rect 8812 22120 9076 22148
rect 8812 22108 8818 22120
rect 2961 22083 3019 22089
rect 2961 22049 2973 22083
rect 3007 22080 3019 22083
rect 3326 22080 3332 22092
rect 3007 22052 3332 22080
rect 3007 22049 3019 22052
rect 2961 22043 3019 22049
rect 3326 22040 3332 22052
rect 3384 22040 3390 22092
rect 3881 22083 3939 22089
rect 3881 22049 3893 22083
rect 3927 22080 3939 22083
rect 4062 22080 4068 22092
rect 3927 22052 4068 22080
rect 3927 22049 3939 22052
rect 3881 22043 3939 22049
rect 4062 22040 4068 22052
rect 4120 22040 4126 22092
rect 5166 22040 5172 22092
rect 5224 22080 5230 22092
rect 5224 22052 5488 22080
rect 5224 22040 5230 22052
rect 4614 21972 4620 22024
rect 4672 22012 4678 22024
rect 4893 22015 4951 22021
rect 4893 22012 4905 22015
rect 4672 21984 4905 22012
rect 4672 21972 4678 21984
rect 4893 21981 4905 21984
rect 4939 21981 4951 22015
rect 4893 21975 4951 21981
rect 5258 21972 5264 22024
rect 5316 21972 5322 22024
rect 2685 21947 2743 21953
rect 2685 21913 2697 21947
rect 2731 21944 2743 21947
rect 4706 21944 4712 21956
rect 2731 21916 4712 21944
rect 2731 21913 2743 21916
rect 2685 21907 2743 21913
rect 4706 21904 4712 21916
rect 4764 21904 4770 21956
rect 4798 21904 4804 21956
rect 4856 21944 4862 21956
rect 5077 21947 5135 21953
rect 5077 21944 5089 21947
rect 4856 21916 5089 21944
rect 4856 21904 4862 21916
rect 5077 21913 5089 21916
rect 5123 21913 5135 21947
rect 5077 21907 5135 21913
rect 5169 21947 5227 21953
rect 5169 21913 5181 21947
rect 5215 21913 5227 21947
rect 5460 21944 5488 22052
rect 5902 22040 5908 22092
rect 5960 22080 5966 22092
rect 6917 22083 6975 22089
rect 6917 22080 6929 22083
rect 5960 22052 6929 22080
rect 5960 22040 5966 22052
rect 6917 22049 6929 22052
rect 6963 22080 6975 22083
rect 6963 22052 7972 22080
rect 6963 22049 6975 22052
rect 6917 22043 6975 22049
rect 7944 22024 7972 22052
rect 8202 22040 8208 22092
rect 8260 22040 8266 22092
rect 8478 22040 8484 22092
rect 8536 22080 8542 22092
rect 8938 22080 8944 22092
rect 8536 22052 8944 22080
rect 8536 22040 8542 22052
rect 8938 22040 8944 22052
rect 8996 22040 9002 22092
rect 9048 22080 9076 22120
rect 11057 22117 11069 22151
rect 11103 22117 11115 22151
rect 11057 22111 11115 22117
rect 11072 22080 11100 22111
rect 12802 22108 12808 22160
rect 12860 22148 12866 22160
rect 12989 22151 13047 22157
rect 12989 22148 13001 22151
rect 12860 22120 13001 22148
rect 12860 22108 12866 22120
rect 12989 22117 13001 22120
rect 13035 22117 13047 22151
rect 12989 22111 13047 22117
rect 9048 22052 11100 22080
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 13648 22080 13676 22188
rect 13814 22176 13820 22228
rect 13872 22176 13878 22228
rect 14936 22188 16988 22216
rect 14826 22108 14832 22160
rect 14884 22108 14890 22160
rect 14936 22080 14964 22188
rect 15562 22148 15568 22160
rect 15488 22120 15568 22148
rect 12115 22052 12480 22080
rect 13648 22052 13860 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 6641 22015 6699 22021
rect 6641 21981 6653 22015
rect 6687 22012 6699 22015
rect 7098 22012 7104 22024
rect 6687 21984 7104 22012
rect 6687 21981 6699 21984
rect 6641 21975 6699 21981
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 7466 21972 7472 22024
rect 7524 21972 7530 22024
rect 7926 21972 7932 22024
rect 7984 21972 7990 22024
rect 8294 21972 8300 22024
rect 8352 22012 8358 22024
rect 9033 22015 9091 22021
rect 9033 22012 9045 22015
rect 8352 21984 9045 22012
rect 8352 21972 8358 21984
rect 9033 21981 9045 21984
rect 9079 21981 9091 22015
rect 9033 21975 9091 21981
rect 10962 21972 10968 22024
rect 11020 22012 11026 22024
rect 11241 22015 11299 22021
rect 11241 22012 11253 22015
rect 11020 21984 11253 22012
rect 11020 21972 11026 21984
rect 11241 21981 11253 21984
rect 11287 21981 11299 22015
rect 11241 21975 11299 21981
rect 6454 21944 6460 21956
rect 5460 21916 6460 21944
rect 5169 21907 5227 21913
rect 5184 21876 5212 21907
rect 6454 21904 6460 21916
rect 6512 21944 6518 21956
rect 6733 21947 6791 21953
rect 6733 21944 6745 21947
rect 6512 21916 6745 21944
rect 6512 21904 6518 21916
rect 6733 21913 6745 21916
rect 6779 21913 6791 21947
rect 6733 21907 6791 21913
rect 5258 21876 5264 21888
rect 5184 21848 5264 21876
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 6273 21879 6331 21885
rect 6273 21845 6285 21879
rect 6319 21876 6331 21879
rect 6546 21876 6552 21888
rect 6319 21848 6552 21876
rect 6319 21845 6331 21848
rect 6273 21839 6331 21845
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 7484 21876 7512 21972
rect 8018 21904 8024 21956
rect 8076 21944 8082 21956
rect 8570 21944 8576 21956
rect 8076 21916 8576 21944
rect 8076 21904 8082 21916
rect 8570 21904 8576 21916
rect 8628 21904 8634 21956
rect 9766 21904 9772 21956
rect 9824 21904 9830 21956
rect 10594 21876 10600 21888
rect 7484 21848 10600 21876
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 10781 21879 10839 21885
rect 10781 21845 10793 21879
rect 10827 21876 10839 21879
rect 11146 21876 11152 21888
rect 10827 21848 11152 21876
rect 10827 21845 10839 21848
rect 10781 21839 10839 21845
rect 11146 21836 11152 21848
rect 11204 21836 11210 21888
rect 11256 21876 11284 21975
rect 11330 21972 11336 22024
rect 11388 21972 11394 22024
rect 11514 21972 11520 22024
rect 11572 21972 11578 22024
rect 11606 21972 11612 22024
rect 11664 21972 11670 22024
rect 11790 21972 11796 22024
rect 11848 21972 11854 22024
rect 11974 21972 11980 22024
rect 12032 21972 12038 22024
rect 12452 22021 12480 22052
rect 12437 22015 12495 22021
rect 12437 21981 12449 22015
rect 12483 21981 12495 22015
rect 12437 21975 12495 21981
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 22012 12771 22015
rect 12894 22012 12900 22024
rect 12759 21984 12900 22012
rect 12759 21981 12771 21984
rect 12713 21975 12771 21981
rect 11885 21947 11943 21953
rect 11885 21913 11897 21947
rect 11931 21944 11943 21947
rect 12158 21944 12164 21956
rect 11931 21916 12164 21944
rect 11931 21913 11943 21916
rect 11885 21907 11943 21913
rect 12158 21904 12164 21916
rect 12216 21904 12222 21956
rect 12253 21947 12311 21953
rect 12253 21913 12265 21947
rect 12299 21944 12311 21947
rect 12342 21944 12348 21956
rect 12299 21916 12348 21944
rect 12299 21913 12311 21916
rect 12253 21907 12311 21913
rect 12342 21904 12348 21916
rect 12400 21904 12406 21956
rect 12636 21944 12664 21975
rect 12894 21972 12900 21984
rect 12952 21972 12958 22024
rect 13173 22015 13231 22021
rect 13173 21981 13185 22015
rect 13219 22012 13231 22015
rect 13354 22012 13360 22024
rect 13219 21984 13360 22012
rect 13219 21981 13231 21984
rect 13173 21975 13231 21981
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13446 21972 13452 22024
rect 13504 22012 13510 22024
rect 13832 22021 13860 22052
rect 14660 22052 14964 22080
rect 15197 22083 15255 22089
rect 13541 22015 13599 22021
rect 13541 22012 13553 22015
rect 13504 21984 13553 22012
rect 13504 21972 13510 21984
rect 13541 21981 13553 21984
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 21981 13783 22015
rect 13725 21975 13783 21981
rect 13817 22015 13875 22021
rect 13817 21981 13829 22015
rect 13863 22012 13875 22015
rect 14660 22012 14688 22052
rect 15197 22049 15209 22083
rect 15243 22080 15255 22083
rect 15381 22083 15439 22089
rect 15381 22080 15393 22083
rect 15243 22052 15393 22080
rect 15243 22049 15255 22052
rect 15197 22043 15255 22049
rect 15381 22049 15393 22052
rect 15427 22049 15439 22083
rect 15381 22043 15439 22049
rect 13863 21984 14688 22012
rect 13863 21981 13875 21984
rect 13817 21975 13875 21981
rect 13262 21944 13268 21956
rect 12636 21916 13268 21944
rect 13262 21904 13268 21916
rect 13320 21904 13326 21956
rect 13740 21944 13768 21975
rect 14734 21972 14740 22024
rect 14792 22012 14798 22024
rect 15013 22015 15071 22021
rect 15013 22012 15025 22015
rect 14792 21984 15025 22012
rect 14792 21972 14798 21984
rect 15013 21981 15025 21984
rect 15059 21981 15071 22015
rect 15013 21975 15071 21981
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 22012 15347 22015
rect 15488 22012 15516 22120
rect 15562 22108 15568 22120
rect 15620 22148 15626 22160
rect 15620 22120 16344 22148
rect 15620 22108 15626 22120
rect 15746 22040 15752 22092
rect 15804 22080 15810 22092
rect 16316 22080 16344 22120
rect 16853 22083 16911 22089
rect 16853 22080 16865 22083
rect 15804 22052 16252 22080
rect 16316 22052 16865 22080
rect 15804 22040 15810 22052
rect 15335 21984 15516 22012
rect 15335 21981 15347 21984
rect 15289 21975 15347 21981
rect 15562 21972 15568 22024
rect 15620 21972 15626 22024
rect 16224 22022 16252 22052
rect 16853 22049 16865 22052
rect 16899 22049 16911 22083
rect 16960 22080 16988 22188
rect 17218 22176 17224 22228
rect 17276 22176 17282 22228
rect 17954 22176 17960 22228
rect 18012 22216 18018 22228
rect 18012 22188 22094 22216
rect 18012 22176 18018 22188
rect 17310 22108 17316 22160
rect 17368 22148 17374 22160
rect 17405 22151 17463 22157
rect 17405 22148 17417 22151
rect 17368 22120 17417 22148
rect 17368 22108 17374 22120
rect 17405 22117 17417 22120
rect 17451 22117 17463 22151
rect 17405 22111 17463 22117
rect 19886 22108 19892 22160
rect 19944 22148 19950 22160
rect 20714 22148 20720 22160
rect 19944 22120 20720 22148
rect 19944 22108 19950 22120
rect 20714 22108 20720 22120
rect 20772 22148 20778 22160
rect 21082 22148 21088 22160
rect 20772 22120 21088 22148
rect 20772 22108 20778 22120
rect 21082 22108 21088 22120
rect 21140 22108 21146 22160
rect 22066 22148 22094 22188
rect 22462 22176 22468 22228
rect 22520 22216 22526 22228
rect 23109 22219 23167 22225
rect 23109 22216 23121 22219
rect 22520 22188 23121 22216
rect 22520 22176 22526 22188
rect 23109 22185 23121 22188
rect 23155 22216 23167 22219
rect 23198 22216 23204 22228
rect 23155 22188 23204 22216
rect 23155 22185 23167 22188
rect 23109 22179 23167 22185
rect 23198 22176 23204 22188
rect 23256 22176 23262 22228
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 24578 22216 24584 22228
rect 23808 22188 24584 22216
rect 23808 22176 23814 22188
rect 24578 22176 24584 22188
rect 24636 22176 24642 22228
rect 35253 22219 35311 22225
rect 35253 22185 35265 22219
rect 35299 22216 35311 22219
rect 35299 22188 35388 22216
rect 35299 22185 35311 22188
rect 35253 22179 35311 22185
rect 23014 22148 23020 22160
rect 22066 22120 23020 22148
rect 23014 22108 23020 22120
rect 23072 22108 23078 22160
rect 19337 22083 19395 22089
rect 19337 22080 19349 22083
rect 16960 22052 19349 22080
rect 16853 22043 16911 22049
rect 19337 22049 19349 22052
rect 19383 22049 19395 22083
rect 19337 22043 19395 22049
rect 19521 22083 19579 22089
rect 19521 22049 19533 22083
rect 19567 22080 19579 22083
rect 21453 22083 21511 22089
rect 19567 22052 19932 22080
rect 19567 22049 19579 22052
rect 19521 22043 19579 22049
rect 19904 22024 19932 22052
rect 21453 22049 21465 22083
rect 21499 22080 21511 22083
rect 21910 22080 21916 22092
rect 21499 22052 21916 22080
rect 21499 22049 21511 22052
rect 21453 22043 21511 22049
rect 21910 22040 21916 22052
rect 21968 22040 21974 22092
rect 23201 22083 23259 22089
rect 23201 22049 23213 22083
rect 23247 22080 23259 22083
rect 23768 22080 23796 22176
rect 35360 22160 35388 22188
rect 25130 22108 25136 22160
rect 25188 22148 25194 22160
rect 25188 22120 27200 22148
rect 25188 22108 25194 22120
rect 23247 22052 23796 22080
rect 23247 22049 23259 22052
rect 23201 22043 23259 22049
rect 26050 22040 26056 22092
rect 26108 22040 26114 22092
rect 26326 22040 26332 22092
rect 26384 22080 26390 22092
rect 27062 22080 27068 22092
rect 26384 22052 27068 22080
rect 26384 22040 26390 22052
rect 27062 22040 27068 22052
rect 27120 22040 27126 22092
rect 27172 22024 27200 22120
rect 32122 22108 32128 22160
rect 32180 22148 32186 22160
rect 32674 22148 32680 22160
rect 32180 22120 32680 22148
rect 32180 22108 32186 22120
rect 32674 22108 32680 22120
rect 32732 22108 32738 22160
rect 35342 22108 35348 22160
rect 35400 22108 35406 22160
rect 27249 22083 27307 22089
rect 27249 22049 27261 22083
rect 27295 22080 27307 22083
rect 27614 22080 27620 22092
rect 27295 22052 27620 22080
rect 27295 22049 27307 22052
rect 27249 22043 27307 22049
rect 27614 22040 27620 22052
rect 27672 22040 27678 22092
rect 27893 22083 27951 22089
rect 27893 22049 27905 22083
rect 27939 22080 27951 22083
rect 30282 22080 30288 22092
rect 27939 22052 30288 22080
rect 27939 22049 27951 22052
rect 27893 22043 27951 22049
rect 30282 22040 30288 22052
rect 30340 22040 30346 22092
rect 30650 22040 30656 22092
rect 30708 22080 30714 22092
rect 35805 22083 35863 22089
rect 35805 22080 35817 22083
rect 30708 22052 35817 22080
rect 30708 22040 30714 22052
rect 35805 22049 35817 22052
rect 35851 22049 35863 22083
rect 35805 22043 35863 22049
rect 15841 22015 15899 22021
rect 15841 21981 15853 22015
rect 15887 21981 15899 22015
rect 15841 21975 15899 21981
rect 16117 22015 16175 22021
rect 16117 21981 16129 22015
rect 16163 21981 16175 22015
rect 16224 22012 16344 22022
rect 16482 22012 16488 22024
rect 16224 21994 16488 22012
rect 16316 21984 16488 21994
rect 16117 21975 16175 21981
rect 14826 21944 14832 21956
rect 13740 21916 14832 21944
rect 14826 21904 14832 21916
rect 14884 21904 14890 21956
rect 15746 21904 15752 21956
rect 15804 21944 15810 21956
rect 15856 21944 15884 21975
rect 15804 21916 15884 21944
rect 15804 21904 15810 21916
rect 13814 21876 13820 21888
rect 11256 21848 13820 21876
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 15838 21836 15844 21888
rect 15896 21876 15902 21888
rect 16025 21879 16083 21885
rect 16025 21876 16037 21879
rect 15896 21848 16037 21876
rect 15896 21836 15902 21848
rect 16025 21845 16037 21848
rect 16071 21845 16083 21879
rect 16132 21876 16160 21975
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 18414 21972 18420 22024
rect 18472 22012 18478 22024
rect 19613 22015 19671 22021
rect 18472 21984 19472 22012
rect 18472 21972 18478 21984
rect 16390 21904 16396 21956
rect 16448 21944 16454 21956
rect 19334 21944 19340 21956
rect 16448 21916 19340 21944
rect 16448 21904 16454 21916
rect 19334 21904 19340 21916
rect 19392 21904 19398 21956
rect 16206 21876 16212 21888
rect 16132 21848 16212 21876
rect 16025 21839 16083 21845
rect 16206 21836 16212 21848
rect 16264 21836 16270 21888
rect 17221 21879 17279 21885
rect 17221 21845 17233 21879
rect 17267 21876 17279 21879
rect 18782 21876 18788 21888
rect 17267 21848 18788 21876
rect 17267 21845 17279 21848
rect 17221 21839 17279 21845
rect 18782 21836 18788 21848
rect 18840 21836 18846 21888
rect 19444 21876 19472 21984
rect 19613 21981 19625 22015
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 19794 22012 19800 22024
rect 19751 21984 19800 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 19628 21944 19656 21975
rect 19794 21972 19800 21984
rect 19852 21972 19858 22024
rect 19886 21972 19892 22024
rect 19944 21972 19950 22024
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 22012 20131 22015
rect 21729 22015 21787 22021
rect 21729 22012 21741 22015
rect 20119 21984 21741 22012
rect 20119 21981 20131 21984
rect 20073 21975 20131 21981
rect 21729 21981 21741 21984
rect 21775 22012 21787 22015
rect 22094 22012 22100 22024
rect 21775 21984 22100 22012
rect 21775 21981 21787 21984
rect 21729 21975 21787 21981
rect 20088 21944 20116 21975
rect 22094 21972 22100 21984
rect 22152 22012 22158 22024
rect 22738 22012 22744 22024
rect 22152 21984 22744 22012
rect 22152 21972 22158 21984
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 23106 21972 23112 22024
rect 23164 22012 23170 22024
rect 23293 22015 23351 22021
rect 23293 22012 23305 22015
rect 23164 21984 23305 22012
rect 23164 21972 23170 21984
rect 23293 21981 23305 21984
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 23477 22015 23535 22021
rect 23477 21981 23489 22015
rect 23523 21981 23535 22015
rect 23477 21975 23535 21981
rect 19628 21916 20116 21944
rect 20254 21904 20260 21956
rect 20312 21944 20318 21956
rect 20990 21944 20996 21956
rect 20312 21916 20996 21944
rect 20312 21904 20318 21916
rect 20990 21904 20996 21916
rect 21048 21904 21054 21956
rect 21244 21947 21302 21953
rect 21244 21913 21256 21947
rect 21290 21944 21302 21947
rect 22833 21947 22891 21953
rect 22833 21944 22845 21947
rect 21290 21916 22845 21944
rect 21290 21913 21302 21916
rect 21244 21907 21302 21913
rect 22833 21913 22845 21916
rect 22879 21913 22891 21947
rect 23492 21944 23520 21975
rect 26234 21972 26240 22024
rect 26292 21972 26298 22024
rect 27154 21972 27160 22024
rect 27212 22012 27218 22024
rect 27525 22015 27583 22021
rect 27525 22012 27537 22015
rect 27212 21984 27537 22012
rect 27212 21972 27218 21984
rect 27525 21981 27537 21984
rect 27571 21981 27583 22015
rect 27525 21975 27583 21981
rect 27709 22015 27767 22021
rect 27709 21981 27721 22015
rect 27755 22012 27767 22015
rect 28166 22012 28172 22024
rect 27755 21984 28172 22012
rect 27755 21981 27767 21984
rect 27709 21975 27767 21981
rect 28166 21972 28172 21984
rect 28224 21972 28230 22024
rect 28261 22015 28319 22021
rect 28261 21981 28273 22015
rect 28307 22012 28319 22015
rect 28994 22012 29000 22024
rect 28307 21984 29000 22012
rect 28307 21981 28319 21984
rect 28261 21975 28319 21981
rect 23750 21944 23756 21956
rect 23492 21916 23756 21944
rect 22833 21907 22891 21913
rect 23750 21904 23756 21916
rect 23808 21904 23814 21956
rect 26970 21904 26976 21956
rect 27028 21944 27034 21956
rect 27387 21947 27445 21953
rect 27387 21944 27399 21947
rect 27028 21916 27399 21944
rect 27028 21904 27034 21916
rect 27387 21913 27399 21916
rect 27433 21913 27445 21947
rect 27387 21907 27445 21913
rect 27617 21947 27675 21953
rect 27617 21913 27629 21947
rect 27663 21913 27675 21947
rect 27617 21907 27675 21913
rect 19981 21879 20039 21885
rect 19981 21876 19993 21879
rect 19444 21848 19993 21876
rect 19981 21845 19993 21848
rect 20027 21845 20039 21879
rect 19981 21839 20039 21845
rect 20162 21836 20168 21888
rect 20220 21876 20226 21888
rect 21085 21879 21143 21885
rect 21085 21876 21097 21879
rect 20220 21848 21097 21876
rect 20220 21836 20226 21848
rect 21085 21845 21097 21848
rect 21131 21845 21143 21879
rect 21085 21839 21143 21845
rect 21361 21879 21419 21885
rect 21361 21845 21373 21879
rect 21407 21876 21419 21879
rect 22002 21876 22008 21888
rect 21407 21848 22008 21876
rect 21407 21845 21419 21848
rect 21361 21839 21419 21845
rect 22002 21836 22008 21848
rect 22060 21836 22066 21888
rect 22462 21836 22468 21888
rect 22520 21876 22526 21888
rect 25774 21876 25780 21888
rect 22520 21848 25780 21876
rect 22520 21836 22526 21848
rect 25774 21836 25780 21848
rect 25832 21836 25838 21888
rect 26234 21836 26240 21888
rect 26292 21876 26298 21888
rect 26418 21876 26424 21888
rect 26292 21848 26424 21876
rect 26292 21836 26298 21848
rect 26418 21836 26424 21848
rect 26476 21836 26482 21888
rect 27632 21876 27660 21907
rect 27798 21904 27804 21956
rect 27856 21944 27862 21956
rect 28276 21944 28304 21975
rect 28994 21972 29000 21984
rect 29052 21972 29058 22024
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 22012 30251 22015
rect 30561 22015 30619 22021
rect 30239 21984 30512 22012
rect 30239 21981 30251 21984
rect 30193 21975 30251 21981
rect 27856 21916 28304 21944
rect 27856 21904 27862 21916
rect 28534 21904 28540 21956
rect 28592 21944 28598 21956
rect 30285 21947 30343 21953
rect 30285 21944 30297 21947
rect 28592 21916 30297 21944
rect 28592 21904 28598 21916
rect 30285 21913 30297 21916
rect 30331 21913 30343 21947
rect 30285 21907 30343 21913
rect 30374 21904 30380 21956
rect 30432 21904 30438 21956
rect 30484 21944 30512 21984
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 33318 22012 33324 22024
rect 30607 21984 33324 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 33318 21972 33324 21984
rect 33376 21972 33382 22024
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 35161 22015 35219 22021
rect 35161 22012 35173 22015
rect 34848 21984 35173 22012
rect 34848 21972 34854 21984
rect 35161 21981 35173 21984
rect 35207 21981 35219 22015
rect 35161 21975 35219 21981
rect 35345 22015 35403 22021
rect 35345 21981 35357 22015
rect 35391 22012 35403 22015
rect 35986 22012 35992 22024
rect 35391 21984 35992 22012
rect 35391 21981 35403 21984
rect 35345 21975 35403 21981
rect 35986 21972 35992 21984
rect 36044 21972 36050 22024
rect 36078 21972 36084 22024
rect 36136 21972 36142 22024
rect 30742 21944 30748 21956
rect 30484 21916 30748 21944
rect 30742 21904 30748 21916
rect 30800 21904 30806 21956
rect 27706 21876 27712 21888
rect 27632 21848 27712 21876
rect 27706 21836 27712 21848
rect 27764 21836 27770 21888
rect 28077 21879 28135 21885
rect 28077 21845 28089 21879
rect 28123 21876 28135 21879
rect 28166 21876 28172 21888
rect 28123 21848 28172 21876
rect 28123 21845 28135 21848
rect 28077 21839 28135 21845
rect 28166 21836 28172 21848
rect 28224 21836 28230 21888
rect 30006 21836 30012 21888
rect 30064 21836 30070 21888
rect 34238 21836 34244 21888
rect 34296 21876 34302 21888
rect 35529 21879 35587 21885
rect 35529 21876 35541 21879
rect 34296 21848 35541 21876
rect 34296 21836 34302 21848
rect 35529 21845 35541 21848
rect 35575 21845 35587 21879
rect 35529 21839 35587 21845
rect 1104 21786 36432 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 36432 21786
rect 1104 21712 36432 21734
rect 4982 21672 4988 21684
rect 4264 21644 4988 21672
rect 2958 21604 2964 21616
rect 2898 21576 2964 21604
rect 2958 21564 2964 21576
rect 3016 21564 3022 21616
rect 3418 21564 3424 21616
rect 3476 21604 3482 21616
rect 4264 21613 4292 21644
rect 4982 21632 4988 21644
rect 5040 21632 5046 21684
rect 5810 21632 5816 21684
rect 5868 21672 5874 21684
rect 5868 21644 8340 21672
rect 5868 21632 5874 21644
rect 4249 21607 4307 21613
rect 3476 21576 4200 21604
rect 3476 21564 3482 21576
rect 4062 21496 4068 21548
rect 4120 21496 4126 21548
rect 4172 21536 4200 21576
rect 4249 21573 4261 21607
rect 4295 21573 4307 21607
rect 4249 21567 4307 21573
rect 4341 21539 4399 21545
rect 4341 21536 4353 21539
rect 4172 21508 4353 21536
rect 4341 21505 4353 21508
rect 4387 21505 4399 21539
rect 4341 21499 4399 21505
rect 4433 21539 4491 21545
rect 4433 21505 4445 21539
rect 4479 21536 4491 21539
rect 4706 21536 4712 21548
rect 4479 21508 4712 21536
rect 4479 21505 4491 21508
rect 4433 21499 4491 21505
rect 4706 21496 4712 21508
rect 4764 21536 4770 21548
rect 5350 21536 5356 21548
rect 4764 21508 5356 21536
rect 4764 21496 4770 21508
rect 5350 21496 5356 21508
rect 5408 21496 5414 21548
rect 6380 21545 6408 21644
rect 8312 21616 8340 21644
rect 8570 21632 8576 21684
rect 8628 21672 8634 21684
rect 8628 21644 11008 21672
rect 8628 21632 8634 21644
rect 6546 21564 6552 21616
rect 6604 21604 6610 21616
rect 6641 21607 6699 21613
rect 6641 21604 6653 21607
rect 6604 21576 6653 21604
rect 6604 21564 6610 21576
rect 6641 21573 6653 21576
rect 6687 21573 6699 21607
rect 6641 21567 6699 21573
rect 7098 21564 7104 21616
rect 7156 21564 7162 21616
rect 8294 21564 8300 21616
rect 8352 21604 8358 21616
rect 8352 21576 8984 21604
rect 8352 21564 8358 21576
rect 8386 21545 8392 21548
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 8384 21536 8392 21545
rect 8347 21508 8392 21536
rect 6365 21499 6423 21505
rect 8384 21499 8392 21508
rect 8386 21496 8392 21499
rect 8444 21496 8450 21548
rect 8481 21539 8539 21545
rect 8481 21505 8493 21539
rect 8527 21505 8539 21539
rect 8481 21499 8539 21505
rect 8573 21539 8631 21545
rect 8573 21505 8585 21539
rect 8619 21536 8631 21539
rect 8662 21536 8668 21548
rect 8619 21508 8668 21536
rect 8619 21505 8631 21508
rect 8573 21499 8631 21505
rect 1394 21428 1400 21480
rect 1452 21428 1458 21480
rect 1673 21471 1731 21477
rect 1673 21437 1685 21471
rect 1719 21468 1731 21471
rect 2130 21468 2136 21480
rect 1719 21440 2136 21468
rect 1719 21437 1731 21440
rect 1673 21431 1731 21437
rect 2130 21428 2136 21440
rect 2188 21428 2194 21480
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21468 3203 21471
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 3191 21440 3893 21468
rect 3191 21437 3203 21440
rect 3145 21431 3203 21437
rect 3881 21437 3893 21440
rect 3927 21468 3939 21471
rect 5258 21468 5264 21480
rect 3927 21440 5264 21468
rect 3927 21437 3939 21440
rect 3881 21431 3939 21437
rect 5258 21428 5264 21440
rect 5316 21428 5322 21480
rect 5534 21428 5540 21480
rect 5592 21468 5598 21480
rect 8496 21468 8524 21499
rect 8662 21496 8668 21508
rect 8720 21496 8726 21548
rect 8754 21496 8760 21548
rect 8812 21496 8818 21548
rect 8956 21545 8984 21576
rect 9766 21564 9772 21616
rect 9824 21564 9830 21616
rect 10980 21613 11008 21644
rect 11146 21632 11152 21684
rect 11204 21632 11210 21684
rect 11330 21632 11336 21684
rect 11388 21672 11394 21684
rect 12437 21675 12495 21681
rect 12437 21672 12449 21675
rect 11388 21644 12449 21672
rect 11388 21632 11394 21644
rect 12437 21641 12449 21644
rect 12483 21641 12495 21675
rect 12437 21635 12495 21641
rect 12605 21675 12663 21681
rect 12605 21641 12617 21675
rect 12651 21672 12663 21675
rect 12710 21672 12716 21684
rect 12651 21644 12716 21672
rect 12651 21641 12663 21644
rect 12605 21635 12663 21641
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 13262 21632 13268 21684
rect 13320 21672 13326 21684
rect 13633 21675 13691 21681
rect 13633 21672 13645 21675
rect 13320 21644 13645 21672
rect 13320 21632 13326 21644
rect 13633 21641 13645 21644
rect 13679 21641 13691 21675
rect 13633 21635 13691 21641
rect 17218 21632 17224 21684
rect 17276 21672 17282 21684
rect 17497 21675 17555 21681
rect 17497 21672 17509 21675
rect 17276 21644 17509 21672
rect 17276 21632 17282 21644
rect 17497 21641 17509 21644
rect 17543 21641 17555 21675
rect 18877 21675 18935 21681
rect 17497 21635 17555 21641
rect 17604 21644 18736 21672
rect 10965 21607 11023 21613
rect 10965 21573 10977 21607
rect 11011 21573 11023 21607
rect 10965 21567 11023 21573
rect 11057 21607 11115 21613
rect 11057 21573 11069 21607
rect 11103 21604 11115 21607
rect 11164 21604 11192 21632
rect 11103 21576 11192 21604
rect 11103 21573 11115 21576
rect 11057 21567 11115 21573
rect 11238 21564 11244 21616
rect 11296 21604 11302 21616
rect 11885 21607 11943 21613
rect 11885 21604 11897 21607
rect 11296 21576 11897 21604
rect 11296 21564 11302 21576
rect 11885 21573 11897 21576
rect 11931 21573 11943 21607
rect 11885 21567 11943 21573
rect 12805 21607 12863 21613
rect 12805 21573 12817 21607
rect 12851 21604 12863 21607
rect 13078 21604 13084 21616
rect 12851 21576 13084 21604
rect 12851 21573 12863 21576
rect 12805 21567 12863 21573
rect 13078 21564 13084 21576
rect 13136 21564 13142 21616
rect 14918 21564 14924 21616
rect 14976 21604 14982 21616
rect 17310 21604 17316 21616
rect 14976 21576 17316 21604
rect 14976 21564 14982 21576
rect 17310 21564 17316 21576
rect 17368 21564 17374 21616
rect 17604 21604 17632 21644
rect 17420 21576 17632 21604
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21505 8907 21539
rect 8849 21499 8907 21505
rect 8941 21539 8999 21545
rect 8941 21505 8953 21539
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21505 11207 21539
rect 11149 21499 11207 21505
rect 5592 21440 8524 21468
rect 5592 21428 5598 21440
rect 8018 21360 8024 21412
rect 8076 21400 8082 21412
rect 8205 21403 8263 21409
rect 8205 21400 8217 21403
rect 8076 21372 8217 21400
rect 8076 21360 8082 21372
rect 8205 21369 8217 21372
rect 8251 21369 8263 21403
rect 8205 21363 8263 21369
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 3237 21335 3295 21341
rect 3237 21332 3249 21335
rect 2832 21304 3249 21332
rect 2832 21292 2838 21304
rect 3237 21301 3249 21304
rect 3283 21301 3295 21335
rect 3237 21295 3295 21301
rect 4617 21335 4675 21341
rect 4617 21301 4629 21335
rect 4663 21332 4675 21335
rect 4798 21332 4804 21344
rect 4663 21304 4804 21332
rect 4663 21301 4675 21304
rect 4617 21295 4675 21301
rect 4798 21292 4804 21304
rect 4856 21292 4862 21344
rect 6730 21292 6736 21344
rect 6788 21332 6794 21344
rect 7650 21332 7656 21344
rect 6788 21304 7656 21332
rect 6788 21292 6794 21304
rect 7650 21292 7656 21304
rect 7708 21332 7714 21344
rect 8113 21335 8171 21341
rect 8113 21332 8125 21335
rect 7708 21304 8125 21332
rect 7708 21292 7714 21304
rect 8113 21301 8125 21304
rect 8159 21301 8171 21335
rect 8864 21332 8892 21499
rect 9217 21471 9275 21477
rect 9217 21437 9229 21471
rect 9263 21468 9275 21471
rect 9766 21468 9772 21480
rect 9263 21440 9772 21468
rect 9263 21437 9275 21440
rect 9217 21431 9275 21437
rect 9766 21428 9772 21440
rect 9824 21428 9830 21480
rect 10689 21471 10747 21477
rect 10689 21437 10701 21471
rect 10735 21468 10747 21471
rect 10796 21468 10824 21499
rect 11054 21468 11060 21480
rect 10735 21440 11060 21468
rect 10735 21437 10747 21440
rect 10689 21431 10747 21437
rect 11054 21428 11060 21440
rect 11112 21428 11118 21480
rect 11164 21468 11192 21499
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 11790 21496 11796 21548
rect 11848 21496 11854 21548
rect 11974 21496 11980 21548
rect 12032 21536 12038 21548
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 12032 21508 12081 21536
rect 12032 21496 12038 21508
rect 12069 21505 12081 21508
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 14185 21539 14243 21545
rect 14185 21505 14197 21539
rect 14231 21536 14243 21539
rect 14642 21536 14648 21548
rect 14231 21508 14648 21536
rect 14231 21505 14243 21508
rect 14185 21499 14243 21505
rect 14642 21496 14648 21508
rect 14700 21496 14706 21548
rect 15562 21496 15568 21548
rect 15620 21536 15626 21548
rect 16574 21536 16580 21548
rect 15620 21508 16580 21536
rect 15620 21496 15626 21508
rect 16574 21496 16580 21508
rect 16632 21536 16638 21548
rect 17221 21539 17279 21545
rect 17221 21536 17233 21539
rect 16632 21508 17233 21536
rect 16632 21496 16638 21508
rect 17221 21505 17233 21508
rect 17267 21536 17279 21539
rect 17420 21536 17448 21576
rect 17678 21564 17684 21616
rect 17736 21604 17742 21616
rect 17862 21604 17868 21616
rect 17736 21576 17868 21604
rect 17736 21564 17742 21576
rect 17862 21564 17868 21576
rect 17920 21604 17926 21616
rect 18601 21607 18659 21613
rect 18601 21604 18613 21607
rect 17920 21576 18613 21604
rect 17920 21564 17926 21576
rect 18601 21573 18613 21576
rect 18647 21573 18659 21607
rect 18601 21567 18659 21573
rect 17267 21508 17448 21536
rect 17267 21505 17279 21508
rect 17221 21499 17279 21505
rect 18230 21496 18236 21548
rect 18288 21496 18294 21548
rect 18381 21539 18439 21545
rect 18381 21505 18393 21539
rect 18427 21536 18439 21539
rect 18427 21505 18460 21536
rect 18381 21499 18460 21505
rect 12342 21468 12348 21480
rect 11164 21440 12348 21468
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 13909 21471 13967 21477
rect 13909 21437 13921 21471
rect 13955 21468 13967 21471
rect 15194 21468 15200 21480
rect 13955 21440 15200 21468
rect 13955 21437 13967 21440
rect 13909 21431 13967 21437
rect 15194 21428 15200 21440
rect 15252 21428 15258 21480
rect 17497 21471 17555 21477
rect 17497 21437 17509 21471
rect 17543 21468 17555 21471
rect 18432 21468 18460 21499
rect 18506 21496 18512 21548
rect 18564 21496 18570 21548
rect 18708 21545 18736 21644
rect 18877 21641 18889 21675
rect 18923 21641 18935 21675
rect 18877 21635 18935 21641
rect 18892 21604 18920 21635
rect 19518 21632 19524 21684
rect 19576 21672 19582 21684
rect 20165 21675 20223 21681
rect 20165 21672 20177 21675
rect 19576 21644 20177 21672
rect 19576 21632 19582 21644
rect 20165 21641 20177 21644
rect 20211 21641 20223 21675
rect 20165 21635 20223 21641
rect 20346 21632 20352 21684
rect 20404 21632 20410 21684
rect 21634 21632 21640 21684
rect 21692 21672 21698 21684
rect 24486 21672 24492 21684
rect 21692 21644 24492 21672
rect 21692 21632 21698 21644
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 26326 21632 26332 21684
rect 26384 21672 26390 21684
rect 29914 21672 29920 21684
rect 26384 21644 29920 21672
rect 26384 21632 26390 21644
rect 29914 21632 29920 21644
rect 29972 21632 29978 21684
rect 35897 21675 35955 21681
rect 35897 21641 35909 21675
rect 35943 21672 35955 21675
rect 36446 21672 36452 21684
rect 35943 21644 36452 21672
rect 35943 21641 35955 21644
rect 35897 21635 35955 21641
rect 36446 21632 36452 21644
rect 36504 21632 36510 21684
rect 18892 21576 19845 21604
rect 18698 21539 18756 21545
rect 18698 21505 18710 21539
rect 18744 21536 18756 21539
rect 19150 21536 19156 21548
rect 18744 21508 19156 21536
rect 18744 21505 18756 21508
rect 18698 21499 18756 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 19242 21496 19248 21548
rect 19300 21536 19306 21548
rect 19429 21539 19487 21545
rect 19429 21536 19441 21539
rect 19300 21508 19441 21536
rect 19300 21496 19306 21508
rect 19429 21505 19441 21508
rect 19475 21505 19487 21539
rect 19429 21499 19487 21505
rect 19702 21496 19708 21548
rect 19760 21496 19766 21548
rect 19817 21545 19845 21576
rect 21082 21564 21088 21616
rect 21140 21604 21146 21616
rect 23829 21607 23887 21613
rect 23829 21604 23841 21607
rect 21140 21576 23841 21604
rect 21140 21564 21146 21576
rect 23829 21573 23841 21576
rect 23875 21604 23887 21607
rect 23875 21573 23888 21604
rect 23829 21567 23888 21573
rect 19797 21539 19855 21545
rect 19797 21505 19809 21539
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20346 21536 20352 21548
rect 20303 21508 20352 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 20441 21539 20499 21545
rect 20441 21505 20453 21539
rect 20487 21536 20499 21539
rect 22002 21536 22008 21548
rect 20487 21508 22008 21536
rect 20487 21505 20499 21508
rect 20441 21499 20499 21505
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 23860 21536 23888 21567
rect 24026 21564 24032 21616
rect 24084 21604 24090 21616
rect 24210 21604 24216 21616
rect 24084 21576 24216 21604
rect 24084 21564 24090 21576
rect 24210 21564 24216 21576
rect 24268 21564 24274 21616
rect 28442 21564 28448 21616
rect 28500 21604 28506 21616
rect 29089 21607 29147 21613
rect 28500 21576 28948 21604
rect 28500 21564 28506 21576
rect 25498 21536 25504 21548
rect 23860 21508 25504 21536
rect 25498 21496 25504 21508
rect 25556 21496 25562 21548
rect 28810 21496 28816 21548
rect 28868 21496 28874 21548
rect 28920 21545 28948 21576
rect 29089 21573 29101 21607
rect 29135 21604 29147 21607
rect 31202 21604 31208 21616
rect 29135 21576 31208 21604
rect 29135 21573 29147 21576
rect 29089 21567 29147 21573
rect 31202 21564 31208 21576
rect 31260 21564 31266 21616
rect 28906 21539 28964 21545
rect 28906 21505 28918 21539
rect 28952 21505 28964 21539
rect 28906 21499 28964 21505
rect 29178 21496 29184 21548
rect 29236 21496 29242 21548
rect 29278 21539 29336 21545
rect 29278 21505 29290 21539
rect 29324 21536 29336 21539
rect 29324 21508 29408 21536
rect 29324 21505 29336 21508
rect 29278 21499 29336 21505
rect 19889 21471 19947 21477
rect 17543 21440 19845 21468
rect 17543 21437 17555 21440
rect 17497 21431 17555 21437
rect 10318 21360 10324 21412
rect 10376 21400 10382 21412
rect 11698 21400 11704 21412
rect 10376 21372 11704 21400
rect 10376 21360 10382 21372
rect 11698 21360 11704 21372
rect 11756 21360 11762 21412
rect 13262 21360 13268 21412
rect 13320 21400 13326 21412
rect 14090 21400 14096 21412
rect 13320 21372 14096 21400
rect 13320 21360 13326 21372
rect 14090 21360 14096 21372
rect 14148 21360 14154 21412
rect 19245 21403 19303 21409
rect 19245 21369 19257 21403
rect 19291 21400 19303 21403
rect 19817 21400 19845 21440
rect 19889 21437 19901 21471
rect 19935 21468 19947 21471
rect 20070 21468 20076 21480
rect 19935 21440 20076 21468
rect 19935 21437 19947 21440
rect 19889 21431 19947 21437
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 20622 21428 20628 21480
rect 20680 21468 20686 21480
rect 22370 21468 22376 21480
rect 20680 21440 22376 21468
rect 20680 21428 20686 21440
rect 22370 21428 22376 21440
rect 22428 21468 22434 21480
rect 24486 21468 24492 21480
rect 22428 21440 24492 21468
rect 22428 21428 22434 21440
rect 24486 21428 24492 21440
rect 24544 21468 24550 21480
rect 25130 21468 25136 21480
rect 24544 21440 25136 21468
rect 24544 21428 24550 21440
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 19291 21372 19748 21400
rect 19817 21372 20944 21400
rect 19291 21369 19303 21372
rect 19245 21363 19303 21369
rect 11238 21332 11244 21344
rect 8864 21304 11244 21332
rect 8113 21295 8171 21301
rect 11238 21292 11244 21304
rect 11296 21292 11302 21344
rect 11330 21292 11336 21344
rect 11388 21292 11394 21344
rect 11514 21292 11520 21344
rect 11572 21292 11578 21344
rect 12526 21292 12532 21344
rect 12584 21332 12590 21344
rect 12621 21335 12679 21341
rect 12621 21332 12633 21335
rect 12584 21304 12633 21332
rect 12584 21292 12590 21304
rect 12621 21301 12633 21304
rect 12667 21301 12679 21335
rect 12621 21295 12679 21301
rect 13538 21292 13544 21344
rect 13596 21332 13602 21344
rect 13817 21335 13875 21341
rect 13817 21332 13829 21335
rect 13596 21304 13829 21332
rect 13596 21292 13602 21304
rect 13817 21301 13829 21304
rect 13863 21332 13875 21335
rect 14458 21332 14464 21344
rect 13863 21304 14464 21332
rect 13863 21301 13875 21304
rect 13817 21295 13875 21301
rect 14458 21292 14464 21304
rect 14516 21292 14522 21344
rect 17310 21292 17316 21344
rect 17368 21292 17374 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19613 21335 19671 21341
rect 19613 21332 19625 21335
rect 19392 21304 19625 21332
rect 19392 21292 19398 21304
rect 19613 21301 19625 21304
rect 19659 21301 19671 21335
rect 19720 21332 19748 21372
rect 20916 21344 20944 21372
rect 22646 21360 22652 21412
rect 22704 21400 22710 21412
rect 22704 21372 23888 21400
rect 22704 21360 22710 21372
rect 19797 21335 19855 21341
rect 19797 21332 19809 21335
rect 19720 21304 19809 21332
rect 19613 21295 19671 21301
rect 19797 21301 19809 21304
rect 19843 21301 19855 21335
rect 19797 21295 19855 21301
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 23106 21332 23112 21344
rect 20956 21304 23112 21332
rect 20956 21292 20962 21304
rect 23106 21292 23112 21304
rect 23164 21292 23170 21344
rect 23658 21292 23664 21344
rect 23716 21292 23722 21344
rect 23860 21341 23888 21372
rect 26050 21360 26056 21412
rect 26108 21400 26114 21412
rect 28534 21400 28540 21412
rect 26108 21372 28540 21400
rect 26108 21360 26114 21372
rect 28534 21360 28540 21372
rect 28592 21360 28598 21412
rect 23845 21335 23903 21341
rect 23845 21301 23857 21335
rect 23891 21332 23903 21335
rect 27706 21332 27712 21344
rect 23891 21304 27712 21332
rect 23891 21301 23903 21304
rect 23845 21295 23903 21301
rect 27706 21292 27712 21304
rect 27764 21292 27770 21344
rect 29380 21332 29408 21508
rect 29546 21496 29552 21548
rect 29604 21496 29610 21548
rect 30098 21496 30104 21548
rect 30156 21536 30162 21548
rect 32766 21536 32772 21548
rect 30156 21508 32772 21536
rect 30156 21496 30162 21508
rect 32766 21496 32772 21508
rect 32824 21496 32830 21548
rect 36078 21496 36084 21548
rect 36136 21496 36142 21548
rect 29457 21403 29515 21409
rect 29457 21369 29469 21403
rect 29503 21400 29515 21403
rect 31202 21400 31208 21412
rect 29503 21372 31208 21400
rect 29503 21369 29515 21372
rect 29457 21363 29515 21369
rect 31202 21360 31208 21372
rect 31260 21360 31266 21412
rect 29733 21335 29791 21341
rect 29733 21332 29745 21335
rect 29380 21304 29745 21332
rect 29733 21301 29745 21304
rect 29779 21332 29791 21335
rect 30742 21332 30748 21344
rect 29779 21304 30748 21332
rect 29779 21301 29791 21304
rect 29733 21295 29791 21301
rect 30742 21292 30748 21304
rect 30800 21292 30806 21344
rect 1104 21242 36432 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 36432 21242
rect 1104 21168 36432 21190
rect 2130 21088 2136 21140
rect 2188 21088 2194 21140
rect 3050 21088 3056 21140
rect 3108 21128 3114 21140
rect 6822 21128 6828 21140
rect 3108 21100 6828 21128
rect 3108 21088 3114 21100
rect 6822 21088 6828 21100
rect 6880 21088 6886 21140
rect 9766 21088 9772 21140
rect 9824 21088 9830 21140
rect 10594 21088 10600 21140
rect 10652 21128 10658 21140
rect 10778 21128 10784 21140
rect 10652 21100 10784 21128
rect 10652 21088 10658 21100
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11330 21088 11336 21140
rect 11388 21128 11394 21140
rect 11885 21131 11943 21137
rect 11388 21100 11652 21128
rect 11388 21088 11394 21100
rect 2866 21020 2872 21072
rect 2924 21060 2930 21072
rect 2924 21032 3280 21060
rect 2924 21020 2930 21032
rect 2222 20952 2228 21004
rect 2280 20992 2286 21004
rect 2593 20995 2651 21001
rect 2593 20992 2605 20995
rect 2280 20964 2605 20992
rect 2280 20952 2286 20964
rect 2593 20961 2605 20964
rect 2639 20961 2651 20995
rect 2593 20955 2651 20961
rect 2682 20952 2688 21004
rect 2740 20952 2746 21004
rect 2501 20927 2559 20933
rect 2501 20893 2513 20927
rect 2547 20924 2559 20927
rect 2774 20924 2780 20936
rect 2547 20896 2780 20924
rect 2547 20893 2559 20896
rect 2501 20887 2559 20893
rect 2774 20884 2780 20896
rect 2832 20884 2838 20936
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 3050 20924 3056 20936
rect 3007 20896 3056 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 3252 20933 3280 21032
rect 6362 21020 6368 21072
rect 6420 21060 6426 21072
rect 6914 21060 6920 21072
rect 6420 21032 6920 21060
rect 6420 21020 6426 21032
rect 6914 21020 6920 21032
rect 6972 21060 6978 21072
rect 6972 21032 7420 21060
rect 6972 21020 6978 21032
rect 4706 20992 4712 21004
rect 3344 20964 4712 20992
rect 3344 20933 3372 20964
rect 4706 20952 4712 20964
rect 4764 20952 4770 21004
rect 5258 20992 5264 21004
rect 4908 20964 5264 20992
rect 3237 20927 3295 20933
rect 3237 20893 3249 20927
rect 3283 20893 3295 20927
rect 3237 20887 3295 20893
rect 3329 20927 3387 20933
rect 3329 20893 3341 20927
rect 3375 20893 3387 20927
rect 3329 20887 3387 20893
rect 4614 20884 4620 20936
rect 4672 20884 4678 20936
rect 4908 20933 4936 20964
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5350 20952 5356 21004
rect 5408 20992 5414 21004
rect 7392 21001 7420 21032
rect 7466 21020 7472 21072
rect 7524 21020 7530 21072
rect 7650 21020 7656 21072
rect 7708 21060 7714 21072
rect 9030 21060 9036 21072
rect 7708 21032 9036 21060
rect 7708 21020 7714 21032
rect 9030 21020 9036 21032
rect 9088 21020 9094 21072
rect 11054 21020 11060 21072
rect 11112 21060 11118 21072
rect 11112 21032 11192 21060
rect 11112 21020 11118 21032
rect 7377 20995 7435 21001
rect 5408 20964 7144 20992
rect 5408 20952 5414 20964
rect 4893 20927 4951 20933
rect 4893 20893 4905 20927
rect 4939 20893 4951 20927
rect 4893 20887 4951 20893
rect 4982 20884 4988 20936
rect 5040 20884 5046 20936
rect 6730 20884 6736 20936
rect 6788 20884 6794 20936
rect 7006 20884 7012 20936
rect 7064 20884 7070 20936
rect 7116 20933 7144 20964
rect 7377 20961 7389 20995
rect 7423 20961 7435 20995
rect 7377 20955 7435 20961
rect 7484 20964 7972 20992
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7484 20924 7512 20964
rect 7147 20896 7512 20924
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7650 20884 7656 20936
rect 7708 20884 7714 20936
rect 7744 20927 7802 20933
rect 7744 20893 7756 20927
rect 7790 20924 7802 20927
rect 7834 20924 7840 20936
rect 7790 20896 7840 20924
rect 7790 20893 7802 20896
rect 7744 20887 7802 20893
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 7944 20924 7972 20964
rect 8386 20952 8392 21004
rect 8444 20992 8450 21004
rect 8757 20995 8815 21001
rect 8757 20992 8769 20995
rect 8444 20964 8769 20992
rect 8444 20952 8450 20964
rect 8757 20961 8769 20964
rect 8803 20992 8815 20995
rect 8938 20992 8944 21004
rect 8803 20964 8944 20992
rect 8803 20961 8815 20964
rect 8757 20955 8815 20961
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 9398 20952 9404 21004
rect 9456 20952 9462 21004
rect 9493 20995 9551 21001
rect 9493 20961 9505 20995
rect 9539 20992 9551 20995
rect 10413 20995 10471 21001
rect 10413 20992 10425 20995
rect 9539 20964 10425 20992
rect 9539 20961 9551 20964
rect 9493 20955 9551 20961
rect 7944 20896 8800 20924
rect 3145 20859 3203 20865
rect 3145 20825 3157 20859
rect 3191 20856 3203 20859
rect 4801 20859 4859 20865
rect 4801 20856 4813 20859
rect 3191 20828 4813 20856
rect 3191 20825 3203 20828
rect 3145 20819 3203 20825
rect 3252 20800 3280 20828
rect 4801 20825 4813 20828
rect 4847 20825 4859 20859
rect 5000 20856 5028 20884
rect 8772 20868 8800 20896
rect 6917 20859 6975 20865
rect 6917 20856 6929 20859
rect 5000 20828 6929 20856
rect 4801 20819 4859 20825
rect 6917 20825 6929 20828
rect 6963 20856 6975 20859
rect 8570 20856 8576 20868
rect 6963 20828 8576 20856
rect 6963 20825 6975 20828
rect 6917 20819 6975 20825
rect 8570 20816 8576 20828
rect 8628 20816 8634 20868
rect 8754 20816 8760 20868
rect 8812 20816 8818 20868
rect 9309 20859 9367 20865
rect 9309 20825 9321 20859
rect 9355 20856 9367 20859
rect 9398 20856 9404 20868
rect 9355 20828 9404 20856
rect 9355 20825 9367 20828
rect 9309 20819 9367 20825
rect 9398 20816 9404 20828
rect 9456 20816 9462 20868
rect 3234 20748 3240 20800
rect 3292 20748 3298 20800
rect 3513 20791 3571 20797
rect 3513 20757 3525 20791
rect 3559 20788 3571 20791
rect 4522 20788 4528 20800
rect 3559 20760 4528 20788
rect 3559 20757 3571 20760
rect 3513 20751 3571 20757
rect 4522 20748 4528 20760
rect 4580 20748 4586 20800
rect 5169 20791 5227 20797
rect 5169 20757 5181 20791
rect 5215 20788 5227 20791
rect 5258 20788 5264 20800
rect 5215 20760 5264 20788
rect 5215 20757 5227 20760
rect 5169 20751 5227 20757
rect 5258 20748 5264 20760
rect 5316 20748 5322 20800
rect 7285 20791 7343 20797
rect 7285 20757 7297 20791
rect 7331 20788 7343 20791
rect 7558 20788 7564 20800
rect 7331 20760 7564 20788
rect 7331 20757 7343 20760
rect 7285 20751 7343 20757
rect 7558 20748 7564 20760
rect 7616 20748 7622 20800
rect 7742 20748 7748 20800
rect 7800 20788 7806 20800
rect 7929 20791 7987 20797
rect 7929 20788 7941 20791
rect 7800 20760 7941 20788
rect 7800 20748 7806 20760
rect 7929 20757 7941 20760
rect 7975 20757 7987 20791
rect 7929 20751 7987 20757
rect 8110 20748 8116 20800
rect 8168 20748 8174 20800
rect 8938 20748 8944 20800
rect 8996 20748 9002 20800
rect 9122 20748 9128 20800
rect 9180 20788 9186 20800
rect 9692 20788 9720 20964
rect 10413 20961 10425 20964
rect 10459 20992 10471 20995
rect 10502 20992 10508 21004
rect 10459 20964 10508 20992
rect 10459 20961 10471 20964
rect 10413 20955 10471 20961
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 11164 21001 11192 21032
rect 11514 21020 11520 21072
rect 11572 21020 11578 21072
rect 11624 21069 11652 21100
rect 11885 21097 11897 21131
rect 11931 21128 11943 21131
rect 12066 21128 12072 21140
rect 11931 21100 12072 21128
rect 11931 21097 11943 21100
rect 11885 21091 11943 21097
rect 12066 21088 12072 21100
rect 12124 21088 12130 21140
rect 12161 21131 12219 21137
rect 12161 21097 12173 21131
rect 12207 21128 12219 21131
rect 12250 21128 12256 21140
rect 12207 21100 12256 21128
rect 12207 21097 12219 21100
rect 12161 21091 12219 21097
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 14093 21131 14151 21137
rect 14093 21128 14105 21131
rect 12360 21100 14105 21128
rect 11609 21063 11667 21069
rect 11609 21029 11621 21063
rect 11655 21029 11667 21063
rect 12360 21060 12388 21100
rect 14093 21097 14105 21100
rect 14139 21097 14151 21131
rect 14093 21091 14151 21097
rect 11609 21023 11667 21029
rect 11900 21032 12388 21060
rect 12437 21063 12495 21069
rect 11149 20995 11207 21001
rect 11149 20961 11161 20995
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 10226 20884 10232 20936
rect 10284 20924 10290 20936
rect 10284 20896 10824 20924
rect 10284 20884 10290 20896
rect 10796 20868 10824 20896
rect 11054 20884 11060 20936
rect 11112 20924 11118 20936
rect 11425 20927 11483 20933
rect 11425 20924 11437 20927
rect 11112 20896 11437 20924
rect 11112 20884 11118 20896
rect 11425 20893 11437 20896
rect 11471 20893 11483 20927
rect 11425 20887 11483 20893
rect 11698 20884 11704 20936
rect 11756 20884 11762 20936
rect 10137 20859 10195 20865
rect 10137 20825 10149 20859
rect 10183 20856 10195 20859
rect 10597 20859 10655 20865
rect 10597 20856 10609 20859
rect 10183 20828 10609 20856
rect 10183 20825 10195 20828
rect 10137 20819 10195 20825
rect 10597 20825 10609 20828
rect 10643 20825 10655 20859
rect 10597 20819 10655 20825
rect 10778 20816 10784 20868
rect 10836 20816 10842 20868
rect 9180 20760 9720 20788
rect 11900 20788 11928 21032
rect 12437 21029 12449 21063
rect 12483 21060 12495 21063
rect 12483 21032 12572 21060
rect 12483 21029 12495 21032
rect 12437 21023 12495 21029
rect 12250 20952 12256 21004
rect 12308 20992 12314 21004
rect 12544 20992 12572 21032
rect 12618 21020 12624 21072
rect 12676 21060 12682 21072
rect 13354 21060 13360 21072
rect 12676 21032 13360 21060
rect 12676 21020 12682 21032
rect 13354 21020 13360 21032
rect 13412 21020 13418 21072
rect 13446 21020 13452 21072
rect 13504 21060 13510 21072
rect 13504 21032 13676 21060
rect 13504 21020 13510 21032
rect 12308 20964 12572 20992
rect 12308 20952 12314 20964
rect 12618 20884 12624 20936
rect 12676 20884 12682 20936
rect 12710 20884 12716 20936
rect 12768 20884 12774 20936
rect 13173 20927 13231 20933
rect 13173 20924 13185 20927
rect 12912 20896 13185 20924
rect 11977 20859 12035 20865
rect 11977 20825 11989 20859
rect 12023 20856 12035 20859
rect 12526 20856 12532 20868
rect 12023 20828 12532 20856
rect 12023 20825 12035 20828
rect 11977 20819 12035 20825
rect 12526 20816 12532 20828
rect 12584 20856 12590 20868
rect 12802 20856 12808 20868
rect 12584 20828 12808 20856
rect 12584 20816 12590 20828
rect 12802 20816 12808 20828
rect 12860 20816 12866 20868
rect 12177 20791 12235 20797
rect 12177 20788 12189 20791
rect 11900 20760 12189 20788
rect 9180 20748 9186 20760
rect 12177 20757 12189 20760
rect 12223 20757 12235 20791
rect 12177 20751 12235 20757
rect 12345 20791 12403 20797
rect 12345 20757 12357 20791
rect 12391 20788 12403 20791
rect 12912 20788 12940 20896
rect 13173 20893 13185 20896
rect 13219 20893 13231 20927
rect 13173 20887 13231 20893
rect 13262 20884 13268 20936
rect 13320 20924 13326 20936
rect 13449 20927 13507 20933
rect 13449 20924 13461 20927
rect 13320 20896 13461 20924
rect 13320 20884 13326 20896
rect 13449 20893 13461 20896
rect 13495 20893 13507 20927
rect 13449 20887 13507 20893
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 12989 20859 13047 20865
rect 12989 20825 13001 20859
rect 13035 20825 13047 20859
rect 12989 20819 13047 20825
rect 12391 20760 12940 20788
rect 13004 20788 13032 20819
rect 13078 20816 13084 20868
rect 13136 20816 13142 20868
rect 13354 20816 13360 20868
rect 13412 20816 13418 20868
rect 13170 20788 13176 20800
rect 13004 20760 13176 20788
rect 12391 20757 12403 20760
rect 12345 20751 12403 20757
rect 13170 20748 13176 20760
rect 13228 20788 13234 20800
rect 13556 20788 13584 20887
rect 13648 20856 13676 21032
rect 14108 20992 14136 21091
rect 17126 21088 17132 21140
rect 17184 21128 17190 21140
rect 17221 21131 17279 21137
rect 17221 21128 17233 21131
rect 17184 21100 17233 21128
rect 17184 21088 17190 21100
rect 17221 21097 17233 21100
rect 17267 21097 17279 21131
rect 17221 21091 17279 21097
rect 17310 21088 17316 21140
rect 17368 21128 17374 21140
rect 18506 21128 18512 21140
rect 17368 21100 18512 21128
rect 17368 21088 17374 21100
rect 18506 21088 18512 21100
rect 18564 21088 18570 21140
rect 19150 21088 19156 21140
rect 19208 21128 19214 21140
rect 19702 21128 19708 21140
rect 19208 21100 19708 21128
rect 19208 21088 19214 21100
rect 19702 21088 19708 21100
rect 19760 21128 19766 21140
rect 20622 21128 20628 21140
rect 19760 21100 20628 21128
rect 19760 21088 19766 21100
rect 20622 21088 20628 21100
rect 20680 21088 20686 21140
rect 21637 21131 21695 21137
rect 21637 21097 21649 21131
rect 21683 21128 21695 21131
rect 21910 21128 21916 21140
rect 21683 21100 21916 21128
rect 21683 21097 21695 21100
rect 21637 21091 21695 21097
rect 21910 21088 21916 21100
rect 21968 21088 21974 21140
rect 22922 21088 22928 21140
rect 22980 21088 22986 21140
rect 23566 21088 23572 21140
rect 23624 21088 23630 21140
rect 23934 21088 23940 21140
rect 23992 21088 23998 21140
rect 25041 21131 25099 21137
rect 25041 21128 25053 21131
rect 24044 21100 25053 21128
rect 16390 21060 16396 21072
rect 15212 21032 16396 21060
rect 15105 20995 15163 21001
rect 15105 20992 15117 20995
rect 14108 20964 15117 20992
rect 15105 20961 15117 20964
rect 15151 20961 15163 20995
rect 15105 20955 15163 20961
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20924 14151 20927
rect 14182 20924 14188 20936
rect 14139 20896 14188 20924
rect 14139 20893 14151 20896
rect 14093 20887 14151 20893
rect 14182 20884 14188 20896
rect 14240 20884 14246 20936
rect 14274 20884 14280 20936
rect 14332 20884 14338 20936
rect 15212 20933 15240 21032
rect 16390 21020 16396 21032
rect 16448 21020 16454 21072
rect 19886 21020 19892 21072
rect 19944 21060 19950 21072
rect 22649 21063 22707 21069
rect 22649 21060 22661 21063
rect 19944 21032 22661 21060
rect 19944 21020 19950 21032
rect 22649 21029 22661 21032
rect 22695 21029 22707 21063
rect 22649 21023 22707 21029
rect 23753 21063 23811 21069
rect 23753 21029 23765 21063
rect 23799 21029 23811 21063
rect 24044 21060 24072 21100
rect 25041 21097 25053 21100
rect 25087 21097 25099 21131
rect 25041 21091 25099 21097
rect 26326 21088 26332 21140
rect 26384 21128 26390 21140
rect 26881 21131 26939 21137
rect 26881 21128 26893 21131
rect 26384 21100 26893 21128
rect 26384 21088 26390 21100
rect 26881 21097 26893 21100
rect 26927 21128 26939 21131
rect 26970 21128 26976 21140
rect 26927 21100 26976 21128
rect 26927 21097 26939 21100
rect 26881 21091 26939 21097
rect 26970 21088 26976 21100
rect 27028 21088 27034 21140
rect 28994 21088 29000 21140
rect 29052 21128 29058 21140
rect 29546 21128 29552 21140
rect 29052 21100 29552 21128
rect 29052 21088 29058 21100
rect 29546 21088 29552 21100
rect 29604 21088 29610 21140
rect 32766 21088 32772 21140
rect 32824 21088 32830 21140
rect 23753 21023 23811 21029
rect 23952 21032 24072 21060
rect 15378 20952 15384 21004
rect 15436 20952 15442 21004
rect 19518 20952 19524 21004
rect 19576 20992 19582 21004
rect 19978 20992 19984 21004
rect 19576 20964 19984 20992
rect 19576 20952 19582 20964
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 23017 20995 23075 21001
rect 23017 20961 23029 20995
rect 23063 20992 23075 20995
rect 23768 20992 23796 21023
rect 23063 20964 23796 20992
rect 23063 20961 23075 20964
rect 23017 20955 23075 20961
rect 15197 20927 15255 20933
rect 15197 20893 15209 20927
rect 15243 20893 15255 20927
rect 15197 20887 15255 20893
rect 15289 20927 15347 20933
rect 15289 20893 15301 20927
rect 15335 20924 15347 20927
rect 15654 20924 15660 20936
rect 15335 20896 15660 20924
rect 15335 20893 15347 20896
rect 15289 20887 15347 20893
rect 13648 20828 14228 20856
rect 13228 20760 13584 20788
rect 13725 20791 13783 20797
rect 13228 20748 13234 20760
rect 13725 20757 13737 20791
rect 13771 20788 13783 20791
rect 14090 20788 14096 20800
rect 13771 20760 14096 20788
rect 13771 20757 13783 20760
rect 13725 20751 13783 20757
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 14200 20788 14228 20828
rect 15304 20788 15332 20887
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 15930 20884 15936 20936
rect 15988 20924 15994 20936
rect 16301 20927 16359 20933
rect 16301 20924 16313 20927
rect 15988 20896 16313 20924
rect 15988 20884 15994 20896
rect 16301 20893 16313 20896
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20924 17003 20927
rect 17034 20924 17040 20936
rect 16991 20896 17040 20924
rect 16991 20893 17003 20896
rect 16945 20887 17003 20893
rect 17034 20884 17040 20896
rect 17092 20884 17098 20936
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 18012 20896 19748 20924
rect 18012 20884 18018 20896
rect 16390 20816 16396 20868
rect 16448 20856 16454 20868
rect 18230 20856 18236 20868
rect 16448 20828 18236 20856
rect 16448 20816 16454 20828
rect 18230 20816 18236 20828
rect 18288 20816 18294 20868
rect 19337 20859 19395 20865
rect 19337 20825 19349 20859
rect 19383 20856 19395 20859
rect 19610 20856 19616 20868
rect 19383 20828 19616 20856
rect 19383 20825 19395 20828
rect 19337 20819 19395 20825
rect 19610 20816 19616 20828
rect 19668 20816 19674 20868
rect 14200 20760 15332 20788
rect 15565 20791 15623 20797
rect 15565 20757 15577 20791
rect 15611 20788 15623 20791
rect 15654 20788 15660 20800
rect 15611 20760 15660 20788
rect 15611 20757 15623 20760
rect 15565 20751 15623 20757
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 15746 20748 15752 20800
rect 15804 20748 15810 20800
rect 17862 20748 17868 20800
rect 17920 20788 17926 20800
rect 19429 20791 19487 20797
rect 19429 20788 19441 20791
rect 17920 20760 19441 20788
rect 17920 20748 17926 20760
rect 19429 20757 19441 20760
rect 19475 20757 19487 20791
rect 19720 20788 19748 20896
rect 19996 20856 20024 20952
rect 21358 20884 21364 20936
rect 21416 20884 21422 20936
rect 21450 20884 21456 20936
rect 21508 20884 21514 20936
rect 21542 20884 21548 20936
rect 21600 20884 21606 20936
rect 22833 20927 22891 20933
rect 22833 20924 22845 20927
rect 22296 20896 22845 20924
rect 21082 20856 21088 20868
rect 19996 20828 21088 20856
rect 21082 20816 21088 20828
rect 21140 20856 21146 20868
rect 21177 20859 21235 20865
rect 21177 20856 21189 20859
rect 21140 20828 21189 20856
rect 21140 20816 21146 20828
rect 21177 20825 21189 20828
rect 21223 20825 21235 20859
rect 21177 20819 21235 20825
rect 22186 20816 22192 20868
rect 22244 20816 22250 20868
rect 22296 20800 22324 20896
rect 22833 20893 22845 20896
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 23032 20896 23336 20924
rect 22373 20859 22431 20865
rect 22373 20825 22385 20859
rect 22419 20856 22431 20859
rect 23032 20856 23060 20896
rect 22419 20828 23060 20856
rect 22419 20825 22431 20828
rect 22373 20819 22431 20825
rect 23106 20816 23112 20868
rect 23164 20816 23170 20868
rect 22094 20788 22100 20800
rect 19720 20760 22100 20788
rect 19429 20751 19487 20757
rect 22094 20748 22100 20760
rect 22152 20748 22158 20800
rect 22278 20748 22284 20800
rect 22336 20788 22342 20800
rect 22557 20791 22615 20797
rect 22557 20788 22569 20791
rect 22336 20760 22569 20788
rect 22336 20748 22342 20760
rect 22557 20757 22569 20760
rect 22603 20757 22615 20791
rect 22557 20751 22615 20757
rect 22830 20748 22836 20800
rect 22888 20788 22894 20800
rect 23201 20791 23259 20797
rect 23201 20788 23213 20791
rect 22888 20760 23213 20788
rect 22888 20748 22894 20760
rect 23201 20757 23213 20760
rect 23247 20757 23259 20791
rect 23308 20788 23336 20896
rect 23382 20884 23388 20936
rect 23440 20884 23446 20936
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20893 23535 20927
rect 23477 20887 23535 20893
rect 23492 20856 23520 20887
rect 23658 20884 23664 20936
rect 23716 20884 23722 20936
rect 23952 20933 23980 21032
rect 24486 21020 24492 21072
rect 24544 21020 24550 21072
rect 24578 21020 24584 21072
rect 24636 21060 24642 21072
rect 29362 21060 29368 21072
rect 24636 21032 24900 21060
rect 24636 21020 24642 21032
rect 24504 20992 24532 21020
rect 24504 20964 24716 20992
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20893 23995 20927
rect 23937 20887 23995 20893
rect 24026 20884 24032 20936
rect 24084 20884 24090 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 24136 20896 24409 20924
rect 24044 20856 24072 20884
rect 23492 20828 24072 20856
rect 23474 20788 23480 20800
rect 23308 20760 23480 20788
rect 23201 20751 23259 20757
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 23658 20748 23664 20800
rect 23716 20788 23722 20800
rect 24136 20788 24164 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 24486 20884 24492 20936
rect 24544 20884 24550 20936
rect 24688 20933 24716 20964
rect 24673 20927 24731 20933
rect 24673 20893 24685 20927
rect 24719 20893 24731 20927
rect 24673 20887 24731 20893
rect 24762 20884 24768 20936
rect 24820 20884 24826 20936
rect 24872 20924 24900 21032
rect 26712 21032 29368 21060
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25004 20964 26280 20992
rect 25004 20952 25010 20964
rect 25225 20927 25283 20933
rect 25225 20924 25237 20927
rect 24872 20896 25237 20924
rect 25225 20893 25237 20896
rect 25271 20893 25283 20927
rect 25225 20887 25283 20893
rect 25498 20884 25504 20936
rect 25556 20884 25562 20936
rect 26252 20933 26280 20964
rect 26237 20927 26295 20933
rect 26237 20893 26249 20927
rect 26283 20893 26295 20927
rect 26237 20887 26295 20893
rect 24213 20859 24271 20865
rect 24213 20825 24225 20859
rect 24259 20856 24271 20859
rect 24949 20859 25007 20865
rect 24949 20856 24961 20859
rect 24259 20828 24961 20856
rect 24259 20825 24271 20828
rect 24213 20819 24271 20825
rect 24949 20825 24961 20828
rect 24995 20825 25007 20859
rect 24949 20819 25007 20825
rect 25314 20816 25320 20868
rect 25372 20856 25378 20868
rect 25409 20859 25467 20865
rect 25409 20856 25421 20859
rect 25372 20828 25421 20856
rect 25372 20816 25378 20828
rect 25409 20825 25421 20828
rect 25455 20856 25467 20859
rect 26050 20856 26056 20868
rect 25455 20828 26056 20856
rect 25455 20825 25467 20828
rect 25409 20819 25467 20825
rect 26050 20816 26056 20828
rect 26108 20816 26114 20868
rect 26712 20865 26740 21032
rect 29362 21020 29368 21032
rect 29420 21020 29426 21072
rect 31662 21020 31668 21072
rect 31720 21060 31726 21072
rect 33134 21060 33140 21072
rect 31720 21032 33140 21060
rect 31720 21020 31726 21032
rect 33134 21020 33140 21032
rect 33192 21020 33198 21072
rect 27246 20952 27252 21004
rect 27304 20992 27310 21004
rect 27304 20964 28488 20992
rect 27304 20952 27310 20964
rect 27982 20884 27988 20936
rect 28040 20884 28046 20936
rect 28350 20884 28356 20936
rect 28408 20884 28414 20936
rect 28460 20933 28488 20964
rect 31202 20952 31208 21004
rect 31260 20992 31266 21004
rect 32861 20995 32919 21001
rect 32861 20992 32873 20995
rect 31260 20964 32873 20992
rect 31260 20952 31266 20964
rect 32861 20961 32873 20964
rect 32907 20961 32919 20995
rect 32861 20955 32919 20961
rect 28445 20927 28503 20933
rect 28445 20893 28457 20927
rect 28491 20893 28503 20927
rect 28445 20887 28503 20893
rect 31478 20884 31484 20936
rect 31536 20884 31542 20936
rect 31662 20884 31668 20936
rect 31720 20884 31726 20936
rect 31757 20927 31815 20933
rect 31757 20893 31769 20927
rect 31803 20924 31815 20927
rect 31938 20924 31944 20936
rect 31803 20896 31944 20924
rect 31803 20893 31815 20896
rect 31757 20887 31815 20893
rect 31938 20884 31944 20896
rect 31996 20884 32002 20936
rect 33042 20884 33048 20936
rect 33100 20884 33106 20936
rect 26697 20859 26755 20865
rect 26697 20825 26709 20859
rect 26743 20825 26755 20859
rect 26697 20819 26755 20825
rect 26913 20859 26971 20865
rect 26913 20825 26925 20859
rect 26959 20856 26971 20859
rect 27246 20856 27252 20868
rect 26959 20828 27252 20856
rect 26959 20825 26971 20828
rect 26913 20819 26971 20825
rect 27246 20816 27252 20828
rect 27304 20816 27310 20868
rect 28166 20865 28172 20868
rect 28143 20859 28172 20865
rect 28143 20825 28155 20859
rect 28143 20819 28172 20825
rect 28166 20816 28172 20819
rect 28224 20816 28230 20868
rect 28258 20816 28264 20868
rect 28316 20816 28322 20868
rect 32030 20816 32036 20868
rect 32088 20856 32094 20868
rect 32769 20859 32827 20865
rect 32769 20856 32781 20859
rect 32088 20828 32781 20856
rect 32088 20816 32094 20828
rect 32769 20825 32781 20828
rect 32815 20825 32827 20859
rect 32769 20819 32827 20825
rect 23716 20760 24164 20788
rect 23716 20748 23722 20760
rect 25774 20748 25780 20800
rect 25832 20788 25838 20800
rect 26329 20791 26387 20797
rect 26329 20788 26341 20791
rect 25832 20760 26341 20788
rect 25832 20748 25838 20760
rect 26329 20757 26341 20760
rect 26375 20757 26387 20791
rect 26329 20751 26387 20757
rect 26786 20748 26792 20800
rect 26844 20788 26850 20800
rect 27065 20791 27123 20797
rect 27065 20788 27077 20791
rect 26844 20760 27077 20788
rect 26844 20748 26850 20760
rect 27065 20757 27077 20760
rect 27111 20757 27123 20791
rect 27065 20751 27123 20757
rect 27706 20748 27712 20800
rect 27764 20788 27770 20800
rect 28350 20788 28356 20800
rect 27764 20760 28356 20788
rect 27764 20748 27770 20760
rect 28350 20748 28356 20760
rect 28408 20748 28414 20800
rect 28629 20791 28687 20797
rect 28629 20757 28641 20791
rect 28675 20788 28687 20791
rect 30282 20788 30288 20800
rect 28675 20760 30288 20788
rect 28675 20757 28687 20760
rect 28629 20751 28687 20757
rect 30282 20748 30288 20760
rect 30340 20748 30346 20800
rect 31294 20748 31300 20800
rect 31352 20748 31358 20800
rect 33229 20791 33287 20797
rect 33229 20757 33241 20791
rect 33275 20788 33287 20791
rect 34606 20788 34612 20800
rect 33275 20760 34612 20788
rect 33275 20757 33287 20760
rect 33229 20751 33287 20757
rect 34606 20748 34612 20760
rect 34664 20748 34670 20800
rect 1104 20698 36432 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 36432 20698
rect 1104 20624 36432 20646
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 7098 20584 7104 20596
rect 3016 20556 7104 20584
rect 3016 20544 3022 20556
rect 7098 20544 7104 20556
rect 7156 20584 7162 20596
rect 7466 20584 7472 20596
rect 7156 20556 7472 20584
rect 7156 20544 7162 20556
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 7745 20587 7803 20593
rect 7745 20553 7757 20587
rect 7791 20584 7803 20587
rect 8110 20584 8116 20596
rect 7791 20556 8116 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 8110 20544 8116 20556
rect 8168 20544 8174 20596
rect 9398 20544 9404 20596
rect 9456 20584 9462 20596
rect 10229 20587 10287 20593
rect 10229 20584 10241 20587
rect 9456 20556 10241 20584
rect 9456 20544 9462 20556
rect 10229 20553 10241 20556
rect 10275 20553 10287 20587
rect 10229 20547 10287 20553
rect 11701 20587 11759 20593
rect 11701 20553 11713 20587
rect 11747 20584 11759 20587
rect 12066 20584 12072 20596
rect 11747 20556 12072 20584
rect 11747 20553 11759 20556
rect 11701 20547 11759 20553
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 13078 20544 13084 20596
rect 13136 20544 13142 20596
rect 13354 20544 13360 20596
rect 13412 20584 13418 20596
rect 13412 20556 14964 20584
rect 13412 20544 13418 20556
rect 7282 20516 7288 20528
rect 6932 20488 7288 20516
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20417 4491 20451
rect 4433 20411 4491 20417
rect 4448 20380 4476 20411
rect 4522 20408 4528 20460
rect 4580 20408 4586 20460
rect 4890 20408 4896 20460
rect 4948 20408 4954 20460
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20448 5595 20451
rect 5810 20448 5816 20460
rect 5583 20420 5816 20448
rect 5583 20417 5595 20420
rect 5537 20411 5595 20417
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 6932 20457 6960 20488
rect 7282 20476 7288 20488
rect 7340 20476 7346 20528
rect 7837 20519 7895 20525
rect 7837 20485 7849 20519
rect 7883 20516 7895 20519
rect 8018 20516 8024 20528
rect 7883 20488 8024 20516
rect 7883 20485 7895 20488
rect 7837 20479 7895 20485
rect 8018 20476 8024 20488
rect 8076 20476 8082 20528
rect 8665 20519 8723 20525
rect 8665 20485 8677 20519
rect 8711 20516 8723 20519
rect 8938 20516 8944 20528
rect 8711 20488 8944 20516
rect 8711 20485 8723 20488
rect 8665 20479 8723 20485
rect 8938 20476 8944 20488
rect 8996 20476 9002 20528
rect 9674 20476 9680 20528
rect 9732 20476 9738 20528
rect 11422 20476 11428 20528
rect 11480 20516 11486 20528
rect 11885 20519 11943 20525
rect 11885 20516 11897 20519
rect 11480 20488 11897 20516
rect 11480 20476 11486 20488
rect 11885 20485 11897 20488
rect 11931 20485 11943 20519
rect 11885 20479 11943 20485
rect 14274 20476 14280 20528
rect 14332 20476 14338 20528
rect 14936 20516 14964 20556
rect 15010 20544 15016 20596
rect 15068 20584 15074 20596
rect 21266 20584 21272 20596
rect 15068 20556 21272 20584
rect 15068 20544 15074 20556
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 22186 20544 22192 20596
rect 22244 20584 22250 20596
rect 22281 20587 22339 20593
rect 22281 20584 22293 20587
rect 22244 20556 22293 20584
rect 22244 20544 22250 20556
rect 22281 20553 22293 20556
rect 22327 20553 22339 20587
rect 22281 20547 22339 20553
rect 24213 20587 24271 20593
rect 24213 20553 24225 20587
rect 24259 20584 24271 20587
rect 24762 20584 24768 20596
rect 24259 20556 24768 20584
rect 24259 20553 24271 20556
rect 24213 20547 24271 20553
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 24946 20544 24952 20596
rect 25004 20544 25010 20596
rect 25130 20544 25136 20596
rect 25188 20584 25194 20596
rect 25774 20584 25780 20596
rect 25188 20556 25780 20584
rect 25188 20544 25194 20556
rect 25774 20544 25780 20556
rect 25832 20544 25838 20596
rect 28166 20584 28172 20596
rect 26620 20556 28172 20584
rect 15473 20519 15531 20525
rect 14936 20488 15148 20516
rect 6917 20451 6975 20457
rect 6917 20417 6929 20451
rect 6963 20417 6975 20451
rect 6917 20411 6975 20417
rect 7006 20408 7012 20460
rect 7064 20408 7070 20460
rect 8202 20408 8208 20460
rect 8260 20448 8266 20460
rect 8389 20451 8447 20457
rect 8389 20448 8401 20451
rect 8260 20420 8401 20448
rect 8260 20408 8266 20420
rect 8389 20417 8401 20420
rect 8435 20417 8447 20451
rect 10686 20448 10692 20460
rect 8389 20411 8447 20417
rect 10152 20420 10692 20448
rect 4614 20380 4620 20392
rect 4448 20352 4620 20380
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 5626 20340 5632 20392
rect 5684 20340 5690 20392
rect 7282 20340 7288 20392
rect 7340 20380 7346 20392
rect 7650 20380 7656 20392
rect 7340 20352 7656 20380
rect 7340 20340 7346 20352
rect 7650 20340 7656 20352
rect 7708 20340 7714 20392
rect 7926 20340 7932 20392
rect 7984 20380 7990 20392
rect 8021 20383 8079 20389
rect 8021 20380 8033 20383
rect 7984 20352 8033 20380
rect 7984 20340 7990 20352
rect 8021 20349 8033 20352
rect 8067 20380 8079 20383
rect 8110 20380 8116 20392
rect 8067 20352 8116 20380
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 6914 20272 6920 20324
rect 6972 20312 6978 20324
rect 8220 20312 8248 20408
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 10152 20389 10180 20420
rect 10686 20408 10692 20420
rect 10744 20448 10750 20460
rect 10781 20451 10839 20457
rect 10781 20448 10793 20451
rect 10744 20420 10793 20448
rect 10744 20408 10750 20420
rect 10781 20417 10793 20420
rect 10827 20417 10839 20451
rect 15120 20448 15148 20488
rect 15473 20485 15485 20519
rect 15519 20516 15531 20519
rect 15746 20516 15752 20528
rect 15519 20488 15752 20516
rect 15519 20485 15531 20488
rect 15473 20479 15531 20485
rect 15746 20476 15752 20488
rect 15804 20476 15810 20528
rect 15930 20476 15936 20528
rect 15988 20476 15994 20528
rect 16114 20476 16120 20528
rect 16172 20525 16178 20528
rect 16172 20519 16191 20525
rect 16179 20485 16191 20519
rect 16172 20479 16191 20485
rect 16172 20476 16178 20479
rect 16482 20476 16488 20528
rect 16540 20516 16546 20528
rect 17497 20519 17555 20525
rect 16540 20488 16804 20516
rect 16540 20476 16546 20488
rect 15565 20451 15623 20457
rect 15565 20448 15577 20451
rect 15120 20420 15577 20448
rect 10781 20411 10839 20417
rect 15565 20417 15577 20420
rect 15611 20417 15623 20451
rect 15565 20411 15623 20417
rect 16666 20408 16672 20460
rect 16724 20408 16730 20460
rect 16776 20448 16804 20488
rect 17497 20485 17509 20519
rect 17543 20516 17555 20519
rect 17586 20516 17592 20528
rect 17543 20488 17592 20516
rect 17543 20485 17555 20488
rect 17497 20479 17555 20485
rect 17586 20476 17592 20488
rect 17644 20476 17650 20528
rect 17681 20519 17739 20525
rect 17681 20485 17693 20519
rect 17727 20485 17739 20519
rect 19981 20519 20039 20525
rect 19981 20516 19993 20519
rect 17681 20479 17739 20485
rect 19306 20488 19993 20516
rect 17696 20448 17724 20479
rect 16776 20420 17724 20448
rect 18414 20408 18420 20460
rect 18472 20448 18478 20460
rect 19306 20448 19334 20488
rect 19981 20485 19993 20488
rect 20027 20485 20039 20519
rect 19981 20479 20039 20485
rect 20346 20476 20352 20528
rect 20404 20476 20410 20528
rect 20898 20476 20904 20528
rect 20956 20476 20962 20528
rect 21117 20519 21175 20525
rect 21117 20485 21129 20519
rect 21163 20516 21175 20519
rect 21358 20516 21364 20528
rect 21163 20488 21364 20516
rect 21163 20485 21175 20488
rect 21117 20479 21175 20485
rect 21358 20476 21364 20488
rect 21416 20476 21422 20528
rect 21542 20476 21548 20528
rect 21600 20516 21606 20528
rect 21821 20519 21879 20525
rect 21821 20516 21833 20519
rect 21600 20488 21833 20516
rect 21600 20476 21606 20488
rect 21821 20485 21833 20488
rect 21867 20485 21879 20519
rect 23382 20516 23388 20528
rect 21821 20479 21879 20485
rect 22388 20488 23388 20516
rect 22388 20460 22416 20488
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 23845 20519 23903 20525
rect 23845 20485 23857 20519
rect 23891 20516 23903 20519
rect 24118 20516 24124 20528
rect 23891 20488 24124 20516
rect 23891 20485 23903 20488
rect 23845 20479 23903 20485
rect 24118 20476 24124 20488
rect 24176 20476 24182 20528
rect 25516 20488 26004 20516
rect 20070 20448 20076 20460
rect 18472 20420 19334 20448
rect 19905 20441 19963 20447
rect 18472 20408 18478 20420
rect 19905 20407 19917 20441
rect 19951 20438 19963 20441
rect 19996 20438 20076 20448
rect 19951 20420 20076 20438
rect 19951 20410 20024 20420
rect 19951 20407 19963 20410
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20448 20223 20451
rect 20438 20448 20444 20460
rect 20211 20420 20444 20448
rect 20211 20417 20223 20420
rect 20165 20411 20223 20417
rect 19905 20401 19963 20407
rect 10137 20383 10195 20389
rect 10137 20380 10149 20383
rect 9732 20352 10149 20380
rect 9732 20340 9738 20352
rect 10137 20349 10149 20352
rect 10183 20349 10195 20383
rect 10137 20343 10195 20349
rect 11609 20383 11667 20389
rect 11609 20349 11621 20383
rect 11655 20380 11667 20383
rect 12066 20380 12072 20392
rect 11655 20352 12072 20380
rect 11655 20349 11667 20352
rect 11609 20343 11667 20349
rect 12066 20340 12072 20352
rect 12124 20340 12130 20392
rect 12526 20340 12532 20392
rect 12584 20340 12590 20392
rect 14090 20340 14096 20392
rect 14148 20380 14154 20392
rect 14737 20383 14795 20389
rect 14737 20380 14749 20383
rect 14148 20352 14749 20380
rect 14148 20340 14154 20352
rect 14737 20349 14749 20352
rect 14783 20349 14795 20383
rect 14737 20343 14795 20349
rect 15010 20340 15016 20392
rect 15068 20340 15074 20392
rect 15654 20340 15660 20392
rect 15712 20340 15718 20392
rect 16758 20340 16764 20392
rect 16816 20380 16822 20392
rect 17034 20380 17040 20392
rect 16816 20352 17040 20380
rect 16816 20340 16822 20352
rect 17034 20340 17040 20352
rect 17092 20340 17098 20392
rect 16390 20312 16396 20324
rect 6972 20284 8248 20312
rect 16132 20284 16396 20312
rect 6972 20272 6978 20284
rect 16132 20256 16160 20284
rect 16390 20272 16396 20284
rect 16448 20272 16454 20324
rect 18138 20312 18144 20324
rect 16868 20284 18144 20312
rect 6733 20247 6791 20253
rect 6733 20213 6745 20247
rect 6779 20244 6791 20247
rect 7006 20244 7012 20256
rect 6779 20216 7012 20244
rect 6779 20213 6791 20216
rect 6733 20207 6791 20213
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 7190 20204 7196 20256
rect 7248 20204 7254 20256
rect 7374 20204 7380 20256
rect 7432 20204 7438 20256
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 9766 20244 9772 20256
rect 7524 20216 9772 20244
rect 7524 20204 7530 20216
rect 9766 20204 9772 20216
rect 9824 20204 9830 20256
rect 12161 20247 12219 20253
rect 12161 20213 12173 20247
rect 12207 20244 12219 20247
rect 12894 20244 12900 20256
rect 12207 20216 12900 20244
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 12894 20204 12900 20216
rect 12952 20204 12958 20256
rect 13262 20204 13268 20256
rect 13320 20204 13326 20256
rect 14550 20204 14556 20256
rect 14608 20244 14614 20256
rect 15105 20247 15163 20253
rect 15105 20244 15117 20247
rect 14608 20216 15117 20244
rect 14608 20204 14614 20216
rect 15105 20213 15117 20216
rect 15151 20213 15163 20247
rect 15105 20207 15163 20213
rect 15194 20204 15200 20256
rect 15252 20244 15258 20256
rect 16022 20244 16028 20256
rect 15252 20216 16028 20244
rect 15252 20204 15258 20216
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 16114 20204 16120 20256
rect 16172 20204 16178 20256
rect 16298 20204 16304 20256
rect 16356 20204 16362 20256
rect 16868 20253 16896 20284
rect 18138 20272 18144 20284
rect 18196 20272 18202 20324
rect 19334 20272 19340 20324
rect 19392 20312 19398 20324
rect 20180 20312 20208 20411
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 21450 20408 21456 20460
rect 21508 20448 21514 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21508 20420 22017 20448
rect 21508 20408 21514 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20448 22155 20451
rect 22370 20448 22376 20460
rect 22143 20420 22376 20448
rect 22143 20417 22155 20420
rect 22097 20411 22155 20417
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 22830 20408 22836 20460
rect 22888 20408 22894 20460
rect 22922 20408 22928 20460
rect 22980 20448 22986 20460
rect 23017 20451 23075 20457
rect 23017 20448 23029 20451
rect 22980 20420 23029 20448
rect 22980 20408 22986 20420
rect 23017 20417 23029 20420
rect 23063 20417 23075 20451
rect 23017 20411 23075 20417
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 24029 20451 24087 20457
rect 24029 20448 24041 20451
rect 23716 20420 24041 20448
rect 23716 20408 23722 20420
rect 24029 20417 24041 20420
rect 24075 20448 24087 20451
rect 24210 20448 24216 20460
rect 24075 20420 24216 20448
rect 24075 20417 24087 20420
rect 24029 20411 24087 20417
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 25516 20457 25544 20488
rect 25976 20460 26004 20488
rect 25133 20451 25191 20457
rect 25133 20417 25145 20451
rect 25179 20448 25191 20451
rect 25501 20451 25559 20457
rect 25179 20420 25452 20448
rect 25179 20417 25191 20420
rect 25133 20411 25191 20417
rect 21818 20340 21824 20392
rect 21876 20380 21882 20392
rect 23566 20380 23572 20392
rect 21876 20352 23572 20380
rect 21876 20340 21882 20352
rect 23566 20340 23572 20352
rect 23624 20340 23630 20392
rect 24302 20340 24308 20392
rect 24360 20380 24366 20392
rect 24762 20380 24768 20392
rect 24360 20352 24768 20380
rect 24360 20340 24366 20352
rect 24762 20340 24768 20352
rect 24820 20380 24826 20392
rect 25317 20383 25375 20389
rect 25317 20380 25329 20383
rect 24820 20352 25329 20380
rect 24820 20340 24826 20352
rect 25317 20349 25329 20352
rect 25363 20349 25375 20383
rect 25317 20343 25375 20349
rect 19392 20284 20208 20312
rect 21269 20315 21327 20321
rect 19392 20272 19398 20284
rect 21269 20281 21281 20315
rect 21315 20312 21327 20315
rect 21450 20312 21456 20324
rect 21315 20284 21456 20312
rect 21315 20281 21327 20284
rect 21269 20275 21327 20281
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 16853 20247 16911 20253
rect 16853 20213 16865 20247
rect 16899 20213 16911 20247
rect 16853 20207 16911 20213
rect 16942 20204 16948 20256
rect 17000 20244 17006 20256
rect 17037 20247 17095 20253
rect 17037 20244 17049 20247
rect 17000 20216 17049 20244
rect 17000 20204 17006 20216
rect 17037 20213 17049 20216
rect 17083 20213 17095 20247
rect 17037 20207 17095 20213
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 17313 20247 17371 20253
rect 17313 20244 17325 20247
rect 17276 20216 17325 20244
rect 17276 20204 17282 20216
rect 17313 20213 17325 20216
rect 17359 20213 17371 20247
rect 17313 20207 17371 20213
rect 17494 20204 17500 20256
rect 17552 20204 17558 20256
rect 21082 20204 21088 20256
rect 21140 20204 21146 20256
rect 21836 20253 21864 20340
rect 22002 20272 22008 20324
rect 22060 20312 22066 20324
rect 22833 20315 22891 20321
rect 22833 20312 22845 20315
rect 22060 20284 22845 20312
rect 22060 20272 22066 20284
rect 22833 20281 22845 20284
rect 22879 20281 22891 20315
rect 25424 20312 25452 20420
rect 25501 20417 25513 20451
rect 25547 20417 25559 20451
rect 25501 20411 25559 20417
rect 25682 20408 25688 20460
rect 25740 20408 25746 20460
rect 25774 20408 25780 20460
rect 25832 20408 25838 20460
rect 25869 20451 25927 20457
rect 25869 20417 25881 20451
rect 25915 20417 25927 20451
rect 25869 20411 25927 20417
rect 25884 20380 25912 20411
rect 25958 20408 25964 20460
rect 26016 20448 26022 20460
rect 26326 20457 26332 20460
rect 26145 20451 26203 20457
rect 26145 20448 26157 20451
rect 26016 20420 26157 20448
rect 26016 20408 26022 20420
rect 26145 20417 26157 20420
rect 26191 20417 26203 20451
rect 26145 20411 26203 20417
rect 26303 20451 26332 20457
rect 26303 20417 26315 20451
rect 26303 20411 26332 20417
rect 26326 20408 26332 20411
rect 26384 20408 26390 20460
rect 26418 20408 26424 20460
rect 26476 20408 26482 20460
rect 26510 20408 26516 20460
rect 26568 20408 26574 20460
rect 26620 20457 26648 20556
rect 26786 20476 26792 20528
rect 26844 20516 26850 20528
rect 27157 20519 27215 20525
rect 27157 20516 27169 20519
rect 26844 20488 27169 20516
rect 26844 20476 26850 20488
rect 27157 20485 27169 20488
rect 27203 20485 27215 20519
rect 27448 20516 27476 20556
rect 28166 20544 28172 20556
rect 28224 20544 28230 20596
rect 33870 20544 33876 20596
rect 33928 20584 33934 20596
rect 34977 20587 35035 20593
rect 34977 20584 34989 20587
rect 33928 20556 34989 20584
rect 33928 20544 33934 20556
rect 34977 20553 34989 20556
rect 35023 20553 35035 20587
rect 34977 20547 35035 20553
rect 27157 20479 27215 20485
rect 27356 20488 27476 20516
rect 27801 20519 27859 20525
rect 26605 20451 26663 20457
rect 26605 20417 26617 20451
rect 26651 20417 26663 20451
rect 26605 20411 26663 20417
rect 26973 20451 27031 20457
rect 26973 20417 26985 20451
rect 27019 20448 27031 20451
rect 27062 20448 27068 20460
rect 27019 20420 27068 20448
rect 27019 20417 27031 20420
rect 26973 20411 27031 20417
rect 26620 20380 26648 20411
rect 27062 20408 27068 20420
rect 27120 20408 27126 20460
rect 27246 20408 27252 20460
rect 27304 20408 27310 20460
rect 27356 20457 27384 20488
rect 27801 20485 27813 20519
rect 27847 20516 27859 20519
rect 28261 20519 28319 20525
rect 28261 20516 28273 20519
rect 27847 20488 28273 20516
rect 27847 20485 27859 20488
rect 27801 20479 27859 20485
rect 28261 20485 28273 20488
rect 28307 20485 28319 20519
rect 28261 20479 28319 20485
rect 27341 20451 27399 20457
rect 27341 20417 27353 20451
rect 27387 20417 27399 20451
rect 27341 20411 27399 20417
rect 27617 20451 27675 20457
rect 27617 20417 27629 20451
rect 27663 20417 27675 20451
rect 27617 20411 27675 20417
rect 25884 20352 26648 20380
rect 26789 20383 26847 20389
rect 26789 20349 26801 20383
rect 26835 20380 26847 20383
rect 27632 20380 27660 20411
rect 26835 20352 27660 20380
rect 26835 20349 26847 20352
rect 26789 20343 26847 20349
rect 26510 20312 26516 20324
rect 25424 20284 26516 20312
rect 22833 20275 22891 20281
rect 26510 20272 26516 20284
rect 26568 20272 26574 20324
rect 27525 20315 27583 20321
rect 27525 20281 27537 20315
rect 27571 20312 27583 20315
rect 27816 20312 27844 20479
rect 29362 20476 29368 20528
rect 29420 20516 29426 20528
rect 32582 20516 32588 20528
rect 29420 20488 32588 20516
rect 29420 20476 29426 20488
rect 32582 20476 32588 20488
rect 32640 20476 32646 20528
rect 28077 20451 28135 20457
rect 28077 20448 28089 20451
rect 27571 20284 27844 20312
rect 27908 20420 28089 20448
rect 27571 20281 27583 20284
rect 27525 20275 27583 20281
rect 21821 20247 21879 20253
rect 21821 20213 21833 20247
rect 21867 20213 21879 20247
rect 21821 20207 21879 20213
rect 26053 20247 26111 20253
rect 26053 20213 26065 20247
rect 26099 20244 26111 20247
rect 27706 20244 27712 20256
rect 26099 20216 27712 20244
rect 26099 20213 26111 20216
rect 26053 20207 26111 20213
rect 27706 20204 27712 20216
rect 27764 20244 27770 20256
rect 27908 20244 27936 20420
rect 28077 20417 28089 20420
rect 28123 20417 28135 20451
rect 28077 20411 28135 20417
rect 30282 20408 30288 20460
rect 30340 20408 30346 20460
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20448 30619 20451
rect 30650 20448 30656 20460
rect 30607 20420 30656 20448
rect 30607 20417 30619 20420
rect 30561 20411 30619 20417
rect 30650 20408 30656 20420
rect 30708 20408 30714 20460
rect 30742 20408 30748 20460
rect 30800 20448 30806 20460
rect 30929 20451 30987 20457
rect 30929 20448 30941 20451
rect 30800 20420 30941 20448
rect 30800 20408 30806 20420
rect 30929 20417 30941 20420
rect 30975 20417 30987 20451
rect 30929 20411 30987 20417
rect 31110 20408 31116 20460
rect 31168 20408 31174 20460
rect 31294 20408 31300 20460
rect 31352 20408 31358 20460
rect 31386 20408 31392 20460
rect 31444 20448 31450 20460
rect 34517 20451 34575 20457
rect 34517 20448 34529 20451
rect 31444 20420 34529 20448
rect 31444 20408 31450 20420
rect 34517 20417 34529 20420
rect 34563 20417 34575 20451
rect 34517 20411 34575 20417
rect 34793 20451 34851 20457
rect 34793 20417 34805 20451
rect 34839 20448 34851 20451
rect 35526 20448 35532 20460
rect 34839 20420 35532 20448
rect 34839 20417 34851 20420
rect 34793 20411 34851 20417
rect 35526 20408 35532 20420
rect 35584 20408 35590 20460
rect 27985 20383 28043 20389
rect 27985 20349 27997 20383
rect 28031 20380 28043 20383
rect 28442 20380 28448 20392
rect 28031 20352 28448 20380
rect 28031 20349 28043 20352
rect 27985 20343 28043 20349
rect 28442 20340 28448 20352
rect 28500 20340 28506 20392
rect 28810 20340 28816 20392
rect 28868 20380 28874 20392
rect 30377 20383 30435 20389
rect 30377 20380 30389 20383
rect 28868 20352 30389 20380
rect 28868 20340 28874 20352
rect 30377 20349 30389 20352
rect 30423 20349 30435 20383
rect 30668 20380 30696 20408
rect 31205 20383 31263 20389
rect 31205 20380 31217 20383
rect 30668 20352 31217 20380
rect 30377 20343 30435 20349
rect 31205 20349 31217 20352
rect 31251 20349 31263 20383
rect 31205 20343 31263 20349
rect 34606 20340 34612 20392
rect 34664 20340 34670 20392
rect 30745 20315 30803 20321
rect 30745 20281 30757 20315
rect 30791 20312 30803 20315
rect 34790 20312 34796 20324
rect 30791 20284 34796 20312
rect 30791 20281 30803 20284
rect 30745 20275 30803 20281
rect 34790 20272 34796 20284
rect 34848 20272 34854 20324
rect 27764 20216 27936 20244
rect 28445 20247 28503 20253
rect 27764 20204 27770 20216
rect 28445 20213 28457 20247
rect 28491 20244 28503 20247
rect 29546 20244 29552 20256
rect 28491 20216 29552 20244
rect 28491 20213 28503 20216
rect 28445 20207 28503 20213
rect 29546 20204 29552 20216
rect 29604 20204 29610 20256
rect 30466 20204 30472 20256
rect 30524 20204 30530 20256
rect 31202 20204 31208 20256
rect 31260 20244 31266 20256
rect 31389 20247 31447 20253
rect 31389 20244 31401 20247
rect 31260 20216 31401 20244
rect 31260 20204 31266 20216
rect 31389 20213 31401 20216
rect 31435 20213 31447 20247
rect 31389 20207 31447 20213
rect 31665 20247 31723 20253
rect 31665 20213 31677 20247
rect 31711 20244 31723 20247
rect 33962 20244 33968 20256
rect 31711 20216 33968 20244
rect 31711 20213 31723 20216
rect 31665 20207 31723 20213
rect 33962 20204 33968 20216
rect 34020 20204 34026 20256
rect 34514 20204 34520 20256
rect 34572 20204 34578 20256
rect 1104 20154 36432 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 36432 20154
rect 1104 20080 36432 20102
rect 4341 20043 4399 20049
rect 4341 20009 4353 20043
rect 4387 20040 4399 20043
rect 4890 20040 4896 20052
rect 4387 20012 4896 20040
rect 4387 20009 4399 20012
rect 4341 20003 4399 20009
rect 4890 20000 4896 20012
rect 4948 20000 4954 20052
rect 5169 20043 5227 20049
rect 5169 20009 5181 20043
rect 5215 20040 5227 20043
rect 6362 20040 6368 20052
rect 5215 20012 6368 20040
rect 5215 20009 5227 20012
rect 5169 20003 5227 20009
rect 6362 20000 6368 20012
rect 6420 20000 6426 20052
rect 6638 20000 6644 20052
rect 6696 20000 6702 20052
rect 6904 20043 6962 20049
rect 6904 20009 6916 20043
rect 6950 20040 6962 20043
rect 7374 20040 7380 20052
rect 6950 20012 7380 20040
rect 6950 20009 6962 20012
rect 6904 20003 6962 20009
rect 7374 20000 7380 20012
rect 7432 20000 7438 20052
rect 8386 20000 8392 20052
rect 8444 20000 8450 20052
rect 8478 20000 8484 20052
rect 8536 20040 8542 20052
rect 8573 20043 8631 20049
rect 8573 20040 8585 20043
rect 8536 20012 8585 20040
rect 8536 20000 8542 20012
rect 8573 20009 8585 20012
rect 8619 20040 8631 20043
rect 9122 20040 9128 20052
rect 8619 20012 9128 20040
rect 8619 20009 8631 20012
rect 8573 20003 8631 20009
rect 9122 20000 9128 20012
rect 9180 20000 9186 20052
rect 9582 20000 9588 20052
rect 9640 20040 9646 20052
rect 9950 20040 9956 20052
rect 9640 20012 9956 20040
rect 9640 20000 9646 20012
rect 9950 20000 9956 20012
rect 10008 20040 10014 20052
rect 11054 20040 11060 20052
rect 10008 20012 11060 20040
rect 10008 20000 10014 20012
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 11425 20043 11483 20049
rect 11425 20009 11437 20043
rect 11471 20040 11483 20043
rect 11790 20040 11796 20052
rect 11471 20012 11796 20040
rect 11471 20009 11483 20012
rect 11425 20003 11483 20009
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 13630 20040 13636 20052
rect 12584 20012 13636 20040
rect 12584 20000 12590 20012
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14332 20012 15516 20040
rect 14332 20000 14338 20012
rect 6656 19972 6684 20000
rect 5920 19944 6684 19972
rect 4430 19904 4436 19916
rect 3988 19876 4436 19904
rect 1394 19796 1400 19848
rect 1452 19796 1458 19848
rect 3694 19796 3700 19848
rect 3752 19836 3758 19848
rect 3988 19845 4016 19876
rect 4430 19864 4436 19876
rect 4488 19864 4494 19916
rect 5074 19864 5080 19916
rect 5132 19864 5138 19916
rect 5920 19913 5948 19944
rect 8202 19932 8208 19984
rect 8260 19972 8266 19984
rect 14292 19972 14320 20000
rect 8260 19944 9720 19972
rect 8260 19932 8266 19944
rect 6362 19913 6368 19916
rect 5905 19907 5963 19913
rect 5905 19873 5917 19907
rect 5951 19873 5963 19907
rect 5905 19867 5963 19873
rect 6319 19907 6368 19913
rect 6319 19873 6331 19907
rect 6365 19873 6368 19907
rect 6319 19867 6368 19873
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 3752 19808 3801 19836
rect 3752 19796 3758 19808
rect 3789 19805 3801 19808
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4246 19836 4252 19848
rect 4203 19808 4252 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 5596 19839 5654 19845
rect 5596 19805 5608 19839
rect 5642 19836 5654 19839
rect 5920 19836 5948 19867
rect 6362 19864 6368 19867
rect 6420 19864 6426 19916
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 6914 19904 6920 19916
rect 6687 19876 6920 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 8846 19904 8852 19916
rect 7340 19876 8852 19904
rect 7340 19864 7346 19876
rect 8846 19864 8852 19876
rect 8904 19864 8910 19916
rect 9692 19913 9720 19944
rect 13280 19944 14320 19972
rect 9401 19907 9459 19913
rect 9401 19904 9413 19907
rect 9324 19876 9413 19904
rect 9324 19848 9352 19876
rect 9401 19873 9413 19876
rect 9447 19873 9459 19907
rect 9401 19867 9459 19873
rect 9677 19907 9735 19913
rect 9677 19873 9689 19907
rect 9723 19904 9735 19907
rect 11885 19907 11943 19913
rect 11885 19904 11897 19907
rect 9723 19876 11897 19904
rect 9723 19873 9735 19876
rect 9677 19867 9735 19873
rect 11885 19873 11897 19876
rect 11931 19873 11943 19907
rect 11885 19867 11943 19873
rect 12161 19907 12219 19913
rect 12161 19873 12173 19907
rect 12207 19904 12219 19907
rect 12250 19904 12256 19916
rect 12207 19876 12256 19904
rect 12207 19873 12219 19876
rect 12161 19867 12219 19873
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 12526 19864 12532 19916
rect 12584 19904 12590 19916
rect 13280 19904 13308 19944
rect 12584 19876 13308 19904
rect 12584 19864 12590 19876
rect 5642 19808 5948 19836
rect 5642 19805 5654 19808
rect 5596 19799 5654 19805
rect 6178 19796 6184 19848
rect 6236 19796 6242 19848
rect 8478 19796 8484 19848
rect 8536 19796 8542 19848
rect 8665 19839 8723 19845
rect 8665 19805 8677 19839
rect 8711 19836 8723 19839
rect 8938 19836 8944 19848
rect 8711 19808 8944 19836
rect 8711 19805 8723 19808
rect 8665 19799 8723 19805
rect 1670 19728 1676 19780
rect 1728 19728 1734 19780
rect 2958 19768 2964 19780
rect 2898 19740 2964 19768
rect 2958 19728 2964 19740
rect 3016 19728 3022 19780
rect 4065 19771 4123 19777
rect 4065 19737 4077 19771
rect 4111 19737 4123 19771
rect 4065 19731 4123 19737
rect 3145 19703 3203 19709
rect 3145 19669 3157 19703
rect 3191 19700 3203 19703
rect 3418 19700 3424 19712
rect 3191 19672 3424 19700
rect 3191 19669 3203 19672
rect 3145 19663 3203 19669
rect 3418 19660 3424 19672
rect 3476 19700 3482 19712
rect 4080 19700 4108 19731
rect 4338 19728 4344 19780
rect 4396 19768 4402 19780
rect 5813 19771 5871 19777
rect 5813 19768 5825 19771
rect 4396 19740 5825 19768
rect 4396 19728 4402 19740
rect 5813 19737 5825 19740
rect 5859 19737 5871 19771
rect 6822 19768 6828 19780
rect 5813 19731 5871 19737
rect 6380 19740 6828 19768
rect 3476 19672 4108 19700
rect 3476 19660 3482 19672
rect 5534 19660 5540 19712
rect 5592 19660 5598 19712
rect 5721 19703 5779 19709
rect 5721 19669 5733 19703
rect 5767 19700 5779 19703
rect 6380 19700 6408 19740
rect 6822 19728 6828 19740
rect 6880 19728 6886 19780
rect 7116 19740 7406 19768
rect 7116 19712 7144 19740
rect 5767 19672 6408 19700
rect 6457 19703 6515 19709
rect 5767 19669 5779 19672
rect 5721 19663 5779 19669
rect 6457 19669 6469 19703
rect 6503 19700 6515 19703
rect 6546 19700 6552 19712
rect 6503 19672 6552 19700
rect 6503 19669 6515 19672
rect 6457 19663 6515 19669
rect 6546 19660 6552 19672
rect 6604 19660 6610 19712
rect 7098 19660 7104 19712
rect 7156 19660 7162 19712
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 8680 19700 8708 19799
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 8846 19728 8852 19780
rect 8904 19768 8910 19780
rect 9232 19768 9260 19799
rect 9306 19796 9312 19848
rect 9364 19796 9370 19848
rect 9493 19839 9551 19845
rect 9493 19836 9505 19839
rect 9416 19808 9505 19836
rect 9416 19780 9444 19808
rect 9493 19805 9505 19808
rect 9539 19805 9551 19839
rect 13280 19822 13308 19876
rect 14185 19907 14243 19913
rect 14185 19873 14197 19907
rect 14231 19904 14243 19907
rect 15010 19904 15016 19916
rect 14231 19876 15016 19904
rect 14231 19873 14243 19876
rect 14185 19867 14243 19873
rect 15010 19864 15016 19876
rect 15068 19864 15074 19916
rect 15488 19904 15516 20012
rect 15930 20000 15936 20052
rect 15988 20000 15994 20052
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 17402 20040 17408 20052
rect 16632 20012 17408 20040
rect 16632 20000 16638 20012
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 20254 20000 20260 20052
rect 20312 20040 20318 20052
rect 20533 20043 20591 20049
rect 20533 20040 20545 20043
rect 20312 20012 20545 20040
rect 20312 20000 20318 20012
rect 20533 20009 20545 20012
rect 20579 20040 20591 20043
rect 22094 20040 22100 20052
rect 20579 20012 22100 20040
rect 20579 20009 20591 20012
rect 20533 20003 20591 20009
rect 22094 20000 22100 20012
rect 22152 20000 22158 20052
rect 26050 20000 26056 20052
rect 26108 20040 26114 20052
rect 27246 20040 27252 20052
rect 26108 20012 27252 20040
rect 26108 20000 26114 20012
rect 27246 20000 27252 20012
rect 27304 20000 27310 20052
rect 28353 20043 28411 20049
rect 28353 20009 28365 20043
rect 28399 20040 28411 20043
rect 28810 20040 28816 20052
rect 28399 20012 28816 20040
rect 28399 20009 28411 20012
rect 28353 20003 28411 20009
rect 28810 20000 28816 20012
rect 28868 20000 28874 20052
rect 29546 20000 29552 20052
rect 29604 20000 29610 20052
rect 30009 20043 30067 20049
rect 30009 20009 30021 20043
rect 30055 20040 30067 20043
rect 31386 20040 31392 20052
rect 30055 20012 31392 20040
rect 30055 20009 30067 20012
rect 30009 20003 30067 20009
rect 31386 20000 31392 20012
rect 31444 20000 31450 20052
rect 33686 20000 33692 20052
rect 33744 20040 33750 20052
rect 33873 20043 33931 20049
rect 33873 20040 33885 20043
rect 33744 20012 33885 20040
rect 33744 20000 33750 20012
rect 33873 20009 33885 20012
rect 33919 20009 33931 20043
rect 33873 20003 33931 20009
rect 15654 19932 15660 19984
rect 15712 19972 15718 19984
rect 19978 19972 19984 19984
rect 15712 19944 19984 19972
rect 15712 19932 15718 19944
rect 19978 19932 19984 19944
rect 20036 19932 20042 19984
rect 21542 19932 21548 19984
rect 21600 19972 21606 19984
rect 21729 19975 21787 19981
rect 21729 19972 21741 19975
rect 21600 19944 21741 19972
rect 21600 19932 21606 19944
rect 21729 19941 21741 19944
rect 21775 19941 21787 19975
rect 21729 19935 21787 19941
rect 26418 19932 26424 19984
rect 26476 19972 26482 19984
rect 31018 19972 31024 19984
rect 26476 19944 31024 19972
rect 26476 19932 26482 19944
rect 31018 19932 31024 19944
rect 31076 19932 31082 19984
rect 15488 19876 15700 19904
rect 9493 19799 9551 19805
rect 8904 19740 9260 19768
rect 8904 19728 8910 19740
rect 9398 19728 9404 19780
rect 9456 19728 9462 19780
rect 9953 19771 10011 19777
rect 9953 19737 9965 19771
rect 9999 19768 10011 19771
rect 10226 19768 10232 19780
rect 9999 19740 10232 19768
rect 9999 19737 10011 19740
rect 9953 19731 10011 19737
rect 10226 19728 10232 19740
rect 10284 19728 10290 19780
rect 14461 19771 14519 19777
rect 10336 19740 10442 19768
rect 7340 19672 8708 19700
rect 7340 19660 7346 19672
rect 8938 19660 8944 19712
rect 8996 19660 9002 19712
rect 9214 19660 9220 19712
rect 9272 19700 9278 19712
rect 10042 19700 10048 19712
rect 9272 19672 10048 19700
rect 9272 19660 9278 19672
rect 10042 19660 10048 19672
rect 10100 19700 10106 19712
rect 10336 19700 10364 19740
rect 14461 19737 14473 19771
rect 14507 19768 14519 19771
rect 14550 19768 14556 19780
rect 14507 19740 14556 19768
rect 14507 19737 14519 19740
rect 14461 19731 14519 19737
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 15672 19768 15700 19876
rect 16114 19864 16120 19916
rect 16172 19864 16178 19916
rect 16209 19907 16267 19913
rect 16209 19873 16221 19907
rect 16255 19904 16267 19907
rect 17862 19904 17868 19916
rect 16255 19876 17868 19904
rect 16255 19873 16267 19876
rect 16209 19867 16267 19873
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16301 19839 16359 19845
rect 16301 19836 16313 19839
rect 15988 19808 16313 19836
rect 15988 19796 15994 19808
rect 16301 19805 16313 19808
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 16390 19796 16396 19848
rect 16448 19796 16454 19848
rect 17126 19836 17132 19848
rect 16500 19808 17132 19836
rect 16500 19768 16528 19808
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17236 19845 17264 19876
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 18138 19864 18144 19916
rect 18196 19904 18202 19916
rect 19058 19904 19064 19916
rect 18196 19876 19064 19904
rect 18196 19864 18202 19876
rect 19058 19864 19064 19876
rect 19116 19904 19122 19916
rect 20806 19904 20812 19916
rect 19116 19876 20812 19904
rect 19116 19864 19122 19876
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 20898 19864 20904 19916
rect 20956 19904 20962 19916
rect 22646 19904 22652 19916
rect 20956 19876 21312 19904
rect 20956 19864 20962 19876
rect 17221 19839 17279 19845
rect 17221 19805 17233 19839
rect 17267 19805 17279 19839
rect 17221 19799 17279 19805
rect 15672 19754 16528 19768
rect 15686 19740 16528 19754
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 16853 19771 16911 19777
rect 16853 19768 16865 19771
rect 16816 19740 16865 19768
rect 16816 19728 16822 19740
rect 16853 19737 16865 19740
rect 16899 19737 16911 19771
rect 16853 19731 16911 19737
rect 17034 19728 17040 19780
rect 17092 19768 17098 19780
rect 17678 19768 17684 19780
rect 17092 19740 17684 19768
rect 17092 19728 17098 19740
rect 17678 19728 17684 19740
rect 17736 19728 17742 19780
rect 18156 19768 18184 19864
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19836 18291 19839
rect 18322 19836 18328 19848
rect 18279 19808 18328 19836
rect 18279 19805 18291 19808
rect 18233 19799 18291 19805
rect 18322 19796 18328 19808
rect 18380 19836 18386 19848
rect 18506 19836 18512 19848
rect 18380 19808 18512 19836
rect 18380 19796 18386 19808
rect 18506 19796 18512 19808
rect 18564 19796 18570 19848
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21284 19845 21312 19876
rect 21376 19876 22652 19904
rect 21376 19848 21404 19876
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 25685 19907 25743 19913
rect 25685 19873 25697 19907
rect 25731 19904 25743 19907
rect 26510 19904 26516 19916
rect 25731 19876 26516 19904
rect 25731 19873 25743 19876
rect 25685 19867 25743 19873
rect 21085 19839 21143 19845
rect 21085 19836 21097 19839
rect 21048 19808 21097 19836
rect 21048 19796 21054 19808
rect 21085 19805 21097 19808
rect 21131 19805 21143 19839
rect 21085 19799 21143 19805
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 18417 19771 18475 19777
rect 18417 19768 18429 19771
rect 18156 19740 18429 19768
rect 18417 19737 18429 19740
rect 18463 19737 18475 19771
rect 18966 19768 18972 19780
rect 18417 19731 18475 19737
rect 18524 19740 18972 19768
rect 10100 19672 10364 19700
rect 10100 19660 10106 19672
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 14366 19700 14372 19712
rect 12124 19672 14372 19700
rect 12124 19660 12130 19672
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 16022 19700 16028 19712
rect 15160 19672 16028 19700
rect 15160 19660 15166 19672
rect 16022 19660 16028 19672
rect 16080 19660 16086 19712
rect 16666 19660 16672 19712
rect 16724 19700 16730 19712
rect 17052 19700 17080 19728
rect 16724 19672 17080 19700
rect 16724 19660 16730 19672
rect 17126 19660 17132 19712
rect 17184 19700 17190 19712
rect 18524 19700 18552 19740
rect 18966 19728 18972 19740
rect 19024 19728 19030 19780
rect 19242 19728 19248 19780
rect 19300 19728 19306 19780
rect 19702 19728 19708 19780
rect 19760 19768 19766 19780
rect 20254 19768 20260 19780
rect 19760 19740 20260 19768
rect 19760 19728 19766 19740
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 21100 19768 21128 19799
rect 21358 19796 21364 19848
rect 21416 19796 21422 19848
rect 21450 19796 21456 19848
rect 21508 19836 21514 19848
rect 25700 19836 25728 19867
rect 26510 19864 26516 19876
rect 26568 19864 26574 19916
rect 29362 19904 29368 19916
rect 28000 19876 29368 19904
rect 21508 19808 25728 19836
rect 25869 19839 25927 19845
rect 21508 19796 21514 19808
rect 25869 19805 25881 19839
rect 25915 19836 25927 19839
rect 25958 19836 25964 19848
rect 25915 19808 25964 19836
rect 25915 19805 25927 19808
rect 25869 19799 25927 19805
rect 25958 19796 25964 19808
rect 26016 19796 26022 19848
rect 27798 19796 27804 19848
rect 27856 19796 27862 19848
rect 28000 19845 28028 19876
rect 29362 19864 29368 19876
rect 29420 19864 29426 19916
rect 29730 19864 29736 19916
rect 29788 19864 29794 19916
rect 33962 19864 33968 19916
rect 34020 19864 34026 19916
rect 35250 19864 35256 19916
rect 35308 19904 35314 19916
rect 35526 19904 35532 19916
rect 35308 19876 35532 19904
rect 35308 19864 35314 19876
rect 35526 19864 35532 19876
rect 35584 19864 35590 19916
rect 27985 19839 28043 19845
rect 27985 19805 27997 19839
rect 28031 19805 28043 19839
rect 27985 19799 28043 19805
rect 28166 19796 28172 19848
rect 28224 19796 28230 19848
rect 29270 19796 29276 19848
rect 29328 19836 29334 19848
rect 29825 19839 29883 19845
rect 29825 19836 29837 19839
rect 29328 19808 29837 19836
rect 29328 19796 29334 19808
rect 29825 19805 29837 19808
rect 29871 19805 29883 19839
rect 29825 19799 29883 19805
rect 34146 19796 34152 19848
rect 34204 19796 34210 19848
rect 23474 19768 23480 19780
rect 21100 19740 23480 19768
rect 23474 19728 23480 19740
rect 23532 19728 23538 19780
rect 28077 19771 28135 19777
rect 28077 19737 28089 19771
rect 28123 19737 28135 19771
rect 28077 19731 28135 19737
rect 17184 19672 18552 19700
rect 17184 19660 17190 19672
rect 18598 19660 18604 19712
rect 18656 19660 18662 19712
rect 18690 19660 18696 19712
rect 18748 19700 18754 19712
rect 23382 19700 23388 19712
rect 18748 19672 23388 19700
rect 18748 19660 18754 19672
rect 23382 19660 23388 19672
rect 23440 19660 23446 19712
rect 26786 19660 26792 19712
rect 26844 19700 26850 19712
rect 28092 19700 28120 19731
rect 28534 19728 28540 19780
rect 28592 19768 28598 19780
rect 29549 19771 29607 19777
rect 29549 19768 29561 19771
rect 28592 19740 29561 19768
rect 28592 19728 28598 19740
rect 29549 19737 29561 19740
rect 29595 19737 29607 19771
rect 29549 19731 29607 19737
rect 33873 19771 33931 19777
rect 33873 19737 33885 19771
rect 33919 19768 33931 19771
rect 33962 19768 33968 19780
rect 33919 19740 33968 19768
rect 33919 19737 33931 19740
rect 33873 19731 33931 19737
rect 33962 19728 33968 19740
rect 34020 19728 34026 19780
rect 26844 19672 28120 19700
rect 26844 19660 26850 19672
rect 34146 19660 34152 19712
rect 34204 19700 34210 19712
rect 34333 19703 34391 19709
rect 34333 19700 34345 19703
rect 34204 19672 34345 19700
rect 34204 19660 34210 19672
rect 34333 19669 34345 19672
rect 34379 19669 34391 19703
rect 34333 19663 34391 19669
rect 1104 19610 36432 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 36432 19610
rect 1104 19536 36432 19558
rect 1670 19456 1676 19508
rect 1728 19496 1734 19508
rect 2041 19499 2099 19505
rect 2041 19496 2053 19499
rect 1728 19468 2053 19496
rect 1728 19456 1734 19468
rect 2041 19465 2053 19468
rect 2087 19465 2099 19499
rect 2041 19459 2099 19465
rect 2130 19456 2136 19508
rect 2188 19496 2194 19508
rect 2501 19499 2559 19505
rect 2501 19496 2513 19499
rect 2188 19468 2513 19496
rect 2188 19456 2194 19468
rect 2501 19465 2513 19468
rect 2547 19496 2559 19499
rect 2590 19496 2596 19508
rect 2547 19468 2596 19496
rect 2547 19465 2559 19468
rect 2501 19459 2559 19465
rect 2590 19456 2596 19468
rect 2648 19456 2654 19508
rect 3510 19456 3516 19508
rect 3568 19496 3574 19508
rect 4062 19496 4068 19508
rect 3568 19468 4068 19496
rect 3568 19456 3574 19468
rect 4062 19456 4068 19468
rect 4120 19496 4126 19508
rect 4338 19496 4344 19508
rect 4120 19468 4344 19496
rect 4120 19456 4126 19468
rect 4338 19456 4344 19468
rect 4396 19456 4402 19508
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 4890 19496 4896 19508
rect 4488 19468 4896 19496
rect 4488 19456 4494 19468
rect 4890 19456 4896 19468
rect 4948 19456 4954 19508
rect 7282 19496 7288 19508
rect 5828 19468 7288 19496
rect 5828 19440 5856 19468
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 7616 19468 8754 19496
rect 7616 19456 7622 19468
rect 3326 19388 3332 19440
rect 3384 19428 3390 19440
rect 3789 19431 3847 19437
rect 3789 19428 3801 19431
rect 3384 19400 3801 19428
rect 3384 19388 3390 19400
rect 3789 19397 3801 19400
rect 3835 19428 3847 19431
rect 4706 19428 4712 19440
rect 3835 19400 4712 19428
rect 3835 19397 3847 19400
rect 3789 19391 3847 19397
rect 4706 19388 4712 19400
rect 4764 19388 4770 19440
rect 5810 19388 5816 19440
rect 5868 19388 5874 19440
rect 6914 19428 6920 19440
rect 6380 19400 6920 19428
rect 2409 19363 2467 19369
rect 2409 19329 2421 19363
rect 2455 19360 2467 19363
rect 2869 19363 2927 19369
rect 2869 19360 2881 19363
rect 2455 19332 2881 19360
rect 2455 19329 2467 19332
rect 2409 19323 2467 19329
rect 2869 19329 2881 19332
rect 2915 19329 2927 19363
rect 2869 19323 2927 19329
rect 3418 19320 3424 19372
rect 3476 19320 3482 19372
rect 3602 19320 3608 19372
rect 3660 19320 3666 19372
rect 3878 19320 3884 19372
rect 3936 19320 3942 19372
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19360 4031 19363
rect 4246 19360 4252 19372
rect 4019 19332 4252 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 4246 19320 4252 19332
rect 4304 19360 4310 19372
rect 4982 19360 4988 19372
rect 4304 19332 4988 19360
rect 4304 19320 4310 19332
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 5442 19320 5448 19372
rect 5500 19320 5506 19372
rect 6380 19369 6408 19400
rect 6914 19388 6920 19400
rect 6972 19388 6978 19440
rect 7926 19428 7932 19440
rect 7866 19400 7932 19428
rect 7926 19388 7932 19400
rect 7984 19388 7990 19440
rect 8386 19428 8392 19440
rect 8128 19400 8392 19428
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 2590 19252 2596 19304
rect 2648 19252 2654 19304
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19292 5687 19295
rect 5718 19292 5724 19304
rect 5675 19264 5724 19292
rect 5675 19261 5687 19264
rect 5629 19255 5687 19261
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 6730 19292 6736 19304
rect 6687 19264 6736 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 6730 19252 6736 19264
rect 6788 19252 6794 19304
rect 8128 19301 8156 19400
rect 8386 19388 8392 19400
rect 8444 19428 8450 19440
rect 8573 19431 8631 19437
rect 8573 19428 8585 19431
rect 8444 19400 8585 19428
rect 8444 19388 8450 19400
rect 8573 19397 8585 19400
rect 8619 19397 8631 19431
rect 8573 19391 8631 19397
rect 8202 19320 8208 19372
rect 8260 19320 8266 19372
rect 8294 19320 8300 19372
rect 8352 19320 8358 19372
rect 8726 19369 8754 19468
rect 9227 19468 10088 19496
rect 9227 19391 9255 19468
rect 9309 19431 9367 19437
rect 9309 19397 9321 19431
rect 9355 19428 9367 19431
rect 10060 19428 10088 19468
rect 10226 19456 10232 19508
rect 10284 19456 10290 19508
rect 12434 19496 12440 19508
rect 10520 19468 12440 19496
rect 10318 19428 10324 19440
rect 9355 19400 9996 19428
rect 10060 19400 10324 19428
rect 9355 19397 9367 19400
rect 9309 19391 9367 19397
rect 9212 19385 9270 19391
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19360 8539 19363
rect 8711 19363 8769 19369
rect 8527 19332 8616 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 8113 19295 8171 19301
rect 8113 19261 8125 19295
rect 8159 19261 8171 19295
rect 8113 19255 8171 19261
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 8588 19224 8616 19332
rect 8711 19329 8723 19363
rect 8757 19360 8769 19363
rect 9212 19360 9224 19385
rect 8757 19351 9224 19360
rect 9258 19351 9270 19385
rect 8757 19345 9270 19351
rect 8757 19332 9255 19345
rect 8757 19329 8769 19332
rect 8711 19323 8769 19329
rect 9398 19320 9404 19372
rect 9456 19320 9462 19372
rect 9539 19363 9597 19369
rect 9539 19329 9551 19363
rect 9585 19360 9597 19363
rect 9674 19360 9680 19372
rect 9585 19332 9680 19360
rect 9585 19329 9597 19332
rect 9539 19323 9597 19329
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 9272 19264 9321 19292
rect 9272 19252 9278 19264
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 9766 19252 9772 19304
rect 9824 19252 9830 19304
rect 9968 19292 9996 19400
rect 10318 19388 10324 19400
rect 10376 19388 10382 19440
rect 10042 19320 10048 19372
rect 10100 19360 10106 19372
rect 10520 19360 10548 19468
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 14182 19496 14188 19508
rect 12544 19468 14188 19496
rect 10689 19431 10747 19437
rect 10689 19397 10701 19431
rect 10735 19428 10747 19431
rect 10778 19428 10784 19440
rect 10735 19400 10784 19428
rect 10735 19397 10747 19400
rect 10689 19391 10747 19397
rect 10778 19388 10784 19400
rect 10836 19388 10842 19440
rect 12345 19431 12403 19437
rect 12345 19397 12357 19431
rect 12391 19428 12403 19431
rect 12544 19428 12572 19468
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 14366 19456 14372 19508
rect 14424 19496 14430 19508
rect 15866 19499 15924 19505
rect 15866 19496 15878 19499
rect 14424 19468 15878 19496
rect 14424 19456 14430 19468
rect 15866 19465 15878 19468
rect 15912 19465 15924 19499
rect 15866 19459 15924 19465
rect 16390 19456 16396 19508
rect 16448 19496 16454 19508
rect 18414 19496 18420 19508
rect 16448 19468 18420 19496
rect 16448 19456 16454 19468
rect 18414 19456 18420 19468
rect 18472 19456 18478 19508
rect 18509 19499 18567 19505
rect 18509 19465 18521 19499
rect 18555 19496 18567 19499
rect 18782 19496 18788 19508
rect 18555 19468 18788 19496
rect 18555 19465 18567 19468
rect 18509 19459 18567 19465
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 19153 19499 19211 19505
rect 19153 19465 19165 19499
rect 19199 19496 19211 19499
rect 19334 19496 19340 19508
rect 19199 19468 19340 19496
rect 19199 19465 19211 19468
rect 19153 19459 19211 19465
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 19886 19496 19892 19508
rect 19843 19468 19892 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 19886 19456 19892 19468
rect 19944 19456 19950 19508
rect 19978 19456 19984 19508
rect 20036 19496 20042 19508
rect 22465 19499 22523 19505
rect 22465 19496 22477 19499
rect 20036 19468 22477 19496
rect 20036 19456 20042 19468
rect 22465 19465 22477 19468
rect 22511 19465 22523 19499
rect 22465 19459 22523 19465
rect 22554 19456 22560 19508
rect 22612 19456 22618 19508
rect 23109 19499 23167 19505
rect 23109 19465 23121 19499
rect 23155 19496 23167 19499
rect 23198 19496 23204 19508
rect 23155 19468 23204 19496
rect 23155 19465 23167 19468
rect 23109 19459 23167 19465
rect 23198 19456 23204 19468
rect 23256 19456 23262 19508
rect 24397 19499 24455 19505
rect 24397 19465 24409 19499
rect 24443 19496 24455 19499
rect 24670 19496 24676 19508
rect 24443 19468 24676 19496
rect 24443 19465 24455 19468
rect 24397 19459 24455 19465
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 30374 19496 30380 19508
rect 25516 19468 30380 19496
rect 13538 19428 13544 19440
rect 12391 19400 12572 19428
rect 12636 19400 13544 19428
rect 12391 19397 12403 19400
rect 12345 19391 12403 19397
rect 12636 19372 12664 19400
rect 13538 19388 13544 19400
rect 13596 19388 13602 19440
rect 13630 19388 13636 19440
rect 13688 19388 13694 19440
rect 13906 19388 13912 19440
rect 13964 19428 13970 19440
rect 14274 19428 14280 19440
rect 13964 19400 14044 19428
rect 13964 19388 13970 19400
rect 10100 19332 10548 19360
rect 10597 19363 10655 19369
rect 10100 19320 10106 19332
rect 10597 19329 10609 19363
rect 10643 19360 10655 19363
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 10643 19332 11529 19360
rect 10643 19329 10655 19332
rect 10597 19323 10655 19329
rect 11517 19329 11529 19332
rect 11563 19329 11575 19363
rect 11517 19323 11575 19329
rect 11790 19320 11796 19372
rect 11848 19360 11854 19372
rect 12069 19363 12127 19369
rect 12069 19360 12081 19363
rect 11848 19332 12081 19360
rect 11848 19320 11854 19332
rect 12069 19329 12081 19332
rect 12115 19329 12127 19363
rect 12069 19323 12127 19329
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19360 12587 19363
rect 12618 19360 12624 19372
rect 12575 19332 12624 19360
rect 12575 19329 12587 19332
rect 12529 19323 12587 19329
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13170 19360 13176 19372
rect 12759 19332 13176 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 13262 19320 13268 19372
rect 13320 19360 13326 19372
rect 13449 19363 13507 19369
rect 13449 19360 13461 19363
rect 13320 19332 13461 19360
rect 13320 19320 13326 19332
rect 13449 19329 13461 19332
rect 13495 19360 13507 19363
rect 13495 19332 13584 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 10686 19292 10692 19304
rect 9968 19264 10692 19292
rect 10686 19252 10692 19264
rect 10744 19252 10750 19304
rect 10870 19252 10876 19304
rect 10928 19252 10934 19304
rect 12802 19252 12808 19304
rect 12860 19292 12866 19304
rect 13081 19295 13139 19301
rect 13081 19292 13093 19295
rect 12860 19264 13093 19292
rect 12860 19252 12866 19264
rect 13081 19261 13093 19264
rect 13127 19261 13139 19295
rect 13081 19255 13139 19261
rect 8754 19224 8760 19236
rect 8352 19196 8760 19224
rect 8352 19184 8358 19196
rect 8754 19184 8760 19196
rect 8812 19224 8818 19236
rect 8812 19196 9633 19224
rect 8812 19184 8818 19196
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4614 19156 4620 19168
rect 4203 19128 4620 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 5721 19159 5779 19165
rect 5721 19125 5733 19159
rect 5767 19156 5779 19159
rect 7190 19156 7196 19168
rect 5767 19128 7196 19156
rect 5767 19125 5779 19128
rect 5721 19119 5779 19125
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 8662 19116 8668 19168
rect 8720 19156 8726 19168
rect 8849 19159 8907 19165
rect 8849 19156 8861 19159
rect 8720 19128 8861 19156
rect 8720 19116 8726 19128
rect 8849 19125 8861 19128
rect 8895 19125 8907 19159
rect 9605 19156 9633 19196
rect 11882 19184 11888 19236
rect 11940 19224 11946 19236
rect 13446 19224 13452 19236
rect 11940 19196 13452 19224
rect 11940 19184 11946 19196
rect 13446 19184 13452 19196
rect 13504 19184 13510 19236
rect 13556 19224 13584 19332
rect 13648 19292 13676 19388
rect 13909 19295 13967 19301
rect 13909 19292 13921 19295
rect 13648 19264 13921 19292
rect 13909 19261 13921 19264
rect 13955 19261 13967 19295
rect 13909 19255 13967 19261
rect 13814 19224 13820 19236
rect 13556 19196 13820 19224
rect 13814 19184 13820 19196
rect 13872 19184 13878 19236
rect 14016 19224 14044 19400
rect 14108 19400 14280 19428
rect 14108 19372 14136 19400
rect 14274 19388 14280 19400
rect 14332 19388 14338 19440
rect 16206 19428 16212 19440
rect 15488 19400 16212 19428
rect 14090 19320 14096 19372
rect 14148 19320 14154 19372
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19360 14427 19363
rect 14550 19360 14556 19372
rect 14415 19332 14556 19360
rect 14415 19329 14427 19332
rect 14369 19323 14427 19329
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 14645 19363 14703 19369
rect 14645 19329 14657 19363
rect 14691 19360 14703 19363
rect 15194 19360 15200 19372
rect 14691 19332 15200 19360
rect 14691 19329 14703 19332
rect 14645 19323 14703 19329
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15488 19369 15516 19400
rect 16206 19388 16212 19400
rect 16264 19388 16270 19440
rect 16316 19400 17080 19428
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 16316 19369 16344 19400
rect 15749 19363 15807 19369
rect 15749 19360 15761 19363
rect 15620 19332 15761 19360
rect 15620 19320 15626 19332
rect 15749 19329 15761 19332
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 14332 19264 14473 19292
rect 14332 19252 14338 19264
rect 14461 19261 14473 19264
rect 14507 19261 14519 19295
rect 16758 19292 16764 19304
rect 16422 19264 16764 19292
rect 14461 19255 14519 19261
rect 16758 19252 16764 19264
rect 16816 19292 16822 19304
rect 16853 19295 16911 19301
rect 16853 19292 16865 19295
rect 16816 19264 16865 19292
rect 16816 19252 16822 19264
rect 16853 19261 16865 19264
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 14369 19227 14427 19233
rect 14369 19224 14381 19227
rect 14016 19196 14381 19224
rect 14369 19193 14381 19196
rect 14415 19193 14427 19227
rect 17052 19224 17080 19400
rect 18598 19388 18604 19440
rect 18656 19428 18662 19440
rect 19521 19431 19579 19437
rect 18656 19400 19288 19428
rect 18656 19388 18662 19400
rect 17126 19320 17132 19372
rect 17184 19320 17190 19372
rect 17678 19320 17684 19372
rect 17736 19360 17742 19372
rect 18509 19363 18567 19369
rect 18509 19360 18521 19363
rect 17736 19332 18521 19360
rect 17736 19320 17742 19332
rect 18509 19329 18521 19332
rect 18555 19329 18567 19363
rect 18509 19323 18567 19329
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19360 18751 19363
rect 18739 19332 18920 19360
rect 18739 19329 18751 19332
rect 18693 19323 18751 19329
rect 18524 19292 18552 19323
rect 18598 19292 18604 19304
rect 18524 19264 18604 19292
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 18892 19292 18920 19332
rect 18966 19320 18972 19372
rect 19024 19320 19030 19372
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19260 19369 19288 19400
rect 19521 19397 19533 19431
rect 19567 19428 19579 19431
rect 20165 19431 20223 19437
rect 20165 19428 20177 19431
rect 19567 19400 20177 19428
rect 19567 19397 19579 19400
rect 19521 19391 19579 19397
rect 20165 19397 20177 19400
rect 20211 19428 20223 19431
rect 20622 19428 20628 19440
rect 20211 19400 20628 19428
rect 20211 19397 20223 19400
rect 20165 19391 20223 19397
rect 20622 19388 20628 19400
rect 20680 19388 20686 19440
rect 22572 19428 22600 19456
rect 22572 19400 22784 19428
rect 19153 19363 19211 19369
rect 19153 19360 19165 19363
rect 19116 19332 19165 19360
rect 19116 19320 19122 19332
rect 19153 19329 19165 19332
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19329 19303 19363
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 19245 19323 19303 19329
rect 19352 19332 19441 19360
rect 19352 19304 19380 19332
rect 19429 19329 19441 19332
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19360 19671 19363
rect 19702 19360 19708 19372
rect 19659 19332 19708 19360
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 19889 19363 19947 19369
rect 19889 19360 19901 19363
rect 19867 19332 19901 19360
rect 19889 19329 19901 19332
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 19334 19292 19340 19304
rect 18892 19264 19340 19292
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 19904 19292 19932 19323
rect 19978 19320 19984 19372
rect 20036 19360 20042 19372
rect 20073 19363 20131 19369
rect 20073 19360 20085 19363
rect 20036 19332 20085 19360
rect 20036 19320 20042 19332
rect 20073 19329 20085 19332
rect 20119 19329 20131 19363
rect 20073 19323 20131 19329
rect 20254 19320 20260 19372
rect 20312 19320 20318 19372
rect 20898 19360 20904 19372
rect 20364 19332 20904 19360
rect 20364 19292 20392 19332
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 22646 19320 22652 19372
rect 22704 19320 22710 19372
rect 22756 19369 22784 19400
rect 22830 19388 22836 19440
rect 22888 19428 22894 19440
rect 23017 19431 23075 19437
rect 23017 19428 23029 19431
rect 22888 19400 23029 19428
rect 22888 19388 22894 19400
rect 23017 19397 23029 19400
rect 23063 19397 23075 19431
rect 23017 19391 23075 19397
rect 23290 19388 23296 19440
rect 23348 19428 23354 19440
rect 23477 19431 23535 19437
rect 23477 19428 23489 19431
rect 23348 19400 23489 19428
rect 23348 19388 23354 19400
rect 23477 19397 23489 19400
rect 23523 19397 23535 19431
rect 24762 19428 24768 19440
rect 23477 19391 23535 19397
rect 24412 19400 24768 19428
rect 24412 19372 24440 19400
rect 24762 19388 24768 19400
rect 24820 19428 24826 19440
rect 25409 19431 25467 19437
rect 25409 19428 25421 19431
rect 24820 19400 25421 19428
rect 24820 19388 24826 19400
rect 25409 19397 25421 19400
rect 25455 19397 25467 19431
rect 25409 19391 25467 19397
rect 22741 19363 22799 19369
rect 22741 19329 22753 19363
rect 22787 19329 22799 19363
rect 22741 19323 22799 19329
rect 22925 19363 22983 19369
rect 22925 19329 22937 19363
rect 22971 19329 22983 19363
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 22925 19323 22983 19329
rect 23124 19332 24041 19360
rect 22940 19306 22978 19323
rect 22950 19292 22978 19306
rect 23124 19292 23152 19332
rect 24029 19329 24041 19332
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 24118 19320 24124 19372
rect 24176 19320 24182 19372
rect 24394 19320 24400 19372
rect 24452 19320 24458 19372
rect 24489 19363 24547 19369
rect 24489 19329 24501 19363
rect 24535 19329 24547 19363
rect 24489 19323 24547 19329
rect 19904 19264 20392 19292
rect 22066 19264 22876 19292
rect 22950 19264 23152 19292
rect 19242 19224 19248 19236
rect 17052 19196 19248 19224
rect 14369 19187 14427 19193
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 20364 19196 20576 19224
rect 12342 19156 12348 19168
rect 9605 19128 12348 19156
rect 8849 19119 8907 19125
rect 12342 19116 12348 19128
rect 12400 19116 12406 19168
rect 12710 19116 12716 19168
rect 12768 19156 12774 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12768 19128 12817 19156
rect 12768 19116 12774 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 12805 19119 12863 19125
rect 12986 19116 12992 19168
rect 13044 19116 13050 19168
rect 13262 19116 13268 19168
rect 13320 19156 13326 19168
rect 13725 19159 13783 19165
rect 13725 19156 13737 19159
rect 13320 19128 13737 19156
rect 13320 19116 13326 19128
rect 13725 19125 13737 19128
rect 13771 19156 13783 19159
rect 16390 19156 16396 19168
rect 13771 19128 16396 19156
rect 13771 19125 13783 19128
rect 13725 19119 13783 19125
rect 16390 19116 16396 19128
rect 16448 19116 16454 19168
rect 16758 19116 16764 19168
rect 16816 19156 16822 19168
rect 20364 19156 20392 19196
rect 16816 19128 20392 19156
rect 16816 19116 16822 19128
rect 20438 19116 20444 19168
rect 20496 19116 20502 19168
rect 20548 19156 20576 19196
rect 21358 19184 21364 19236
rect 21416 19224 21422 19236
rect 22066 19224 22094 19264
rect 22848 19224 22876 19264
rect 23290 19252 23296 19304
rect 23348 19252 23354 19304
rect 23382 19252 23388 19304
rect 23440 19252 23446 19304
rect 24504 19292 24532 19323
rect 25222 19320 25228 19372
rect 25280 19320 25286 19372
rect 25516 19369 25544 19468
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 33137 19499 33195 19505
rect 33137 19465 33149 19499
rect 33183 19496 33195 19499
rect 33962 19496 33968 19508
rect 33183 19468 33968 19496
rect 33183 19465 33195 19468
rect 33137 19459 33195 19465
rect 33962 19456 33968 19468
rect 34020 19456 34026 19508
rect 27798 19388 27804 19440
rect 27856 19428 27862 19440
rect 29638 19428 29644 19440
rect 27856 19400 29644 19428
rect 27856 19388 27862 19400
rect 25501 19363 25559 19369
rect 25501 19329 25513 19363
rect 25547 19329 25559 19363
rect 25501 19323 25559 19329
rect 27890 19320 27896 19372
rect 27948 19320 27954 19372
rect 28092 19369 28120 19400
rect 29638 19388 29644 19400
rect 29696 19388 29702 19440
rect 28041 19363 28120 19369
rect 28041 19329 28053 19363
rect 28087 19332 28120 19363
rect 28169 19363 28227 19369
rect 28087 19329 28099 19332
rect 28041 19323 28099 19329
rect 28169 19329 28181 19363
rect 28215 19329 28227 19363
rect 28169 19323 28227 19329
rect 25041 19295 25099 19301
rect 25041 19292 25053 19295
rect 24504 19264 25053 19292
rect 25041 19261 25053 19264
rect 25087 19261 25099 19295
rect 28184 19292 28212 19323
rect 28258 19320 28264 19372
rect 28316 19320 28322 19372
rect 28399 19363 28457 19369
rect 28399 19329 28411 19363
rect 28445 19360 28457 19363
rect 28994 19360 29000 19372
rect 28445 19332 29000 19360
rect 28445 19329 28457 19332
rect 28399 19323 28457 19329
rect 28994 19320 29000 19332
rect 29052 19320 29058 19372
rect 32766 19320 32772 19372
rect 32824 19320 32830 19372
rect 34422 19360 34428 19372
rect 32968 19332 34428 19360
rect 32968 19304 32996 19332
rect 34422 19320 34428 19332
rect 34480 19320 34486 19372
rect 29086 19292 29092 19304
rect 28184 19264 29092 19292
rect 25041 19255 25099 19261
rect 29086 19252 29092 19264
rect 29144 19292 29150 19304
rect 29822 19292 29828 19304
rect 29144 19264 29828 19292
rect 29144 19252 29150 19264
rect 29822 19252 29828 19264
rect 29880 19252 29886 19304
rect 30190 19252 30196 19304
rect 30248 19292 30254 19304
rect 32858 19292 32864 19304
rect 30248 19264 32864 19292
rect 30248 19252 30254 19264
rect 32858 19252 32864 19264
rect 32916 19252 32922 19304
rect 32950 19252 32956 19304
rect 33008 19252 33014 19304
rect 26694 19224 26700 19236
rect 21416 19196 22094 19224
rect 22388 19196 22692 19224
rect 22848 19196 26700 19224
rect 21416 19184 21422 19196
rect 22388 19156 22416 19196
rect 22664 19165 22692 19196
rect 26694 19184 26700 19196
rect 26752 19224 26758 19236
rect 30466 19224 30472 19236
rect 26752 19196 30472 19224
rect 26752 19184 26758 19196
rect 30466 19184 30472 19196
rect 30524 19184 30530 19236
rect 20548 19128 22416 19156
rect 22649 19159 22707 19165
rect 22649 19125 22661 19159
rect 22695 19125 22707 19159
rect 22649 19119 22707 19125
rect 24213 19159 24271 19165
rect 24213 19125 24225 19159
rect 24259 19156 24271 19159
rect 24302 19156 24308 19168
rect 24259 19128 24308 19156
rect 24259 19125 24271 19128
rect 24213 19119 24271 19125
rect 24302 19116 24308 19128
rect 24360 19116 24366 19168
rect 24394 19116 24400 19168
rect 24452 19156 24458 19168
rect 25774 19156 25780 19168
rect 24452 19128 25780 19156
rect 24452 19116 24458 19128
rect 25774 19116 25780 19128
rect 25832 19116 25838 19168
rect 27982 19116 27988 19168
rect 28040 19156 28046 19168
rect 28166 19156 28172 19168
rect 28040 19128 28172 19156
rect 28040 19116 28046 19128
rect 28166 19116 28172 19128
rect 28224 19116 28230 19168
rect 28534 19116 28540 19168
rect 28592 19116 28598 19168
rect 30006 19116 30012 19168
rect 30064 19156 30070 19168
rect 30558 19156 30564 19168
rect 30064 19128 30564 19156
rect 30064 19116 30070 19128
rect 30558 19116 30564 19128
rect 30616 19156 30622 19168
rect 32769 19159 32827 19165
rect 32769 19156 32781 19159
rect 30616 19128 32781 19156
rect 30616 19116 30622 19128
rect 32769 19125 32781 19128
rect 32815 19125 32827 19159
rect 32769 19119 32827 19125
rect 1104 19066 36432 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 36432 19066
rect 1104 18992 36432 19014
rect 3145 18955 3203 18961
rect 3145 18921 3157 18955
rect 3191 18952 3203 18955
rect 3510 18952 3516 18964
rect 3191 18924 3516 18952
rect 3191 18921 3203 18924
rect 3145 18915 3203 18921
rect 3510 18912 3516 18924
rect 3568 18952 3574 18964
rect 3878 18952 3884 18964
rect 3568 18924 3884 18952
rect 3568 18912 3574 18924
rect 3878 18912 3884 18924
rect 3936 18912 3942 18964
rect 4893 18955 4951 18961
rect 4893 18921 4905 18955
rect 4939 18952 4951 18955
rect 5442 18952 5448 18964
rect 4939 18924 5448 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 6730 18912 6736 18964
rect 6788 18912 6794 18964
rect 8754 18952 8760 18964
rect 6840 18924 8760 18952
rect 4614 18844 4620 18896
rect 4672 18844 4678 18896
rect 6638 18844 6644 18896
rect 6696 18884 6702 18896
rect 6840 18884 6868 18924
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 9398 18912 9404 18964
rect 9456 18952 9462 18964
rect 9858 18952 9864 18964
rect 9456 18924 9864 18952
rect 9456 18912 9462 18924
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10686 18912 10692 18964
rect 10744 18952 10750 18964
rect 10744 18924 11652 18952
rect 10744 18912 10750 18924
rect 6696 18856 6868 18884
rect 6696 18844 6702 18856
rect 6914 18844 6920 18896
rect 6972 18884 6978 18896
rect 6972 18856 8524 18884
rect 6972 18844 6978 18856
rect 4632 18816 4660 18844
rect 4356 18788 4660 18816
rect 1394 18708 1400 18760
rect 1452 18708 1458 18760
rect 2774 18708 2780 18760
rect 2832 18708 2838 18760
rect 4356 18757 4384 18788
rect 4982 18776 4988 18828
rect 5040 18816 5046 18828
rect 5442 18816 5448 18828
rect 5040 18788 5448 18816
rect 5040 18776 5046 18788
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 7006 18776 7012 18828
rect 7064 18816 7070 18828
rect 7285 18819 7343 18825
rect 7285 18816 7297 18819
rect 7064 18788 7297 18816
rect 7064 18776 7070 18788
rect 7285 18785 7297 18788
rect 7331 18816 7343 18819
rect 8297 18819 8355 18825
rect 7331 18788 8248 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 4341 18751 4399 18757
rect 4341 18717 4353 18751
rect 4387 18717 4399 18751
rect 4341 18711 4399 18717
rect 4430 18708 4436 18760
rect 4488 18708 4494 18760
rect 4617 18751 4675 18757
rect 4617 18717 4629 18751
rect 4663 18717 4675 18751
rect 4617 18711 4675 18717
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4890 18748 4896 18760
rect 4755 18720 4896 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 1670 18640 1676 18692
rect 1728 18640 1734 18692
rect 4632 18680 4660 18711
rect 4890 18708 4896 18720
rect 4948 18748 4954 18760
rect 7193 18751 7251 18757
rect 4948 18720 7052 18748
rect 4948 18708 4954 18720
rect 5350 18680 5356 18692
rect 4632 18652 5356 18680
rect 5350 18640 5356 18652
rect 5408 18640 5414 18692
rect 7024 18612 7052 18720
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 8018 18748 8024 18760
rect 7239 18720 8024 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 8018 18708 8024 18720
rect 8076 18708 8082 18760
rect 7101 18683 7159 18689
rect 7101 18649 7113 18683
rect 7147 18680 7159 18683
rect 7653 18683 7711 18689
rect 7653 18680 7665 18683
rect 7147 18652 7665 18680
rect 7147 18649 7159 18652
rect 7101 18643 7159 18649
rect 7653 18649 7665 18652
rect 7699 18649 7711 18683
rect 8220 18680 8248 18788
rect 8297 18785 8309 18819
rect 8343 18816 8355 18819
rect 8386 18816 8392 18828
rect 8343 18788 8392 18816
rect 8343 18785 8355 18788
rect 8297 18779 8355 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 8496 18816 8524 18856
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 8496 18788 8953 18816
rect 8941 18785 8953 18788
rect 8987 18785 8999 18819
rect 8941 18779 8999 18785
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 9582 18816 9588 18828
rect 9272 18788 9588 18816
rect 9272 18776 9278 18788
rect 9582 18776 9588 18788
rect 9640 18776 9646 18828
rect 10686 18776 10692 18828
rect 10744 18816 10750 18828
rect 11146 18816 11152 18828
rect 10744 18788 11152 18816
rect 10744 18776 10750 18788
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 11425 18819 11483 18825
rect 11425 18785 11437 18819
rect 11471 18816 11483 18819
rect 11624 18816 11652 18924
rect 12066 18912 12072 18964
rect 12124 18952 12130 18964
rect 12124 18924 13584 18952
rect 12124 18912 12130 18924
rect 12434 18884 12440 18896
rect 11471 18788 11652 18816
rect 11716 18856 12440 18884
rect 11471 18785 11483 18788
rect 11425 18779 11483 18785
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18748 8631 18751
rect 8754 18748 8760 18760
rect 8619 18720 8760 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11716 18757 11744 18856
rect 12434 18844 12440 18856
rect 12492 18884 12498 18896
rect 12492 18856 12572 18884
rect 12492 18844 12498 18856
rect 12544 18816 12572 18856
rect 12710 18844 12716 18896
rect 12768 18884 12774 18896
rect 13265 18887 13323 18893
rect 13265 18884 13277 18887
rect 12768 18856 13277 18884
rect 12768 18844 12774 18856
rect 13265 18853 13277 18856
rect 13311 18853 13323 18887
rect 13265 18847 13323 18853
rect 12544 18788 13308 18816
rect 11701 18751 11759 18757
rect 11701 18748 11713 18751
rect 11112 18720 11713 18748
rect 11112 18708 11118 18720
rect 11701 18717 11713 18720
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 11790 18708 11796 18760
rect 11848 18708 11854 18760
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 11940 18720 11989 18748
rect 11940 18708 11946 18720
rect 11977 18717 11989 18720
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 12066 18708 12072 18760
rect 12124 18708 12130 18760
rect 12345 18751 12403 18757
rect 12345 18748 12357 18751
rect 12175 18720 12357 18748
rect 8220 18652 9168 18680
rect 7653 18643 7711 18649
rect 8386 18612 8392 18624
rect 7024 18584 8392 18612
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 8665 18615 8723 18621
rect 8665 18581 8677 18615
rect 8711 18612 8723 18615
rect 8846 18612 8852 18624
rect 8711 18584 8852 18612
rect 8711 18581 8723 18584
rect 8665 18575 8723 18581
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 9140 18612 9168 18652
rect 9214 18640 9220 18692
rect 9272 18640 9278 18692
rect 9766 18640 9772 18692
rect 9824 18640 9830 18692
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 10781 18683 10839 18689
rect 10781 18680 10793 18683
rect 10560 18652 10793 18680
rect 10560 18640 10566 18652
rect 10781 18649 10793 18652
rect 10827 18649 10839 18683
rect 10781 18643 10839 18649
rect 11238 18640 11244 18692
rect 11296 18680 11302 18692
rect 12175 18680 12203 18720
rect 12345 18717 12357 18720
rect 12391 18717 12403 18751
rect 12345 18711 12403 18717
rect 12529 18751 12587 18757
rect 12529 18717 12541 18751
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 11296 18652 12203 18680
rect 11296 18640 11302 18652
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 12544 18680 12572 18711
rect 12802 18708 12808 18760
rect 12860 18708 12866 18760
rect 13078 18708 13084 18760
rect 13136 18708 13142 18760
rect 13280 18757 13308 18788
rect 13265 18751 13323 18757
rect 13265 18717 13277 18751
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 13446 18708 13452 18760
rect 13504 18708 13510 18760
rect 13556 18757 13584 18924
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 14090 18952 14096 18964
rect 13688 18924 14096 18952
rect 13688 18912 13694 18924
rect 14090 18912 14096 18924
rect 14148 18952 14154 18964
rect 15378 18952 15384 18964
rect 14148 18924 15384 18952
rect 14148 18912 14154 18924
rect 15378 18912 15384 18924
rect 15436 18912 15442 18964
rect 16758 18912 16764 18964
rect 16816 18952 16822 18964
rect 17037 18955 17095 18961
rect 17037 18952 17049 18955
rect 16816 18924 17049 18952
rect 16816 18912 16822 18924
rect 17037 18921 17049 18924
rect 17083 18921 17095 18955
rect 17037 18915 17095 18921
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 21729 18955 21787 18961
rect 21729 18952 21741 18955
rect 20956 18924 21741 18952
rect 20956 18912 20962 18924
rect 21729 18921 21741 18924
rect 21775 18952 21787 18955
rect 21818 18952 21824 18964
rect 21775 18924 21824 18952
rect 21775 18921 21787 18924
rect 21729 18915 21787 18921
rect 21818 18912 21824 18924
rect 21876 18912 21882 18964
rect 23106 18912 23112 18964
rect 23164 18912 23170 18964
rect 24302 18912 24308 18964
rect 24360 18952 24366 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 24360 18924 24409 18952
rect 24360 18912 24366 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24397 18915 24455 18921
rect 26513 18955 26571 18961
rect 26513 18921 26525 18955
rect 26559 18952 26571 18955
rect 28718 18952 28724 18964
rect 26559 18924 28724 18952
rect 26559 18921 26571 18924
rect 26513 18915 26571 18921
rect 28718 18912 28724 18924
rect 28776 18952 28782 18964
rect 29178 18952 29184 18964
rect 28776 18924 29184 18952
rect 28776 18912 28782 18924
rect 29178 18912 29184 18924
rect 29236 18912 29242 18964
rect 30190 18912 30196 18964
rect 30248 18912 30254 18964
rect 30650 18912 30656 18964
rect 30708 18912 30714 18964
rect 33686 18912 33692 18964
rect 33744 18952 33750 18964
rect 34701 18955 34759 18961
rect 34701 18952 34713 18955
rect 33744 18924 34713 18952
rect 33744 18912 33750 18924
rect 34701 18921 34713 18924
rect 34747 18921 34759 18955
rect 34701 18915 34759 18921
rect 16666 18884 16672 18896
rect 14660 18856 16672 18884
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18717 13599 18751
rect 13541 18711 13599 18717
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18748 14519 18751
rect 14660 18748 14688 18856
rect 16666 18844 16672 18856
rect 16724 18844 16730 18896
rect 18141 18887 18199 18893
rect 18141 18853 18153 18887
rect 18187 18884 18199 18887
rect 26145 18887 26203 18893
rect 26145 18884 26157 18887
rect 18187 18856 26157 18884
rect 18187 18853 18199 18856
rect 18141 18847 18199 18853
rect 26145 18853 26157 18856
rect 26191 18853 26203 18887
rect 28166 18884 28172 18896
rect 26145 18847 26203 18853
rect 27816 18856 28172 18884
rect 15930 18816 15936 18828
rect 14752 18788 15936 18816
rect 14752 18757 14780 18788
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 16209 18819 16267 18825
rect 16209 18785 16221 18819
rect 16255 18816 16267 18819
rect 16574 18816 16580 18828
rect 16255 18788 16580 18816
rect 16255 18785 16267 18788
rect 16209 18779 16267 18785
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 21266 18776 21272 18828
rect 21324 18816 21330 18828
rect 22002 18816 22008 18828
rect 21324 18788 22008 18816
rect 21324 18776 21330 18788
rect 22002 18776 22008 18788
rect 22060 18816 22066 18828
rect 22833 18819 22891 18825
rect 22833 18816 22845 18819
rect 22060 18788 22845 18816
rect 22060 18776 22066 18788
rect 22833 18785 22845 18788
rect 22879 18785 22891 18819
rect 22833 18779 22891 18785
rect 23216 18788 26004 18816
rect 14507 18720 14688 18748
rect 14737 18751 14795 18757
rect 14507 18717 14519 18720
rect 14461 18711 14519 18717
rect 14737 18717 14749 18751
rect 14783 18717 14795 18751
rect 14737 18711 14795 18717
rect 12308 18652 12572 18680
rect 12713 18683 12771 18689
rect 12308 18640 12314 18652
rect 12713 18649 12725 18683
rect 12759 18680 12771 18683
rect 13170 18680 13176 18692
rect 12759 18652 13176 18680
rect 12759 18649 12771 18652
rect 12713 18643 12771 18649
rect 13170 18640 13176 18652
rect 13228 18640 13234 18692
rect 9858 18612 9864 18624
rect 9140 18584 9864 18612
rect 9858 18572 9864 18584
rect 9916 18612 9922 18624
rect 10870 18612 10876 18624
rect 9916 18584 10876 18612
rect 9916 18572 9922 18584
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 12342 18572 12348 18624
rect 12400 18612 12406 18624
rect 12897 18615 12955 18621
rect 12897 18612 12909 18615
rect 12400 18584 12909 18612
rect 12400 18572 12406 18584
rect 12897 18581 12909 18584
rect 12943 18581 12955 18615
rect 13556 18612 13584 18711
rect 15746 18708 15752 18760
rect 15804 18708 15810 18760
rect 16114 18708 16120 18760
rect 16172 18708 16178 18760
rect 16666 18708 16672 18760
rect 16724 18748 16730 18760
rect 17034 18748 17040 18760
rect 16724 18720 17040 18748
rect 16724 18708 16730 18720
rect 17034 18708 17040 18720
rect 17092 18708 17098 18760
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 17773 18751 17831 18757
rect 17773 18748 17785 18751
rect 17451 18720 17785 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 17773 18717 17785 18720
rect 17819 18717 17831 18751
rect 17773 18711 17831 18717
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18748 18107 18751
rect 18138 18748 18144 18760
rect 18095 18720 18144 18748
rect 18095 18717 18107 18720
rect 18049 18711 18107 18717
rect 14182 18640 14188 18692
rect 14240 18680 14246 18692
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 14240 18652 14381 18680
rect 14240 18640 14246 18652
rect 14369 18649 14381 18652
rect 14415 18680 14427 18683
rect 14550 18680 14556 18692
rect 14415 18652 14556 18680
rect 14415 18649 14427 18652
rect 14369 18643 14427 18649
rect 14550 18640 14556 18652
rect 14608 18640 14614 18692
rect 17678 18640 17684 18692
rect 17736 18680 17742 18692
rect 17972 18680 18000 18711
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 18230 18708 18236 18760
rect 18288 18708 18294 18760
rect 21542 18708 21548 18760
rect 21600 18708 21606 18760
rect 21910 18708 21916 18760
rect 21968 18708 21974 18760
rect 22094 18708 22100 18760
rect 22152 18708 22158 18760
rect 23216 18748 23244 18788
rect 22756 18720 23244 18748
rect 17736 18652 18000 18680
rect 17736 18640 17742 18652
rect 18598 18640 18604 18692
rect 18656 18680 18662 18692
rect 22756 18680 22784 18720
rect 23290 18708 23296 18760
rect 23348 18708 23354 18760
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18717 23443 18751
rect 23385 18711 23443 18717
rect 18656 18652 22784 18680
rect 23400 18680 23428 18711
rect 23474 18708 23480 18760
rect 23532 18708 23538 18760
rect 23569 18751 23627 18757
rect 23569 18717 23581 18751
rect 23615 18748 23627 18751
rect 23937 18751 23995 18757
rect 23615 18720 23888 18748
rect 23615 18717 23627 18720
rect 23569 18711 23627 18717
rect 23658 18680 23664 18692
rect 23400 18652 23664 18680
rect 18656 18640 18662 18652
rect 23658 18640 23664 18652
rect 23716 18680 23722 18692
rect 23753 18683 23811 18689
rect 23753 18680 23765 18683
rect 23716 18652 23765 18680
rect 23716 18640 23722 18652
rect 23753 18649 23765 18652
rect 23799 18649 23811 18683
rect 23753 18643 23811 18649
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 13556 18584 15577 18612
rect 12897 18575 12955 18581
rect 15565 18581 15577 18584
rect 15611 18581 15623 18615
rect 15565 18575 15623 18581
rect 15749 18615 15807 18621
rect 15749 18581 15761 18615
rect 15795 18612 15807 18615
rect 16206 18612 16212 18624
rect 15795 18584 16212 18612
rect 15795 18581 15807 18584
rect 15749 18575 15807 18581
rect 16206 18572 16212 18584
rect 16264 18572 16270 18624
rect 16850 18572 16856 18624
rect 16908 18572 16914 18624
rect 21266 18572 21272 18624
rect 21324 18612 21330 18624
rect 21361 18615 21419 18621
rect 21361 18612 21373 18615
rect 21324 18584 21373 18612
rect 21324 18572 21330 18584
rect 21361 18581 21373 18584
rect 21407 18581 21419 18615
rect 21361 18575 21419 18581
rect 23290 18572 23296 18624
rect 23348 18612 23354 18624
rect 23860 18612 23888 18720
rect 23937 18717 23949 18751
rect 23983 18748 23995 18751
rect 24302 18748 24308 18760
rect 23983 18720 24308 18748
rect 23983 18717 23995 18720
rect 23937 18711 23995 18717
rect 24302 18708 24308 18720
rect 24360 18708 24366 18760
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24121 18683 24179 18689
rect 24121 18649 24133 18683
rect 24167 18680 24179 18683
rect 24210 18680 24216 18692
rect 24167 18652 24216 18680
rect 24167 18649 24179 18652
rect 24121 18643 24179 18649
rect 24210 18640 24216 18652
rect 24268 18640 24274 18692
rect 24596 18680 24624 18711
rect 24670 18708 24676 18760
rect 24728 18708 24734 18760
rect 24872 18757 24900 18788
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 24857 18751 24915 18757
rect 24857 18717 24869 18751
rect 24903 18717 24915 18751
rect 24857 18711 24915 18717
rect 24780 18680 24808 18711
rect 25222 18708 25228 18760
rect 25280 18748 25286 18760
rect 25685 18751 25743 18757
rect 25685 18748 25697 18751
rect 25280 18720 25697 18748
rect 25280 18708 25286 18720
rect 25685 18717 25697 18720
rect 25731 18717 25743 18751
rect 25685 18711 25743 18717
rect 25777 18751 25835 18757
rect 25777 18717 25789 18751
rect 25823 18717 25835 18751
rect 25777 18711 25835 18717
rect 25590 18680 25596 18692
rect 24596 18652 24716 18680
rect 24780 18652 25596 18680
rect 23348 18584 23888 18612
rect 24688 18612 24716 18652
rect 25590 18640 25596 18652
rect 25648 18640 25654 18692
rect 25792 18680 25820 18711
rect 25866 18708 25872 18760
rect 25924 18708 25930 18760
rect 25976 18757 26004 18788
rect 26050 18776 26056 18828
rect 26108 18816 26114 18828
rect 26605 18819 26663 18825
rect 26605 18816 26617 18819
rect 26108 18788 26617 18816
rect 26108 18776 26114 18788
rect 26605 18785 26617 18788
rect 26651 18785 26663 18819
rect 26605 18779 26663 18785
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18748 26019 18751
rect 26329 18751 26387 18757
rect 26329 18748 26341 18751
rect 26007 18720 26341 18748
rect 26007 18717 26019 18720
rect 25961 18711 26019 18717
rect 26329 18717 26341 18720
rect 26375 18717 26387 18751
rect 26329 18711 26387 18717
rect 26694 18708 26700 18760
rect 26752 18708 26758 18760
rect 26881 18751 26939 18757
rect 26881 18717 26893 18751
rect 26927 18748 26939 18751
rect 27062 18748 27068 18760
rect 26927 18720 27068 18748
rect 26927 18717 26939 18720
rect 26881 18711 26939 18717
rect 27062 18708 27068 18720
rect 27120 18708 27126 18760
rect 27522 18708 27528 18760
rect 27580 18708 27586 18760
rect 27614 18708 27620 18760
rect 27672 18708 27678 18760
rect 27816 18757 27844 18856
rect 28166 18844 28172 18856
rect 28224 18884 28230 18896
rect 28902 18884 28908 18896
rect 28224 18856 28908 18884
rect 28224 18844 28230 18856
rect 28902 18844 28908 18856
rect 28960 18844 28966 18896
rect 33594 18884 33600 18896
rect 31726 18856 33600 18884
rect 28920 18816 28948 18844
rect 28920 18788 30972 18816
rect 27801 18751 27859 18757
rect 27801 18717 27813 18751
rect 27847 18717 27859 18751
rect 27801 18711 27859 18717
rect 27982 18708 27988 18760
rect 28040 18757 28046 18760
rect 28040 18748 28048 18757
rect 28040 18720 28085 18748
rect 28040 18711 28048 18720
rect 28040 18708 28046 18711
rect 29546 18708 29552 18760
rect 29604 18708 29610 18760
rect 29638 18708 29644 18760
rect 29696 18748 29702 18760
rect 29696 18720 29741 18748
rect 29696 18708 29702 18720
rect 29822 18708 29828 18760
rect 29880 18708 29886 18760
rect 30055 18751 30113 18757
rect 30055 18717 30067 18751
rect 30101 18748 30113 18751
rect 30742 18748 30748 18760
rect 30101 18720 30748 18748
rect 30101 18717 30113 18720
rect 30055 18711 30113 18717
rect 30742 18708 30748 18720
rect 30800 18748 30806 18760
rect 30837 18751 30895 18757
rect 30837 18748 30849 18751
rect 30800 18720 30849 18748
rect 30800 18708 30806 18720
rect 30837 18717 30849 18720
rect 30883 18717 30895 18751
rect 30944 18748 30972 18788
rect 31205 18751 31263 18757
rect 30944 18720 31064 18748
rect 30837 18711 30895 18717
rect 26050 18680 26056 18692
rect 25792 18652 26056 18680
rect 26050 18640 26056 18652
rect 26108 18640 26114 18692
rect 27430 18640 27436 18692
rect 27488 18680 27494 18692
rect 27893 18683 27951 18689
rect 27893 18680 27905 18683
rect 27488 18652 27905 18680
rect 27488 18640 27494 18652
rect 27893 18649 27905 18652
rect 27939 18649 27951 18683
rect 28258 18680 28264 18692
rect 27893 18643 27951 18649
rect 28092 18652 28264 18680
rect 24946 18612 24952 18624
rect 24688 18584 24952 18612
rect 23348 18572 23354 18584
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 25498 18572 25504 18624
rect 25556 18572 25562 18624
rect 25866 18572 25872 18624
rect 25924 18612 25930 18624
rect 27065 18615 27123 18621
rect 27065 18612 27077 18615
rect 25924 18584 27077 18612
rect 25924 18572 25930 18584
rect 27065 18581 27077 18584
rect 27111 18612 27123 18615
rect 28092 18612 28120 18652
rect 28258 18640 28264 18652
rect 28316 18680 28322 18692
rect 29917 18683 29975 18689
rect 28316 18652 29776 18680
rect 28316 18640 28322 18652
rect 27111 18584 28120 18612
rect 28169 18615 28227 18621
rect 27111 18581 27123 18584
rect 27065 18575 27123 18581
rect 28169 18581 28181 18615
rect 28215 18612 28227 18615
rect 28902 18612 28908 18624
rect 28215 18584 28908 18612
rect 28215 18581 28227 18584
rect 28169 18575 28227 18581
rect 28902 18572 28908 18584
rect 28960 18572 28966 18624
rect 29748 18612 29776 18652
rect 29917 18649 29929 18683
rect 29963 18649 29975 18683
rect 29917 18643 29975 18649
rect 29932 18612 29960 18643
rect 30466 18640 30472 18692
rect 30524 18680 30530 18692
rect 31036 18689 31064 18720
rect 31205 18717 31217 18751
rect 31251 18748 31263 18751
rect 31726 18748 31754 18856
rect 33594 18844 33600 18856
rect 33652 18844 33658 18896
rect 32858 18776 32864 18828
rect 32916 18816 32922 18828
rect 34793 18819 34851 18825
rect 34793 18816 34805 18819
rect 32916 18788 34805 18816
rect 32916 18776 32922 18788
rect 34793 18785 34805 18788
rect 34839 18785 34851 18819
rect 34793 18779 34851 18785
rect 31251 18720 31754 18748
rect 31251 18717 31263 18720
rect 31205 18711 31263 18717
rect 33226 18708 33232 18760
rect 33284 18748 33290 18760
rect 34701 18751 34759 18757
rect 34701 18748 34713 18751
rect 33284 18720 34713 18748
rect 33284 18708 33290 18720
rect 34701 18717 34713 18720
rect 34747 18717 34759 18751
rect 34701 18711 34759 18717
rect 34977 18751 35035 18757
rect 34977 18717 34989 18751
rect 35023 18748 35035 18751
rect 35342 18748 35348 18760
rect 35023 18720 35348 18748
rect 35023 18717 35035 18720
rect 34977 18711 35035 18717
rect 35342 18708 35348 18720
rect 35400 18708 35406 18760
rect 30929 18683 30987 18689
rect 30929 18680 30941 18683
rect 30524 18652 30941 18680
rect 30524 18640 30530 18652
rect 30929 18649 30941 18652
rect 30975 18649 30987 18683
rect 30929 18643 30987 18649
rect 31021 18683 31079 18689
rect 31021 18649 31033 18683
rect 31067 18680 31079 18683
rect 33686 18680 33692 18692
rect 31067 18652 33692 18680
rect 31067 18649 31079 18652
rect 31021 18643 31079 18649
rect 33686 18640 33692 18652
rect 33744 18640 33750 18692
rect 29748 18584 29960 18612
rect 30098 18572 30104 18624
rect 30156 18612 30162 18624
rect 33318 18612 33324 18624
rect 30156 18584 33324 18612
rect 30156 18572 30162 18584
rect 33318 18572 33324 18584
rect 33376 18572 33382 18624
rect 35161 18615 35219 18621
rect 35161 18581 35173 18615
rect 35207 18612 35219 18615
rect 35342 18612 35348 18624
rect 35207 18584 35348 18612
rect 35207 18581 35219 18584
rect 35161 18575 35219 18581
rect 35342 18572 35348 18584
rect 35400 18572 35406 18624
rect 1104 18522 36432 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 36432 18522
rect 1104 18448 36432 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 2041 18411 2099 18417
rect 2041 18408 2053 18411
rect 1728 18380 2053 18408
rect 1728 18368 1734 18380
rect 2041 18377 2053 18380
rect 2087 18377 2099 18411
rect 2041 18371 2099 18377
rect 5442 18368 5448 18420
rect 5500 18408 5506 18420
rect 7558 18408 7564 18420
rect 5500 18380 7564 18408
rect 5500 18368 5506 18380
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18272 2467 18275
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 2455 18244 2881 18272
rect 2455 18241 2467 18244
rect 2409 18235 2467 18241
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 3510 18232 3516 18284
rect 3568 18232 3574 18284
rect 6748 18281 6776 18380
rect 7558 18368 7564 18380
rect 7616 18368 7622 18420
rect 7742 18368 7748 18420
rect 7800 18368 7806 18420
rect 7834 18368 7840 18420
rect 7892 18368 7898 18420
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 8478 18408 8484 18420
rect 8251 18380 8484 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 9033 18411 9091 18417
rect 9033 18377 9045 18411
rect 9079 18408 9091 18411
rect 9214 18408 9220 18420
rect 9079 18380 9220 18408
rect 9079 18377 9091 18380
rect 9033 18371 9091 18377
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 9401 18411 9459 18417
rect 9401 18377 9413 18411
rect 9447 18408 9459 18411
rect 10502 18408 10508 18420
rect 9447 18380 10508 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 11241 18411 11299 18417
rect 10612 18380 10916 18408
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18340 6883 18343
rect 7098 18340 7104 18352
rect 6871 18312 7104 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 8312 18312 8800 18340
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18272 7067 18275
rect 8312 18272 8340 18312
rect 7055 18244 8340 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 2498 18164 2504 18216
rect 2556 18164 2562 18216
rect 2590 18164 2596 18216
rect 2648 18164 2654 18216
rect 5718 18164 5724 18216
rect 5776 18204 5782 18216
rect 7024 18204 7052 18235
rect 8386 18232 8392 18284
rect 8444 18232 8450 18284
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18272 8539 18275
rect 8570 18272 8576 18284
rect 8527 18244 8576 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 8662 18232 8668 18284
rect 8720 18232 8726 18284
rect 8772 18281 8800 18312
rect 9490 18300 9496 18352
rect 9548 18300 9554 18352
rect 10042 18300 10048 18352
rect 10100 18300 10106 18352
rect 10134 18300 10140 18352
rect 10192 18340 10198 18352
rect 10612 18349 10640 18380
rect 10229 18343 10287 18349
rect 10229 18340 10241 18343
rect 10192 18312 10241 18340
rect 10192 18300 10198 18312
rect 10229 18309 10241 18312
rect 10275 18309 10287 18343
rect 10229 18303 10287 18309
rect 10597 18343 10655 18349
rect 10597 18309 10609 18343
rect 10643 18309 10655 18343
rect 10597 18303 10655 18309
rect 10781 18343 10839 18349
rect 10781 18309 10793 18343
rect 10827 18309 10839 18343
rect 10888 18340 10916 18380
rect 11241 18377 11253 18411
rect 11287 18408 11299 18411
rect 11882 18408 11888 18420
rect 11287 18380 11888 18408
rect 11287 18377 11299 18380
rect 11241 18371 11299 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12802 18408 12808 18420
rect 12406 18380 12808 18408
rect 11422 18340 11428 18352
rect 10888 18312 11428 18340
rect 10781 18303 10839 18309
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18272 8815 18275
rect 8938 18272 8944 18284
rect 8803 18244 8944 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10686 18272 10692 18284
rect 10367 18244 10692 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 5776 18176 7052 18204
rect 8021 18207 8079 18213
rect 5776 18164 5782 18176
rect 8021 18173 8033 18207
rect 8067 18204 8079 18207
rect 8846 18204 8852 18216
rect 8067 18176 8852 18204
rect 8067 18173 8079 18176
rect 8021 18167 8079 18173
rect 8846 18164 8852 18176
rect 8904 18164 8910 18216
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 9858 18204 9864 18216
rect 9723 18176 9864 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10226 18164 10232 18216
rect 10284 18204 10290 18216
rect 10336 18204 10364 18235
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 10796 18272 10824 18303
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 10796 18244 10916 18272
rect 10888 18213 10916 18244
rect 10962 18232 10968 18284
rect 11020 18272 11026 18284
rect 11057 18275 11115 18281
rect 11057 18272 11069 18275
rect 11020 18244 11069 18272
rect 11020 18232 11026 18244
rect 11057 18241 11069 18244
rect 11103 18241 11115 18275
rect 11057 18235 11115 18241
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 11882 18272 11888 18284
rect 11379 18244 11888 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 11882 18232 11888 18244
rect 11940 18272 11946 18284
rect 12066 18272 12072 18284
rect 11940 18244 12072 18272
rect 11940 18232 11946 18244
rect 12066 18232 12072 18244
rect 12124 18232 12130 18284
rect 12158 18232 12164 18284
rect 12216 18272 12222 18284
rect 12406 18272 12434 18380
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 13078 18368 13084 18420
rect 13136 18408 13142 18420
rect 13265 18411 13323 18417
rect 13265 18408 13277 18411
rect 13136 18380 13277 18408
rect 13136 18368 13142 18380
rect 13265 18377 13277 18380
rect 13311 18377 13323 18411
rect 13265 18371 13323 18377
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 15746 18408 15752 18420
rect 13872 18380 15752 18408
rect 13872 18368 13878 18380
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 20809 18411 20867 18417
rect 20809 18377 20821 18411
rect 20855 18408 20867 18411
rect 21450 18408 21456 18420
rect 20855 18380 21456 18408
rect 20855 18377 20867 18380
rect 20809 18371 20867 18377
rect 21450 18368 21456 18380
rect 21508 18408 21514 18420
rect 21508 18380 22232 18408
rect 21508 18368 21514 18380
rect 13096 18340 13124 18368
rect 16850 18340 16856 18352
rect 12544 18312 13124 18340
rect 13188 18312 16856 18340
rect 12544 18281 12572 18312
rect 12216 18244 12434 18272
rect 12529 18275 12587 18281
rect 12216 18232 12222 18244
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 12710 18232 12716 18284
rect 12768 18232 12774 18284
rect 12986 18232 12992 18284
rect 13044 18272 13050 18284
rect 13188 18272 13216 18312
rect 13464 18281 13492 18312
rect 16850 18300 16856 18312
rect 16908 18300 16914 18352
rect 20993 18343 21051 18349
rect 20993 18309 21005 18343
rect 21039 18340 21051 18343
rect 21039 18312 21312 18340
rect 21039 18309 21051 18312
rect 20993 18303 21051 18309
rect 21284 18284 21312 18312
rect 22002 18300 22008 18352
rect 22060 18340 22066 18352
rect 22204 18340 22232 18380
rect 23014 18368 23020 18420
rect 23072 18368 23078 18420
rect 24305 18411 24363 18417
rect 24305 18377 24317 18411
rect 24351 18408 24363 18411
rect 24578 18408 24584 18420
rect 24351 18380 24584 18408
rect 24351 18377 24363 18380
rect 24305 18371 24363 18377
rect 24578 18368 24584 18380
rect 24636 18368 24642 18420
rect 25774 18368 25780 18420
rect 25832 18408 25838 18420
rect 26053 18411 26111 18417
rect 26053 18408 26065 18411
rect 25832 18380 26065 18408
rect 25832 18368 25838 18380
rect 26053 18377 26065 18380
rect 26099 18408 26111 18411
rect 26694 18408 26700 18420
rect 26099 18380 26700 18408
rect 26099 18377 26111 18380
rect 26053 18371 26111 18377
rect 26694 18368 26700 18380
rect 26752 18368 26758 18420
rect 27614 18368 27620 18420
rect 27672 18408 27678 18420
rect 27801 18411 27859 18417
rect 27801 18408 27813 18411
rect 27672 18380 27813 18408
rect 27672 18368 27678 18380
rect 27801 18377 27813 18380
rect 27847 18408 27859 18411
rect 27890 18408 27896 18420
rect 27847 18380 27896 18408
rect 27847 18377 27859 18380
rect 27801 18371 27859 18377
rect 27890 18368 27896 18380
rect 27948 18368 27954 18420
rect 30742 18368 30748 18420
rect 30800 18408 30806 18420
rect 31570 18408 31576 18420
rect 30800 18380 31576 18408
rect 30800 18368 30806 18380
rect 31570 18368 31576 18380
rect 31628 18368 31634 18420
rect 31846 18368 31852 18420
rect 31904 18408 31910 18420
rect 34057 18411 34115 18417
rect 31904 18380 33916 18408
rect 31904 18368 31910 18380
rect 23169 18343 23227 18349
rect 23169 18340 23181 18343
rect 22060 18300 22094 18340
rect 22204 18312 23181 18340
rect 23169 18309 23181 18312
rect 23215 18309 23227 18343
rect 23169 18303 23227 18309
rect 23385 18343 23443 18349
rect 23385 18309 23397 18343
rect 23431 18309 23443 18343
rect 23385 18303 23443 18309
rect 13044 18244 13216 18272
rect 13265 18275 13323 18281
rect 13044 18232 13050 18244
rect 13265 18241 13277 18275
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18241 13507 18275
rect 13449 18235 13507 18241
rect 10284 18176 10364 18204
rect 10873 18207 10931 18213
rect 10284 18164 10290 18176
rect 10873 18173 10885 18207
rect 10919 18204 10931 18207
rect 10919 18176 11008 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 7193 18139 7251 18145
rect 7193 18105 7205 18139
rect 7239 18136 7251 18139
rect 9122 18136 9128 18148
rect 7239 18108 9128 18136
rect 7239 18105 7251 18108
rect 7193 18099 7251 18105
rect 9122 18096 9128 18108
rect 9180 18096 9186 18148
rect 9692 18108 10640 18136
rect 9692 18080 9720 18108
rect 7374 18028 7380 18080
rect 7432 18028 7438 18080
rect 8386 18028 8392 18080
rect 8444 18068 8450 18080
rect 9214 18068 9220 18080
rect 8444 18040 9220 18068
rect 8444 18028 8450 18040
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 9674 18028 9680 18080
rect 9732 18028 9738 18080
rect 9861 18071 9919 18077
rect 9861 18037 9873 18071
rect 9907 18068 9919 18071
rect 10042 18068 10048 18080
rect 9907 18040 10048 18068
rect 9907 18037 9919 18040
rect 9861 18031 9919 18037
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 10612 18077 10640 18108
rect 10597 18071 10655 18077
rect 10597 18037 10609 18071
rect 10643 18068 10655 18071
rect 10686 18068 10692 18080
rect 10643 18040 10692 18068
rect 10643 18037 10655 18040
rect 10597 18031 10655 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 10980 18068 11008 18176
rect 11146 18164 11152 18216
rect 11204 18204 11210 18216
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 11204 18176 11529 18204
rect 11204 18164 11210 18176
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 11517 18167 11575 18173
rect 12250 18164 12256 18216
rect 12308 18164 12314 18216
rect 13170 18164 13176 18216
rect 13228 18204 13234 18216
rect 13280 18204 13308 18235
rect 13538 18232 13544 18284
rect 13596 18272 13602 18284
rect 13725 18275 13783 18281
rect 13725 18272 13737 18275
rect 13596 18244 13737 18272
rect 13596 18232 13602 18244
rect 13725 18241 13737 18244
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 13998 18232 14004 18284
rect 14056 18232 14062 18284
rect 21082 18232 21088 18284
rect 21140 18232 21146 18284
rect 21266 18232 21272 18284
rect 21324 18232 21330 18284
rect 21358 18232 21364 18284
rect 21416 18232 21422 18284
rect 22066 18272 22094 18300
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 22066 18244 22201 18272
rect 22189 18241 22201 18244
rect 22235 18241 22247 18275
rect 23400 18272 23428 18303
rect 23474 18300 23480 18352
rect 23532 18340 23538 18352
rect 23532 18312 23796 18340
rect 23532 18300 23538 18312
rect 23768 18284 23796 18312
rect 24210 18300 24216 18352
rect 24268 18340 24274 18352
rect 24857 18343 24915 18349
rect 24857 18340 24869 18343
rect 24268 18312 24869 18340
rect 24268 18300 24274 18312
rect 24857 18309 24869 18312
rect 24903 18309 24915 18343
rect 24857 18303 24915 18309
rect 27062 18300 27068 18352
rect 27120 18340 27126 18352
rect 27433 18343 27491 18349
rect 27120 18312 27200 18340
rect 27120 18300 27126 18312
rect 23658 18272 23664 18284
rect 23400 18244 23664 18272
rect 22189 18235 22247 18241
rect 23658 18232 23664 18244
rect 23716 18232 23722 18284
rect 23750 18232 23756 18284
rect 23808 18272 23814 18284
rect 23845 18275 23903 18281
rect 23845 18272 23857 18275
rect 23808 18244 23857 18272
rect 23808 18232 23814 18244
rect 23845 18241 23857 18244
rect 23891 18241 23903 18275
rect 23845 18235 23903 18241
rect 23934 18232 23940 18284
rect 23992 18232 23998 18284
rect 24029 18275 24087 18281
rect 24029 18241 24041 18275
rect 24075 18272 24087 18275
rect 24118 18272 24124 18284
rect 24075 18244 24124 18272
rect 24075 18241 24087 18244
rect 24029 18235 24087 18241
rect 24118 18232 24124 18244
rect 24176 18232 24182 18284
rect 24489 18275 24547 18281
rect 24489 18241 24501 18275
rect 24535 18241 24547 18275
rect 24489 18235 24547 18241
rect 15654 18204 15660 18216
rect 13228 18176 15660 18204
rect 13228 18164 13234 18176
rect 15654 18164 15660 18176
rect 15712 18164 15718 18216
rect 21726 18164 21732 18216
rect 21784 18204 21790 18216
rect 24504 18204 24532 18235
rect 25406 18232 25412 18284
rect 25464 18232 25470 18284
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18241 25559 18275
rect 25501 18235 25559 18241
rect 21784 18176 24532 18204
rect 21784 18164 21790 18176
rect 24854 18164 24860 18216
rect 24912 18204 24918 18216
rect 25038 18204 25044 18216
rect 24912 18176 25044 18204
rect 24912 18164 24918 18176
rect 25038 18164 25044 18176
rect 25096 18204 25102 18216
rect 25516 18204 25544 18235
rect 25590 18232 25596 18284
rect 25648 18272 25654 18284
rect 25685 18275 25743 18281
rect 25685 18272 25697 18275
rect 25648 18244 25697 18272
rect 25648 18232 25654 18244
rect 25685 18241 25697 18244
rect 25731 18241 25743 18275
rect 25685 18235 25743 18241
rect 25777 18275 25835 18281
rect 25777 18241 25789 18275
rect 25823 18272 25835 18275
rect 26050 18272 26056 18284
rect 25823 18244 26056 18272
rect 25823 18241 25835 18244
rect 25777 18235 25835 18241
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 26142 18232 26148 18284
rect 26200 18232 26206 18284
rect 25096 18176 25544 18204
rect 27172 18204 27200 18312
rect 27433 18309 27445 18343
rect 27479 18340 27491 18343
rect 28166 18340 28172 18352
rect 27479 18312 28172 18340
rect 27479 18309 27491 18312
rect 27433 18303 27491 18309
rect 28166 18300 28172 18312
rect 28224 18300 28230 18352
rect 32493 18343 32551 18349
rect 32493 18340 32505 18343
rect 28276 18312 32505 18340
rect 27249 18275 27307 18281
rect 27249 18241 27261 18275
rect 27295 18272 27307 18275
rect 27338 18272 27344 18284
rect 27295 18244 27344 18272
rect 27295 18241 27307 18244
rect 27249 18235 27307 18241
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 27522 18232 27528 18284
rect 27580 18232 27586 18284
rect 27617 18275 27675 18281
rect 27617 18241 27629 18275
rect 27663 18272 27675 18275
rect 27798 18272 27804 18284
rect 27663 18244 27804 18272
rect 27663 18241 27675 18244
rect 27617 18235 27675 18241
rect 27798 18232 27804 18244
rect 27856 18232 27862 18284
rect 28166 18204 28172 18216
rect 27172 18176 28172 18204
rect 25096 18164 25102 18176
rect 28166 18164 28172 18176
rect 28224 18164 28230 18216
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 13078 18136 13084 18148
rect 12584 18108 13084 18136
rect 12584 18096 12590 18108
rect 13078 18096 13084 18108
rect 13136 18096 13142 18148
rect 14001 18139 14059 18145
rect 14001 18105 14013 18139
rect 14047 18136 14059 18139
rect 18046 18136 18052 18148
rect 14047 18108 18052 18136
rect 14047 18105 14059 18108
rect 14001 18099 14059 18105
rect 18046 18096 18052 18108
rect 18104 18096 18110 18148
rect 21085 18139 21143 18145
rect 21085 18105 21097 18139
rect 21131 18136 21143 18139
rect 21174 18136 21180 18148
rect 21131 18108 21180 18136
rect 21131 18105 21143 18108
rect 21085 18099 21143 18105
rect 21174 18096 21180 18108
rect 21232 18096 21238 18148
rect 24670 18096 24676 18148
rect 24728 18136 24734 18148
rect 24728 18108 25544 18136
rect 24728 18096 24734 18108
rect 11146 18068 11152 18080
rect 10980 18040 11152 18068
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 12805 18071 12863 18077
rect 12805 18068 12817 18071
rect 11388 18040 12817 18068
rect 11388 18028 11394 18040
rect 12805 18037 12817 18040
rect 12851 18037 12863 18071
rect 12805 18031 12863 18037
rect 20622 18028 20628 18080
rect 20680 18028 20686 18080
rect 20809 18071 20867 18077
rect 20809 18037 20821 18071
rect 20855 18068 20867 18071
rect 22002 18068 22008 18080
rect 20855 18040 22008 18068
rect 20855 18037 20867 18040
rect 20809 18031 20867 18037
rect 22002 18028 22008 18040
rect 22060 18068 22066 18080
rect 23201 18071 23259 18077
rect 23201 18068 23213 18071
rect 22060 18040 23213 18068
rect 22060 18028 22066 18040
rect 23201 18037 23213 18040
rect 23247 18068 23259 18071
rect 24394 18068 24400 18080
rect 23247 18040 24400 18068
rect 23247 18037 23259 18040
rect 23201 18031 23259 18037
rect 24394 18028 24400 18040
rect 24452 18028 24458 18080
rect 25225 18071 25283 18077
rect 25225 18037 25237 18071
rect 25271 18068 25283 18071
rect 25406 18068 25412 18080
rect 25271 18040 25412 18068
rect 25271 18037 25283 18040
rect 25225 18031 25283 18037
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 25516 18068 25544 18108
rect 25682 18096 25688 18148
rect 25740 18136 25746 18148
rect 28276 18136 28304 18312
rect 32493 18309 32505 18312
rect 32539 18309 32551 18343
rect 33594 18340 33600 18352
rect 32493 18303 32551 18309
rect 32692 18312 33600 18340
rect 28994 18232 29000 18284
rect 29052 18272 29058 18284
rect 29638 18272 29644 18284
rect 29052 18244 29644 18272
rect 29052 18232 29058 18244
rect 29638 18232 29644 18244
rect 29696 18272 29702 18284
rect 32692 18281 32720 18312
rect 33594 18300 33600 18312
rect 33652 18300 33658 18352
rect 33686 18300 33692 18352
rect 33744 18300 33750 18352
rect 32263 18275 32321 18281
rect 32263 18272 32275 18275
rect 29696 18244 32275 18272
rect 29696 18232 29702 18244
rect 32263 18241 32275 18244
rect 32309 18241 32321 18275
rect 32263 18235 32321 18241
rect 32401 18275 32459 18281
rect 32401 18241 32413 18275
rect 32447 18241 32459 18275
rect 32401 18235 32459 18241
rect 32676 18275 32734 18281
rect 32676 18241 32688 18275
rect 32722 18241 32734 18275
rect 32676 18235 32734 18241
rect 32416 18204 32444 18235
rect 32766 18232 32772 18284
rect 32824 18232 32830 18284
rect 32950 18232 32956 18284
rect 33008 18232 33014 18284
rect 33318 18232 33324 18284
rect 33376 18272 33382 18284
rect 33505 18275 33563 18281
rect 33505 18272 33517 18275
rect 33376 18244 33517 18272
rect 33376 18232 33382 18244
rect 33505 18241 33517 18244
rect 33551 18241 33563 18275
rect 33505 18235 33563 18241
rect 33778 18232 33784 18284
rect 33836 18232 33842 18284
rect 33888 18281 33916 18380
rect 34057 18377 34069 18411
rect 34103 18377 34115 18411
rect 34057 18371 34115 18377
rect 34072 18340 34100 18371
rect 35250 18368 35256 18420
rect 35308 18368 35314 18420
rect 34330 18340 34336 18352
rect 34072 18312 34336 18340
rect 34330 18300 34336 18312
rect 34388 18340 34394 18352
rect 35069 18343 35127 18349
rect 35069 18340 35081 18343
rect 34388 18312 35081 18340
rect 34388 18300 34394 18312
rect 35069 18309 35081 18312
rect 35115 18309 35127 18343
rect 35069 18303 35127 18309
rect 35342 18300 35348 18352
rect 35400 18300 35406 18352
rect 33873 18275 33931 18281
rect 33873 18241 33885 18275
rect 33919 18241 33931 18275
rect 33873 18235 33931 18241
rect 34885 18275 34943 18281
rect 34885 18241 34897 18275
rect 34931 18241 34943 18275
rect 34885 18235 34943 18241
rect 33229 18207 33287 18213
rect 33229 18204 33241 18207
rect 31726 18176 33241 18204
rect 31726 18136 31754 18176
rect 33229 18173 33241 18176
rect 33275 18173 33287 18207
rect 33229 18167 33287 18173
rect 25740 18108 28304 18136
rect 28368 18108 31754 18136
rect 25740 18096 25746 18108
rect 28368 18068 28396 18108
rect 31938 18096 31944 18148
rect 31996 18136 32002 18148
rect 32125 18139 32183 18145
rect 32125 18136 32137 18139
rect 31996 18108 32137 18136
rect 31996 18096 32002 18108
rect 32125 18105 32137 18108
rect 32171 18136 32183 18139
rect 34900 18136 34928 18235
rect 35434 18232 35440 18284
rect 35492 18272 35498 18284
rect 35529 18275 35587 18281
rect 35529 18272 35541 18275
rect 35492 18244 35541 18272
rect 35492 18232 35498 18244
rect 35529 18241 35541 18244
rect 35575 18241 35587 18275
rect 35529 18235 35587 18241
rect 32171 18108 34928 18136
rect 32171 18105 32183 18108
rect 32125 18099 32183 18105
rect 25516 18040 28396 18068
rect 29822 18028 29828 18080
rect 29880 18068 29886 18080
rect 31202 18068 31208 18080
rect 29880 18040 31208 18068
rect 29880 18028 29886 18040
rect 31202 18028 31208 18040
rect 31260 18028 31266 18080
rect 34606 18028 34612 18080
rect 34664 18068 34670 18080
rect 35713 18071 35771 18077
rect 35713 18068 35725 18071
rect 34664 18040 35725 18068
rect 34664 18028 34670 18040
rect 35713 18037 35725 18040
rect 35759 18037 35771 18071
rect 35713 18031 35771 18037
rect 1104 17978 36432 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 36432 17978
rect 1104 17904 36432 17926
rect 3326 17864 3332 17876
rect 2884 17836 3332 17864
rect 2314 17620 2320 17672
rect 2372 17660 2378 17672
rect 2593 17663 2651 17669
rect 2593 17660 2605 17663
rect 2372 17632 2605 17660
rect 2372 17620 2378 17632
rect 2593 17629 2605 17632
rect 2639 17629 2651 17663
rect 2593 17623 2651 17629
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17660 2835 17663
rect 2884 17660 2912 17836
rect 3326 17824 3332 17836
rect 3384 17824 3390 17876
rect 4433 17867 4491 17873
rect 4433 17833 4445 17867
rect 4479 17864 4491 17867
rect 4614 17864 4620 17876
rect 4479 17836 4620 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5810 17864 5816 17876
rect 4724 17836 5816 17864
rect 4338 17728 4344 17740
rect 2976 17700 4344 17728
rect 2976 17669 3004 17700
rect 4338 17688 4344 17700
rect 4396 17688 4402 17740
rect 4724 17728 4752 17836
rect 5810 17824 5816 17836
rect 5868 17824 5874 17876
rect 7098 17824 7104 17876
rect 7156 17824 7162 17876
rect 10137 17867 10195 17873
rect 10137 17833 10149 17867
rect 10183 17864 10195 17867
rect 11238 17864 11244 17876
rect 10183 17836 11244 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 11238 17824 11244 17836
rect 11296 17864 11302 17876
rect 11333 17867 11391 17873
rect 11333 17864 11345 17867
rect 11296 17836 11345 17864
rect 11296 17824 11302 17836
rect 11333 17833 11345 17836
rect 11379 17833 11391 17867
rect 11333 17827 11391 17833
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 11701 17867 11759 17873
rect 11701 17864 11713 17867
rect 11480 17836 11713 17864
rect 11480 17824 11486 17836
rect 11701 17833 11713 17836
rect 11747 17864 11759 17867
rect 12158 17864 12164 17876
rect 11747 17836 12164 17864
rect 11747 17833 11759 17836
rect 11701 17827 11759 17833
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 12434 17824 12440 17876
rect 12492 17824 12498 17876
rect 13998 17824 14004 17876
rect 14056 17864 14062 17876
rect 14093 17867 14151 17873
rect 14093 17864 14105 17867
rect 14056 17836 14105 17864
rect 14056 17824 14062 17836
rect 14093 17833 14105 17836
rect 14139 17833 14151 17867
rect 14093 17827 14151 17833
rect 14369 17867 14427 17873
rect 14369 17833 14381 17867
rect 14415 17864 14427 17867
rect 14642 17864 14648 17876
rect 14415 17836 14648 17864
rect 14415 17833 14427 17836
rect 14369 17827 14427 17833
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 15102 17824 15108 17876
rect 15160 17864 15166 17876
rect 18598 17864 18604 17876
rect 15160 17836 18604 17864
rect 15160 17824 15166 17836
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 18693 17867 18751 17873
rect 18693 17833 18705 17867
rect 18739 17864 18751 17867
rect 18874 17864 18880 17876
rect 18739 17836 18880 17864
rect 18739 17833 18751 17836
rect 18693 17827 18751 17833
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 21634 17864 21640 17876
rect 20772 17836 21640 17864
rect 20772 17824 20778 17836
rect 21634 17824 21640 17836
rect 21692 17864 21698 17876
rect 22005 17867 22063 17873
rect 22005 17864 22017 17867
rect 21692 17836 22017 17864
rect 21692 17824 21698 17836
rect 22005 17833 22017 17836
rect 22051 17833 22063 17867
rect 22005 17827 22063 17833
rect 22370 17824 22376 17876
rect 22428 17824 22434 17876
rect 23658 17824 23664 17876
rect 23716 17864 23722 17876
rect 24670 17864 24676 17876
rect 23716 17836 24676 17864
rect 23716 17824 23722 17836
rect 24670 17824 24676 17836
rect 24728 17824 24734 17876
rect 24946 17824 24952 17876
rect 25004 17864 25010 17876
rect 25774 17864 25780 17876
rect 25004 17836 25780 17864
rect 25004 17824 25010 17836
rect 25774 17824 25780 17836
rect 25832 17824 25838 17876
rect 28902 17824 28908 17876
rect 28960 17864 28966 17876
rect 30377 17867 30435 17873
rect 30377 17864 30389 17867
rect 28960 17836 30389 17864
rect 28960 17824 28966 17836
rect 30377 17833 30389 17836
rect 30423 17833 30435 17867
rect 30377 17827 30435 17833
rect 31478 17824 31484 17876
rect 31536 17864 31542 17876
rect 31662 17864 31668 17876
rect 31536 17836 31668 17864
rect 31536 17824 31542 17836
rect 31662 17824 31668 17836
rect 31720 17824 31726 17876
rect 34330 17824 34336 17876
rect 34388 17824 34394 17876
rect 34514 17824 34520 17876
rect 34572 17824 34578 17876
rect 4632 17700 4752 17728
rect 7116 17728 7144 17824
rect 9030 17756 9036 17808
rect 9088 17796 9094 17808
rect 9217 17799 9275 17805
rect 9217 17796 9229 17799
rect 9088 17768 9229 17796
rect 9088 17756 9094 17768
rect 9217 17765 9229 17768
rect 9263 17765 9275 17799
rect 9217 17759 9275 17765
rect 10226 17756 10232 17808
rect 10284 17756 10290 17808
rect 10686 17756 10692 17808
rect 10744 17796 10750 17808
rect 14734 17796 14740 17808
rect 10744 17768 12204 17796
rect 10744 17756 10750 17768
rect 7745 17731 7803 17737
rect 7745 17728 7757 17731
rect 7116 17700 7757 17728
rect 2823 17632 2912 17660
rect 2961 17663 3019 17669
rect 2823 17629 2835 17632
rect 2777 17623 2835 17629
rect 2961 17629 2973 17663
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 3418 17620 3424 17672
rect 3476 17660 3482 17672
rect 3786 17660 3792 17672
rect 3476 17632 3792 17660
rect 3476 17620 3482 17632
rect 3786 17620 3792 17632
rect 3844 17660 3850 17672
rect 3881 17663 3939 17669
rect 3881 17660 3893 17663
rect 3844 17632 3893 17660
rect 3844 17620 3850 17632
rect 3881 17629 3893 17632
rect 3927 17629 3939 17663
rect 3881 17623 3939 17629
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4295 17629 4318 17660
rect 4249 17623 4318 17629
rect 2869 17595 2927 17601
rect 2869 17561 2881 17595
rect 2915 17592 2927 17595
rect 3050 17592 3056 17604
rect 2915 17564 3056 17592
rect 2915 17561 2927 17564
rect 2869 17555 2927 17561
rect 3050 17552 3056 17564
rect 3108 17552 3114 17604
rect 3234 17552 3240 17604
rect 3292 17592 3298 17604
rect 3602 17592 3608 17604
rect 3292 17564 3608 17592
rect 3292 17552 3298 17564
rect 3602 17552 3608 17564
rect 3660 17592 3666 17604
rect 4065 17595 4123 17601
rect 4065 17592 4077 17595
rect 3660 17564 4077 17592
rect 3660 17552 3666 17564
rect 4065 17561 4077 17564
rect 4111 17561 4123 17595
rect 4065 17555 4123 17561
rect 4154 17552 4160 17604
rect 4212 17552 4218 17604
rect 4290 17592 4318 17623
rect 4522 17620 4528 17672
rect 4580 17660 4586 17672
rect 4632 17669 4660 17700
rect 7745 17697 7757 17700
rect 7791 17697 7803 17731
rect 7745 17691 7803 17697
rect 8478 17688 8484 17740
rect 8536 17688 8542 17740
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 9309 17731 9367 17737
rect 9309 17728 9321 17731
rect 8628 17700 9321 17728
rect 8628 17688 8634 17700
rect 9309 17697 9321 17700
rect 9355 17697 9367 17731
rect 9309 17691 9367 17697
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10235 17728 10263 17756
rect 9732 17700 10088 17728
rect 10235 17700 10364 17728
rect 9732 17688 9738 17700
rect 4617 17663 4675 17669
rect 4617 17660 4629 17663
rect 4580 17632 4629 17660
rect 4580 17620 4586 17632
rect 4617 17629 4629 17632
rect 4663 17629 4675 17663
rect 4617 17623 4675 17629
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 4798 17620 4804 17672
rect 4856 17620 4862 17672
rect 4890 17620 4896 17672
rect 4948 17620 4954 17672
rect 5350 17620 5356 17672
rect 5408 17620 5414 17672
rect 6638 17620 6644 17672
rect 6696 17660 6702 17672
rect 7926 17660 7932 17672
rect 6696 17632 7932 17660
rect 6696 17620 6702 17632
rect 7926 17620 7932 17632
rect 7984 17620 7990 17672
rect 8941 17663 8999 17669
rect 8941 17660 8953 17663
rect 8128 17632 8953 17660
rect 5077 17595 5135 17601
rect 4290 17564 4936 17592
rect 3145 17527 3203 17533
rect 3145 17493 3157 17527
rect 3191 17524 3203 17527
rect 4798 17524 4804 17536
rect 3191 17496 4804 17524
rect 3191 17493 3203 17496
rect 3145 17487 3203 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 4908 17524 4936 17564
rect 5077 17561 5089 17595
rect 5123 17592 5135 17595
rect 5534 17592 5540 17604
rect 5123 17564 5540 17592
rect 5123 17561 5135 17564
rect 5077 17555 5135 17561
rect 5534 17552 5540 17564
rect 5592 17552 5598 17604
rect 5626 17552 5632 17604
rect 5684 17552 5690 17604
rect 7742 17552 7748 17604
rect 7800 17592 7806 17604
rect 8128 17592 8156 17632
rect 8941 17629 8953 17632
rect 8987 17629 8999 17663
rect 8941 17623 8999 17629
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17660 9459 17663
rect 9447 17632 9812 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 7800 17564 8156 17592
rect 8297 17595 8355 17601
rect 7800 17552 7806 17564
rect 8297 17561 8309 17595
rect 8343 17592 8355 17595
rect 9030 17592 9036 17604
rect 8343 17564 9036 17592
rect 8343 17561 8355 17564
rect 8297 17555 8355 17561
rect 9030 17552 9036 17564
rect 9088 17592 9094 17604
rect 9490 17592 9496 17604
rect 9088 17564 9496 17592
rect 9088 17552 9094 17564
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 5902 17524 5908 17536
rect 4908 17496 5908 17524
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 7190 17484 7196 17536
rect 7248 17484 7254 17536
rect 7558 17484 7564 17536
rect 7616 17524 7622 17536
rect 7929 17527 7987 17533
rect 7929 17524 7941 17527
rect 7616 17496 7941 17524
rect 7616 17484 7622 17496
rect 7929 17493 7941 17496
rect 7975 17493 7987 17527
rect 7929 17487 7987 17493
rect 8389 17527 8447 17533
rect 8389 17493 8401 17527
rect 8435 17524 8447 17527
rect 9306 17524 9312 17536
rect 8435 17496 9312 17524
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 9674 17484 9680 17536
rect 9732 17484 9738 17536
rect 9784 17524 9812 17632
rect 9858 17620 9864 17672
rect 9916 17620 9922 17672
rect 10060 17669 10088 17700
rect 10336 17669 10364 17700
rect 10410 17688 10416 17740
rect 10468 17728 10474 17740
rect 10468 17700 12112 17728
rect 10468 17688 10474 17700
rect 10045 17663 10103 17669
rect 10321 17663 10379 17669
rect 10045 17629 10057 17663
rect 10091 17629 10103 17663
rect 10220 17657 10278 17663
rect 10220 17654 10232 17657
rect 10045 17623 10103 17629
rect 10152 17626 10232 17654
rect 10152 17536 10180 17626
rect 10220 17623 10232 17626
rect 10266 17623 10278 17657
rect 10321 17629 10333 17663
rect 10367 17629 10379 17663
rect 10321 17623 10379 17629
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17660 10563 17663
rect 10686 17660 10692 17672
rect 10551 17632 10692 17660
rect 10551 17629 10563 17632
rect 10505 17623 10563 17629
rect 10220 17617 10278 17623
rect 10686 17620 10692 17632
rect 10744 17620 10750 17672
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17629 10931 17663
rect 10873 17623 10931 17629
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17662 11115 17663
rect 11103 17660 11284 17662
rect 11422 17660 11428 17672
rect 11103 17634 11428 17660
rect 11103 17629 11115 17634
rect 11256 17632 11428 17634
rect 11057 17623 11115 17629
rect 10042 17524 10048 17536
rect 9784 17496 10048 17524
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 10134 17484 10140 17536
rect 10192 17484 10198 17536
rect 10502 17484 10508 17536
rect 10560 17484 10566 17536
rect 10686 17484 10692 17536
rect 10744 17524 10750 17536
rect 10781 17527 10839 17533
rect 10781 17524 10793 17527
rect 10744 17496 10793 17524
rect 10744 17484 10750 17496
rect 10781 17493 10793 17496
rect 10827 17493 10839 17527
rect 10888 17524 10916 17623
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 11514 17620 11520 17672
rect 11572 17620 11578 17672
rect 11882 17669 11888 17672
rect 11880 17660 11888 17669
rect 11843 17632 11888 17660
rect 11880 17623 11888 17632
rect 11882 17620 11888 17623
rect 11940 17620 11946 17672
rect 11146 17552 11152 17604
rect 11204 17552 11210 17604
rect 11333 17595 11391 17601
rect 11333 17561 11345 17595
rect 11379 17592 11391 17595
rect 11532 17592 11560 17620
rect 11379 17564 11560 17592
rect 11379 17561 11391 17564
rect 11333 17555 11391 17561
rect 11348 17524 11376 17555
rect 11790 17552 11796 17604
rect 11848 17592 11854 17604
rect 12084 17601 12112 17700
rect 12176 17672 12204 17768
rect 13004 17768 14740 17796
rect 13004 17672 13032 17768
rect 14734 17756 14740 17768
rect 14792 17756 14798 17808
rect 14918 17756 14924 17808
rect 14976 17796 14982 17808
rect 20257 17799 20315 17805
rect 20257 17796 20269 17799
rect 14976 17768 20269 17796
rect 14976 17756 14982 17768
rect 20257 17765 20269 17768
rect 20303 17765 20315 17799
rect 20257 17759 20315 17765
rect 21818 17756 21824 17808
rect 21876 17796 21882 17808
rect 22388 17796 22416 17824
rect 21876 17768 22416 17796
rect 22741 17799 22799 17805
rect 21876 17756 21882 17768
rect 22741 17765 22753 17799
rect 22787 17796 22799 17799
rect 23014 17796 23020 17808
rect 22787 17768 23020 17796
rect 22787 17765 22799 17768
rect 22741 17759 22799 17765
rect 23014 17756 23020 17768
rect 23072 17756 23078 17808
rect 23477 17799 23535 17805
rect 23477 17765 23489 17799
rect 23523 17796 23535 17799
rect 24486 17796 24492 17808
rect 23523 17768 24492 17796
rect 23523 17765 23535 17768
rect 23477 17759 23535 17765
rect 24486 17756 24492 17768
rect 24544 17756 24550 17808
rect 25130 17756 25136 17808
rect 25188 17796 25194 17808
rect 25188 17768 31708 17796
rect 25188 17756 25194 17768
rect 31680 17740 31708 17768
rect 14553 17731 14611 17737
rect 14553 17697 14565 17731
rect 14599 17697 14611 17731
rect 17221 17731 17279 17737
rect 17221 17728 17233 17731
rect 14553 17691 14611 17697
rect 14752 17700 17233 17728
rect 12158 17620 12164 17672
rect 12216 17669 12222 17672
rect 12216 17663 12255 17669
rect 12243 17629 12255 17663
rect 12216 17623 12255 17629
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 12434 17660 12440 17672
rect 12391 17632 12440 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 12216 17620 12222 17623
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 12618 17620 12624 17672
rect 12676 17620 12682 17672
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17660 12863 17663
rect 12986 17660 12992 17672
rect 12851 17632 12992 17660
rect 12851 17629 12863 17632
rect 12805 17623 12863 17629
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 14458 17620 14464 17672
rect 14516 17620 14522 17672
rect 14568 17660 14596 17691
rect 14752 17660 14780 17700
rect 14568 17632 14780 17660
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17660 14887 17663
rect 15010 17660 15016 17672
rect 14875 17632 15016 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15378 17620 15384 17672
rect 15436 17660 15442 17672
rect 15657 17663 15715 17669
rect 15657 17660 15669 17663
rect 15436 17632 15669 17660
rect 15436 17620 15442 17632
rect 15657 17629 15669 17632
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 15746 17620 15752 17672
rect 15804 17620 15810 17672
rect 15948 17669 15976 17700
rect 17221 17697 17233 17700
rect 17267 17697 17279 17731
rect 17221 17691 17279 17697
rect 17586 17688 17592 17740
rect 17644 17728 17650 17740
rect 17644 17700 18552 17728
rect 17644 17688 17650 17700
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 16022 17620 16028 17672
rect 16080 17620 16086 17672
rect 17402 17620 17408 17672
rect 17460 17620 17466 17672
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17629 17555 17663
rect 17497 17623 17555 17629
rect 11977 17595 12035 17601
rect 11977 17592 11989 17595
rect 11848 17564 11989 17592
rect 11848 17552 11854 17564
rect 11977 17561 11989 17564
rect 12023 17561 12035 17595
rect 11977 17555 12035 17561
rect 12069 17595 12127 17601
rect 12069 17561 12081 17595
rect 12115 17592 12127 17595
rect 13170 17592 13176 17604
rect 12115 17564 13176 17592
rect 12115 17561 12127 17564
rect 12069 17555 12127 17561
rect 13170 17552 13176 17564
rect 13228 17552 13234 17604
rect 15028 17592 15056 17620
rect 16942 17592 16948 17604
rect 15028 17564 16948 17592
rect 16942 17552 16948 17564
rect 17000 17552 17006 17604
rect 17512 17592 17540 17623
rect 17678 17620 17684 17672
rect 17736 17620 17742 17672
rect 18524 17669 18552 17700
rect 20530 17688 20536 17740
rect 20588 17688 20594 17740
rect 22002 17688 22008 17740
rect 22060 17688 22066 17740
rect 26970 17728 26976 17740
rect 23492 17700 26976 17728
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17660 17831 17663
rect 18509 17663 18567 17669
rect 17819 17632 18276 17660
rect 17819 17629 17831 17632
rect 17773 17623 17831 17629
rect 17954 17592 17960 17604
rect 17512 17564 17960 17592
rect 17954 17552 17960 17564
rect 18012 17552 18018 17604
rect 18248 17601 18276 17632
rect 18509 17629 18521 17663
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17660 18843 17663
rect 18966 17660 18972 17672
rect 18831 17632 18972 17660
rect 18831 17629 18843 17632
rect 18785 17623 18843 17629
rect 18049 17595 18107 17601
rect 18049 17561 18061 17595
rect 18095 17561 18107 17595
rect 18049 17555 18107 17561
rect 18233 17595 18291 17601
rect 18233 17561 18245 17595
rect 18279 17592 18291 17595
rect 18325 17595 18383 17601
rect 18325 17592 18337 17595
rect 18279 17564 18337 17592
rect 18279 17561 18291 17564
rect 18233 17555 18291 17561
rect 18325 17561 18337 17564
rect 18371 17561 18383 17595
rect 18524 17592 18552 17623
rect 18966 17620 18972 17632
rect 19024 17620 19030 17672
rect 20254 17620 20260 17672
rect 20312 17660 20318 17672
rect 20548 17660 20576 17688
rect 20312 17632 20576 17660
rect 20993 17663 21051 17669
rect 20312 17620 20318 17632
rect 20993 17629 21005 17663
rect 21039 17660 21051 17663
rect 21174 17660 21180 17672
rect 21039 17632 21180 17660
rect 21039 17629 21051 17632
rect 20993 17623 21051 17629
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 21358 17620 21364 17672
rect 21416 17620 21422 17672
rect 21450 17620 21456 17672
rect 21508 17620 21514 17672
rect 22020 17660 22048 17688
rect 21988 17635 22048 17660
rect 21959 17632 22048 17635
rect 21959 17629 22017 17632
rect 19886 17592 19892 17604
rect 18524 17564 19892 17592
rect 18325 17555 18383 17561
rect 10888 17496 11376 17524
rect 10781 17487 10839 17493
rect 11422 17484 11428 17536
rect 11480 17524 11486 17536
rect 11517 17527 11575 17533
rect 11517 17524 11529 17527
rect 11480 17496 11529 17524
rect 11480 17484 11486 17496
rect 11517 17493 11529 17496
rect 11563 17493 11575 17527
rect 11517 17487 11575 17493
rect 14737 17527 14795 17533
rect 14737 17493 14749 17527
rect 14783 17524 14795 17527
rect 15102 17524 15108 17536
rect 14783 17496 15108 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 15378 17484 15384 17536
rect 15436 17524 15442 17536
rect 15473 17527 15531 17533
rect 15473 17524 15485 17527
rect 15436 17496 15485 17524
rect 15436 17484 15442 17496
rect 15473 17493 15485 17496
rect 15519 17493 15531 17527
rect 15473 17487 15531 17493
rect 17034 17484 17040 17536
rect 17092 17524 17098 17536
rect 17865 17527 17923 17533
rect 17865 17524 17877 17527
rect 17092 17496 17877 17524
rect 17092 17484 17098 17496
rect 17865 17493 17877 17496
rect 17911 17493 17923 17527
rect 18064 17524 18092 17555
rect 19886 17552 19892 17564
rect 19944 17552 19950 17604
rect 21959 17595 21971 17629
rect 22005 17595 22017 17629
rect 22554 17620 22560 17672
rect 22612 17660 22618 17672
rect 22649 17663 22707 17669
rect 22649 17660 22661 17663
rect 22612 17632 22661 17660
rect 22612 17620 22618 17632
rect 22649 17629 22661 17632
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 22830 17620 22836 17672
rect 22888 17620 22894 17672
rect 22925 17663 22983 17669
rect 22925 17629 22937 17663
rect 22971 17660 22983 17663
rect 23014 17660 23020 17672
rect 22971 17632 23020 17660
rect 22971 17629 22983 17632
rect 22925 17623 22983 17629
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 23106 17620 23112 17672
rect 23164 17660 23170 17672
rect 23492 17660 23520 17700
rect 26970 17688 26976 17700
rect 27028 17688 27034 17740
rect 29546 17688 29552 17740
rect 29604 17728 29610 17740
rect 30469 17731 30527 17737
rect 30469 17728 30481 17731
rect 29604 17700 30481 17728
rect 29604 17688 29610 17700
rect 30469 17697 30481 17700
rect 30515 17697 30527 17731
rect 30469 17691 30527 17697
rect 31662 17688 31668 17740
rect 31720 17688 31726 17740
rect 23164 17632 23520 17660
rect 23164 17620 23170 17632
rect 23750 17620 23756 17672
rect 23808 17660 23814 17672
rect 27430 17660 27436 17672
rect 23808 17632 27436 17660
rect 23808 17620 23814 17632
rect 21959 17589 22017 17595
rect 22094 17552 22100 17604
rect 22152 17592 22158 17604
rect 23860 17601 23888 17632
rect 27430 17620 27436 17632
rect 27488 17620 27494 17672
rect 28810 17620 28816 17672
rect 28868 17620 28874 17672
rect 22189 17595 22247 17601
rect 22189 17592 22201 17595
rect 22152 17564 22201 17592
rect 22152 17552 22158 17564
rect 22189 17561 22201 17564
rect 22235 17561 22247 17595
rect 23845 17595 23903 17601
rect 22189 17555 22247 17561
rect 22296 17564 23688 17592
rect 21082 17524 21088 17536
rect 18064 17496 21088 17524
rect 17865 17487 17923 17493
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 21818 17484 21824 17536
rect 21876 17484 21882 17536
rect 22002 17484 22008 17536
rect 22060 17524 22066 17536
rect 22296 17524 22324 17564
rect 22060 17496 22324 17524
rect 22060 17484 22066 17496
rect 22830 17484 22836 17536
rect 22888 17524 22894 17536
rect 23660 17533 23688 17564
rect 23845 17561 23857 17595
rect 23891 17561 23903 17595
rect 29270 17592 29276 17604
rect 23845 17555 23903 17561
rect 28966 17564 29276 17592
rect 23109 17527 23167 17533
rect 23109 17524 23121 17527
rect 22888 17496 23121 17524
rect 22888 17484 22894 17496
rect 23109 17493 23121 17496
rect 23155 17493 23167 17527
rect 23109 17487 23167 17493
rect 23645 17527 23703 17533
rect 23645 17493 23657 17527
rect 23691 17524 23703 17527
rect 28966 17524 28994 17564
rect 29270 17552 29276 17564
rect 29328 17552 29334 17604
rect 29564 17533 29592 17688
rect 29638 17620 29644 17672
rect 29696 17660 29702 17672
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 29696 17632 29745 17660
rect 29696 17620 29702 17632
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 30098 17620 30104 17672
rect 30156 17620 30162 17672
rect 30377 17663 30435 17669
rect 30377 17629 30389 17663
rect 30423 17629 30435 17663
rect 30377 17623 30435 17629
rect 29822 17552 29828 17604
rect 29880 17552 29886 17604
rect 29917 17595 29975 17601
rect 29917 17561 29929 17595
rect 29963 17592 29975 17595
rect 30006 17592 30012 17604
rect 29963 17564 30012 17592
rect 29963 17561 29975 17564
rect 29917 17555 29975 17561
rect 30006 17552 30012 17564
rect 30064 17552 30070 17604
rect 30392 17592 30420 17623
rect 30558 17620 30564 17672
rect 30616 17660 30622 17672
rect 30653 17663 30711 17669
rect 30653 17660 30665 17663
rect 30616 17632 30665 17660
rect 30616 17620 30622 17632
rect 30653 17629 30665 17632
rect 30699 17629 30711 17663
rect 30653 17623 30711 17629
rect 32766 17620 32772 17672
rect 32824 17660 32830 17672
rect 34149 17663 34207 17669
rect 34149 17660 34161 17663
rect 32824 17632 34161 17660
rect 32824 17620 32830 17632
rect 34149 17629 34161 17632
rect 34195 17629 34207 17663
rect 34149 17623 34207 17629
rect 34241 17663 34299 17669
rect 34241 17629 34253 17663
rect 34287 17629 34299 17663
rect 34241 17623 34299 17629
rect 30116 17564 30420 17592
rect 23691 17496 28994 17524
rect 29549 17527 29607 17533
rect 23691 17493 23703 17496
rect 23645 17487 23703 17493
rect 29549 17493 29561 17527
rect 29595 17493 29607 17527
rect 29549 17487 29607 17493
rect 29638 17484 29644 17536
rect 29696 17524 29702 17536
rect 30116 17524 30144 17564
rect 30466 17552 30472 17604
rect 30524 17592 30530 17604
rect 34256 17592 34284 17623
rect 30524 17564 34284 17592
rect 30524 17552 30530 17564
rect 29696 17496 30144 17524
rect 30193 17527 30251 17533
rect 29696 17484 29702 17496
rect 30193 17493 30205 17527
rect 30239 17524 30251 17527
rect 30282 17524 30288 17536
rect 30239 17496 30288 17524
rect 30239 17493 30251 17496
rect 30193 17487 30251 17493
rect 30282 17484 30288 17496
rect 30340 17484 30346 17536
rect 1104 17434 36432 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 36432 17434
rect 1104 17360 36432 17382
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3145 17323 3203 17329
rect 3145 17320 3157 17323
rect 3108 17292 3157 17320
rect 3108 17280 3114 17292
rect 3145 17289 3157 17292
rect 3191 17289 3203 17323
rect 3145 17283 3203 17289
rect 2774 17144 2780 17196
rect 2832 17144 2838 17196
rect 3160 17184 3188 17283
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4525 17323 4583 17329
rect 4525 17320 4537 17323
rect 4304 17292 4537 17320
rect 4304 17280 4310 17292
rect 4525 17289 4537 17292
rect 4571 17289 4583 17323
rect 5534 17320 5540 17332
rect 4525 17283 4583 17289
rect 4632 17292 5540 17320
rect 3602 17212 3608 17264
rect 3660 17252 3666 17264
rect 4157 17255 4215 17261
rect 4157 17252 4169 17255
rect 3660 17224 4169 17252
rect 3660 17212 3666 17224
rect 4157 17221 4169 17224
rect 4203 17252 4215 17255
rect 4632 17252 4660 17292
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 5626 17280 5632 17332
rect 5684 17320 5690 17332
rect 6365 17323 6423 17329
rect 6365 17320 6377 17323
rect 5684 17292 6377 17320
rect 5684 17280 5690 17292
rect 6365 17289 6377 17292
rect 6411 17289 6423 17323
rect 6365 17283 6423 17289
rect 6733 17323 6791 17329
rect 6733 17289 6745 17323
rect 6779 17320 6791 17323
rect 7190 17320 7196 17332
rect 6779 17292 7196 17320
rect 6779 17289 6791 17292
rect 6733 17283 6791 17289
rect 7190 17280 7196 17292
rect 7248 17280 7254 17332
rect 7926 17280 7932 17332
rect 7984 17320 7990 17332
rect 9033 17323 9091 17329
rect 7984 17292 8892 17320
rect 7984 17280 7990 17292
rect 4203 17224 4660 17252
rect 4203 17221 4215 17224
rect 4157 17215 4215 17221
rect 4798 17212 4804 17264
rect 4856 17252 4862 17264
rect 4856 17224 5028 17252
rect 4856 17212 4862 17224
rect 3789 17187 3847 17193
rect 3789 17184 3801 17187
rect 3160 17156 3801 17184
rect 3789 17153 3801 17156
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 3970 17144 3976 17196
rect 4028 17144 4034 17196
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17153 4307 17187
rect 4249 17147 4307 17153
rect 1394 17076 1400 17128
rect 1452 17076 1458 17128
rect 1670 17076 1676 17128
rect 1728 17076 1734 17128
rect 4264 17116 4292 17147
rect 4338 17144 4344 17196
rect 4396 17144 4402 17196
rect 4522 17144 4528 17196
rect 4580 17184 4586 17196
rect 5000 17193 5028 17224
rect 5350 17212 5356 17264
rect 5408 17252 5414 17264
rect 6914 17252 6920 17264
rect 5408 17224 6920 17252
rect 5408 17212 5414 17224
rect 6914 17212 6920 17224
rect 6972 17252 6978 17264
rect 6972 17224 7328 17252
rect 6972 17212 6978 17224
rect 4893 17187 4951 17193
rect 4893 17184 4905 17187
rect 4580 17156 4905 17184
rect 4580 17144 4586 17156
rect 4893 17153 4905 17156
rect 4939 17153 4951 17187
rect 4893 17147 4951 17153
rect 4985 17187 5043 17193
rect 4985 17153 4997 17187
rect 5031 17153 5043 17187
rect 4985 17147 5043 17153
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17184 5227 17187
rect 5445 17187 5503 17193
rect 5445 17184 5457 17187
rect 5215 17156 5457 17184
rect 5215 17153 5227 17156
rect 5169 17147 5227 17153
rect 5445 17153 5457 17156
rect 5491 17153 5503 17187
rect 5445 17147 5503 17153
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 5718 17184 5724 17196
rect 5675 17156 5724 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 5810 17144 5816 17196
rect 5868 17144 5874 17196
rect 5902 17144 5908 17196
rect 5960 17144 5966 17196
rect 7300 17193 7328 17224
rect 7558 17212 7564 17264
rect 7616 17212 7622 17264
rect 8864 17252 8892 17292
rect 9033 17289 9045 17323
rect 9079 17320 9091 17323
rect 9306 17320 9312 17332
rect 9079 17292 9312 17320
rect 9079 17289 9091 17292
rect 9033 17283 9091 17289
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 9766 17320 9772 17332
rect 9416 17292 9772 17320
rect 9416 17252 9444 17292
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 9950 17280 9956 17332
rect 10008 17280 10014 17332
rect 10042 17280 10048 17332
rect 10100 17320 10106 17332
rect 10594 17320 10600 17332
rect 10100 17292 10600 17320
rect 10100 17280 10106 17292
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11388 17292 11621 17320
rect 11388 17280 11394 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 11698 17280 11704 17332
rect 11756 17320 11762 17332
rect 11977 17323 12035 17329
rect 11977 17320 11989 17323
rect 11756 17292 11989 17320
rect 11756 17280 11762 17292
rect 11977 17289 11989 17292
rect 12023 17289 12035 17323
rect 11977 17283 12035 17289
rect 12158 17280 12164 17332
rect 12216 17280 12222 17332
rect 12618 17280 12624 17332
rect 12676 17280 12682 17332
rect 15286 17280 15292 17332
rect 15344 17280 15350 17332
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 24949 17323 25007 17329
rect 24949 17320 24961 17323
rect 21416 17292 24961 17320
rect 21416 17280 21422 17292
rect 24949 17289 24961 17292
rect 24995 17289 25007 17323
rect 24949 17283 25007 17289
rect 27893 17323 27951 17329
rect 27893 17289 27905 17323
rect 27939 17320 27951 17323
rect 30650 17320 30656 17332
rect 27939 17292 30656 17320
rect 27939 17289 27951 17292
rect 27893 17283 27951 17289
rect 30650 17280 30656 17292
rect 30708 17280 30714 17332
rect 30745 17323 30803 17329
rect 30745 17289 30757 17323
rect 30791 17320 30803 17323
rect 31941 17323 31999 17329
rect 30791 17292 31754 17320
rect 30791 17289 30803 17292
rect 30745 17283 30803 17289
rect 8786 17224 9444 17252
rect 9493 17255 9551 17261
rect 9493 17221 9505 17255
rect 9539 17252 9551 17255
rect 9539 17224 10364 17252
rect 9539 17221 9551 17224
rect 9493 17215 9551 17221
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 8846 17144 8852 17196
rect 8904 17184 8910 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8904 17156 9229 17184
rect 8904 17144 8910 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 9309 17187 9367 17193
rect 9309 17153 9321 17187
rect 9355 17153 9367 17187
rect 9583 17187 9641 17193
rect 9583 17184 9595 17187
rect 9309 17147 9367 17153
rect 9508 17156 9595 17184
rect 4798 17116 4804 17128
rect 4264 17088 4804 17116
rect 4798 17076 4804 17088
rect 4856 17076 4862 17128
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17116 5135 17119
rect 5258 17116 5264 17128
rect 5123 17088 5264 17116
rect 5123 17085 5135 17088
rect 5077 17079 5135 17085
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 6454 17076 6460 17128
rect 6512 17116 6518 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6512 17088 6837 17116
rect 6512 17076 6518 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7006 17076 7012 17128
rect 7064 17076 7070 17128
rect 3237 17051 3295 17057
rect 3237 17048 3249 17051
rect 2746 17020 3249 17048
rect 2314 16940 2320 16992
rect 2372 16980 2378 16992
rect 2746 16980 2774 17020
rect 3237 17017 3249 17020
rect 3283 17017 3295 17051
rect 3237 17011 3295 17017
rect 4062 17008 4068 17060
rect 4120 17048 4126 17060
rect 5353 17051 5411 17057
rect 5353 17048 5365 17051
rect 4120 17020 5365 17048
rect 4120 17008 4126 17020
rect 5353 17017 5365 17020
rect 5399 17017 5411 17051
rect 9324 17048 9352 17147
rect 9508 17128 9536 17156
rect 9583 17153 9595 17156
rect 9629 17153 9641 17187
rect 9583 17147 9641 17153
rect 9709 17187 9767 17193
rect 9709 17153 9721 17187
rect 9755 17184 9767 17187
rect 9950 17184 9956 17196
rect 9755 17156 9956 17184
rect 9755 17153 9767 17156
rect 9709 17147 9767 17153
rect 9950 17144 9956 17156
rect 10008 17184 10014 17196
rect 10336 17193 10364 17224
rect 10410 17212 10416 17264
rect 10468 17252 10474 17264
rect 10686 17252 10692 17264
rect 10468 17224 10692 17252
rect 10468 17212 10474 17224
rect 10686 17212 10692 17224
rect 10744 17212 10750 17264
rect 12526 17252 12532 17264
rect 11532 17224 12532 17252
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 10008 17156 10149 17184
rect 10008 17144 10014 17156
rect 10137 17153 10149 17156
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10502 17184 10508 17196
rect 10367 17156 10508 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 11532 17193 11560 17224
rect 12526 17212 12532 17224
rect 12584 17212 12590 17264
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 11793 17187 11851 17193
rect 11793 17153 11805 17187
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 12437 17187 12495 17193
rect 12437 17153 12449 17187
rect 12483 17184 12495 17187
rect 12636 17184 12664 17280
rect 13538 17212 13544 17264
rect 13596 17252 13602 17264
rect 13596 17224 16252 17252
rect 13596 17212 13602 17224
rect 12483 17156 12664 17184
rect 12713 17187 12771 17193
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 12713 17153 12725 17187
rect 12759 17184 12771 17187
rect 12802 17184 12808 17196
rect 12759 17156 12808 17184
rect 12759 17153 12771 17156
rect 12713 17147 12771 17153
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 10229 17119 10287 17125
rect 10229 17116 10241 17119
rect 9548 17088 10241 17116
rect 9548 17076 9554 17088
rect 10229 17085 10241 17088
rect 10275 17085 10287 17119
rect 10229 17079 10287 17085
rect 10413 17119 10471 17125
rect 10413 17085 10425 17119
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 10318 17048 10324 17060
rect 9324 17020 10324 17048
rect 5353 17011 5411 17017
rect 10318 17008 10324 17020
rect 10376 17048 10382 17060
rect 10428 17048 10456 17079
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11238 17116 11244 17128
rect 11112 17088 11244 17116
rect 11112 17076 11118 17088
rect 11238 17076 11244 17088
rect 11296 17116 11302 17128
rect 11808 17116 11836 17147
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 15105 17187 15163 17193
rect 13648 17156 15056 17184
rect 11296 17088 11836 17116
rect 12161 17119 12219 17125
rect 11296 17076 11302 17088
rect 12161 17085 12173 17119
rect 12207 17116 12219 17119
rect 12986 17116 12992 17128
rect 12207 17088 12992 17116
rect 12207 17085 12219 17088
rect 12161 17079 12219 17085
rect 12986 17076 12992 17088
rect 13044 17076 13050 17128
rect 10376 17020 10456 17048
rect 12345 17051 12403 17057
rect 10376 17008 10382 17020
rect 12345 17017 12357 17051
rect 12391 17048 12403 17051
rect 13648 17048 13676 17156
rect 12391 17020 13676 17048
rect 15028 17048 15056 17156
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15120 17116 15148 17147
rect 15378 17144 15384 17196
rect 15436 17144 15442 17196
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 16224 17193 16252 17224
rect 17586 17212 17592 17264
rect 17644 17252 17650 17264
rect 17681 17255 17739 17261
rect 17681 17252 17693 17255
rect 17644 17224 17693 17252
rect 17644 17212 17650 17224
rect 17681 17221 17693 17224
rect 17727 17221 17739 17255
rect 17681 17215 17739 17221
rect 17865 17255 17923 17261
rect 17865 17221 17877 17255
rect 17911 17252 17923 17255
rect 17954 17252 17960 17264
rect 17911 17224 17960 17252
rect 17911 17221 17923 17224
rect 17865 17215 17923 17221
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 21910 17252 21916 17264
rect 19536 17224 21916 17252
rect 16209 17187 16267 17193
rect 15712 17156 16160 17184
rect 15712 17144 15718 17156
rect 16132 17125 16160 17156
rect 16209 17153 16221 17187
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 16298 17144 16304 17196
rect 16356 17144 16362 17196
rect 19536 17193 19564 17224
rect 21910 17212 21916 17224
rect 21968 17212 21974 17264
rect 22020 17224 22232 17252
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17184 19855 17187
rect 19886 17184 19892 17196
rect 19843 17156 19892 17184
rect 19843 17153 19855 17156
rect 19797 17147 19855 17153
rect 19886 17144 19892 17156
rect 19944 17184 19950 17196
rect 20165 17187 20223 17193
rect 19944 17156 20116 17184
rect 19944 17144 19950 17156
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15120 17088 15853 17116
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 16025 17119 16083 17125
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17116 16175 17119
rect 18046 17116 18052 17128
rect 16163 17088 18052 17116
rect 16163 17085 16175 17088
rect 16117 17079 16175 17085
rect 15194 17048 15200 17060
rect 15028 17020 15200 17048
rect 12391 17017 12403 17020
rect 12345 17011 12403 17017
rect 15194 17008 15200 17020
rect 15252 17008 15258 17060
rect 16040 17048 16068 17079
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19392 17088 19717 17116
rect 19392 17076 19398 17088
rect 19705 17085 19717 17088
rect 19751 17116 19763 17119
rect 19981 17119 20039 17125
rect 19981 17116 19993 17119
rect 19751 17088 19993 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 19981 17085 19993 17088
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 16390 17048 16396 17060
rect 16040 17020 16396 17048
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 19613 17051 19671 17057
rect 19613 17017 19625 17051
rect 19659 17048 19671 17051
rect 19886 17048 19892 17060
rect 19659 17020 19892 17048
rect 19659 17017 19671 17020
rect 19613 17011 19671 17017
rect 19886 17008 19892 17020
rect 19944 17008 19950 17060
rect 2372 16952 2774 16980
rect 2372 16940 2378 16952
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 4798 16980 4804 16992
rect 4212 16952 4804 16980
rect 4212 16940 4218 16952
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 9861 16983 9919 16989
rect 9861 16949 9873 16983
rect 9907 16980 9919 16983
rect 10134 16980 10140 16992
rect 9907 16952 10140 16980
rect 9907 16949 9919 16952
rect 9861 16943 9919 16949
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 13872 16952 15117 16980
rect 13872 16940 13878 16952
rect 15105 16949 15117 16952
rect 15151 16949 15163 16983
rect 15105 16943 15163 16949
rect 19334 16940 19340 16992
rect 19392 16940 19398 16992
rect 20088 16980 20116 17156
rect 20165 17153 20177 17187
rect 20211 17184 20223 17187
rect 20990 17184 20996 17196
rect 20211 17156 20996 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 22020 17184 22048 17224
rect 21928 17156 22048 17184
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17116 20499 17119
rect 20714 17116 20720 17128
rect 20487 17088 20720 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 21082 17076 21088 17128
rect 21140 17116 21146 17128
rect 21821 17119 21879 17125
rect 21821 17116 21833 17119
rect 21140 17088 21833 17116
rect 21140 17076 21146 17088
rect 21821 17085 21833 17088
rect 21867 17085 21879 17119
rect 21821 17079 21879 17085
rect 20162 17008 20168 17060
rect 20220 17048 20226 17060
rect 20349 17051 20407 17057
rect 20349 17048 20361 17051
rect 20220 17020 20361 17048
rect 20220 17008 20226 17020
rect 20349 17017 20361 17020
rect 20395 17048 20407 17051
rect 21928 17048 21956 17156
rect 22094 17144 22100 17196
rect 22152 17144 22158 17196
rect 22204 17193 22232 17224
rect 26326 17212 26332 17264
rect 26384 17252 26390 17264
rect 27525 17255 27583 17261
rect 27525 17252 27537 17255
rect 26384 17224 27537 17252
rect 26384 17212 26390 17224
rect 27525 17221 27537 17224
rect 27571 17252 27583 17255
rect 30006 17252 30012 17264
rect 27571 17224 30012 17252
rect 27571 17221 27583 17224
rect 27525 17215 27583 17221
rect 30006 17212 30012 17224
rect 30064 17212 30070 17264
rect 30282 17212 30288 17264
rect 30340 17212 30346 17264
rect 31726 17252 31754 17292
rect 31941 17289 31953 17323
rect 31987 17320 31999 17323
rect 32030 17320 32036 17332
rect 31987 17292 32036 17320
rect 31987 17289 31999 17292
rect 31941 17283 31999 17289
rect 32030 17280 32036 17292
rect 32088 17320 32094 17332
rect 32950 17320 32956 17332
rect 32088 17292 32956 17320
rect 32088 17280 32094 17292
rect 32950 17280 32956 17292
rect 33008 17280 33014 17332
rect 30392 17224 31340 17252
rect 31726 17224 32168 17252
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 22281 17187 22339 17193
rect 22281 17153 22293 17187
rect 22327 17153 22339 17187
rect 22281 17147 22339 17153
rect 22459 17187 22517 17193
rect 22459 17153 22471 17187
rect 22505 17184 22517 17187
rect 22646 17184 22652 17196
rect 22505 17156 22652 17184
rect 22505 17153 22517 17156
rect 22459 17147 22517 17153
rect 22296 17116 22324 17147
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 23382 17144 23388 17196
rect 23440 17144 23446 17196
rect 24394 17144 24400 17196
rect 24452 17184 24458 17196
rect 25130 17184 25136 17196
rect 24452 17156 25136 17184
rect 24452 17144 24458 17156
rect 25130 17144 25136 17156
rect 25188 17144 25194 17196
rect 25225 17187 25283 17193
rect 25225 17153 25237 17187
rect 25271 17184 25283 17187
rect 25314 17184 25320 17196
rect 25271 17156 25320 17184
rect 25271 17153 25283 17156
rect 25225 17147 25283 17153
rect 25314 17144 25320 17156
rect 25372 17144 25378 17196
rect 25409 17187 25467 17193
rect 25409 17153 25421 17187
rect 25455 17184 25467 17187
rect 25498 17184 25504 17196
rect 25455 17156 25504 17184
rect 25455 17153 25467 17156
rect 25409 17147 25467 17153
rect 25498 17144 25504 17156
rect 25556 17144 25562 17196
rect 27338 17144 27344 17196
rect 27396 17144 27402 17196
rect 27614 17144 27620 17196
rect 27672 17144 27678 17196
rect 27709 17187 27767 17193
rect 27709 17153 27721 17187
rect 27755 17184 27767 17187
rect 27798 17184 27804 17196
rect 27755 17156 27804 17184
rect 27755 17153 27767 17156
rect 27709 17147 27767 17153
rect 27798 17144 27804 17156
rect 27856 17144 27862 17196
rect 27982 17144 27988 17196
rect 28040 17144 28046 17196
rect 30190 17144 30196 17196
rect 30248 17184 30254 17196
rect 30392 17184 30420 17224
rect 30248 17156 30420 17184
rect 30248 17144 30254 17156
rect 30558 17144 30564 17196
rect 30616 17144 30622 17196
rect 31312 17193 31340 17224
rect 31478 17193 31484 17196
rect 31297 17187 31355 17193
rect 31297 17153 31309 17187
rect 31343 17153 31355 17187
rect 31297 17147 31355 17153
rect 31445 17187 31484 17193
rect 31445 17153 31457 17187
rect 31445 17147 31484 17153
rect 31478 17144 31484 17147
rect 31536 17144 31542 17196
rect 31573 17187 31631 17193
rect 31573 17153 31585 17187
rect 31619 17153 31631 17187
rect 31573 17147 31631 17153
rect 22554 17116 22560 17128
rect 22296 17088 22560 17116
rect 22554 17076 22560 17088
rect 22612 17076 22618 17128
rect 28810 17076 28816 17128
rect 28868 17076 28874 17128
rect 30469 17119 30527 17125
rect 30469 17085 30481 17119
rect 30515 17085 30527 17119
rect 30469 17079 30527 17085
rect 20395 17020 21956 17048
rect 25317 17051 25375 17057
rect 20395 17017 20407 17020
rect 20349 17011 20407 17017
rect 25317 17017 25329 17051
rect 25363 17048 25375 17051
rect 25958 17048 25964 17060
rect 25363 17020 25964 17048
rect 25363 17017 25375 17020
rect 25317 17011 25375 17017
rect 25958 17008 25964 17020
rect 26016 17008 26022 17060
rect 30484 17048 30512 17079
rect 30650 17076 30656 17128
rect 30708 17116 30714 17128
rect 31202 17116 31208 17128
rect 30708 17088 31208 17116
rect 30708 17076 30714 17088
rect 31202 17076 31208 17088
rect 31260 17116 31266 17128
rect 31588 17116 31616 17147
rect 31662 17144 31668 17196
rect 31720 17144 31726 17196
rect 31846 17193 31852 17196
rect 31803 17187 31852 17193
rect 31803 17153 31815 17187
rect 31849 17153 31852 17187
rect 31803 17147 31852 17153
rect 31846 17144 31852 17147
rect 31904 17144 31910 17196
rect 32140 17193 32168 17224
rect 32125 17187 32183 17193
rect 32125 17153 32137 17187
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 32214 17144 32220 17196
rect 32272 17144 32278 17196
rect 32306 17144 32312 17196
rect 32364 17184 32370 17196
rect 32490 17184 32496 17196
rect 32364 17156 32496 17184
rect 32364 17144 32370 17156
rect 32490 17144 32496 17156
rect 32548 17144 32554 17196
rect 31260 17088 31616 17116
rect 31680 17116 31708 17144
rect 32030 17116 32036 17128
rect 31680 17088 32036 17116
rect 31260 17076 31266 17088
rect 32030 17076 32036 17088
rect 32088 17076 32094 17128
rect 31938 17048 31944 17060
rect 30484 17020 31944 17048
rect 31938 17008 31944 17020
rect 31996 17008 32002 17060
rect 34698 17048 34704 17060
rect 32232 17020 34704 17048
rect 21266 16980 21272 16992
rect 20088 16952 21272 16980
rect 21266 16940 21272 16952
rect 21324 16980 21330 16992
rect 22554 16980 22560 16992
rect 21324 16952 22560 16980
rect 21324 16940 21330 16952
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 27246 16940 27252 16992
rect 27304 16980 27310 16992
rect 28442 16980 28448 16992
rect 27304 16952 28448 16980
rect 27304 16940 27310 16952
rect 28442 16940 28448 16952
rect 28500 16980 28506 16992
rect 29638 16980 29644 16992
rect 28500 16952 29644 16980
rect 28500 16940 28506 16952
rect 29638 16940 29644 16952
rect 29696 16940 29702 16992
rect 29730 16940 29736 16992
rect 29788 16980 29794 16992
rect 32232 16989 32260 17020
rect 34698 17008 34704 17020
rect 34756 17008 34762 17060
rect 30377 16983 30435 16989
rect 30377 16980 30389 16983
rect 29788 16952 30389 16980
rect 29788 16940 29794 16952
rect 30377 16949 30389 16952
rect 30423 16949 30435 16983
rect 30377 16943 30435 16949
rect 32217 16983 32275 16989
rect 32217 16949 32229 16983
rect 32263 16949 32275 16983
rect 32217 16943 32275 16949
rect 32306 16940 32312 16992
rect 32364 16980 32370 16992
rect 32493 16983 32551 16989
rect 32493 16980 32505 16983
rect 32364 16952 32505 16980
rect 32364 16940 32370 16952
rect 32493 16949 32505 16952
rect 32539 16949 32551 16983
rect 32493 16943 32551 16949
rect 1104 16890 36432 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 36432 16890
rect 1104 16816 36432 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1949 16779 2007 16785
rect 1949 16776 1961 16779
rect 1728 16748 1961 16776
rect 1728 16736 1734 16748
rect 1949 16745 1961 16748
rect 1995 16745 2007 16779
rect 1949 16739 2007 16745
rect 3145 16779 3203 16785
rect 3145 16745 3157 16779
rect 3191 16776 3203 16779
rect 3694 16776 3700 16788
rect 3191 16748 3700 16776
rect 3191 16745 3203 16748
rect 3145 16739 3203 16745
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 4430 16736 4436 16788
rect 4488 16776 4494 16788
rect 5718 16776 5724 16788
rect 4488 16748 5724 16776
rect 4488 16736 4494 16748
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 6086 16736 6092 16788
rect 6144 16736 6150 16788
rect 9766 16736 9772 16788
rect 9824 16736 9830 16788
rect 10318 16736 10324 16788
rect 10376 16736 10382 16788
rect 10689 16779 10747 16785
rect 10689 16745 10701 16779
rect 10735 16776 10747 16779
rect 11606 16776 11612 16788
rect 10735 16748 11612 16776
rect 10735 16745 10747 16748
rect 10689 16739 10747 16745
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 12802 16736 12808 16788
rect 12860 16736 12866 16788
rect 20622 16736 20628 16788
rect 20680 16776 20686 16788
rect 20990 16776 20996 16788
rect 20680 16748 20996 16776
rect 20680 16736 20686 16748
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 24397 16779 24455 16785
rect 24397 16776 24409 16779
rect 24084 16748 24409 16776
rect 24084 16736 24090 16748
rect 24397 16745 24409 16748
rect 24443 16745 24455 16779
rect 24397 16739 24455 16745
rect 25222 16736 25228 16788
rect 25280 16776 25286 16788
rect 25590 16776 25596 16788
rect 25280 16748 25596 16776
rect 25280 16736 25286 16748
rect 25590 16736 25596 16748
rect 25648 16736 25654 16788
rect 25869 16779 25927 16785
rect 25869 16745 25881 16779
rect 25915 16776 25927 16779
rect 26234 16776 26240 16788
rect 25915 16748 26240 16776
rect 25915 16745 25927 16748
rect 25869 16739 25927 16745
rect 26234 16736 26240 16748
rect 26292 16736 26298 16788
rect 26326 16736 26332 16788
rect 26384 16776 26390 16788
rect 26973 16779 27031 16785
rect 26973 16776 26985 16779
rect 26384 16748 26985 16776
rect 26384 16736 26390 16748
rect 26973 16745 26985 16748
rect 27019 16745 27031 16779
rect 27614 16776 27620 16788
rect 26973 16739 27031 16745
rect 27080 16748 27620 16776
rect 2222 16668 2228 16720
rect 2280 16708 2286 16720
rect 5902 16708 5908 16720
rect 2280 16680 2452 16708
rect 2280 16668 2286 16680
rect 2424 16652 2452 16680
rect 3896 16680 5908 16708
rect 2406 16600 2412 16652
rect 2464 16600 2470 16652
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16640 2559 16643
rect 2590 16640 2596 16652
rect 2547 16612 2596 16640
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 2590 16600 2596 16612
rect 2648 16600 2654 16652
rect 3896 16640 3924 16680
rect 3712 16612 3924 16640
rect 2314 16532 2320 16584
rect 2372 16532 2378 16584
rect 3326 16532 3332 16584
rect 3384 16532 3390 16584
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 3712 16572 3740 16612
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 4890 16640 4896 16652
rect 4396 16612 4896 16640
rect 4396 16600 4402 16612
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 5092 16640 5120 16680
rect 5001 16612 5120 16640
rect 3651 16544 3740 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 4430 16532 4436 16584
rect 4488 16572 4494 16584
rect 5001 16581 5029 16612
rect 5828 16581 5856 16680
rect 5902 16668 5908 16680
rect 5960 16708 5966 16720
rect 8386 16708 8392 16720
rect 5960 16680 8392 16708
rect 5960 16668 5966 16680
rect 8386 16668 8392 16680
rect 8444 16708 8450 16720
rect 12526 16708 12532 16720
rect 8444 16680 12532 16708
rect 8444 16668 8450 16680
rect 6454 16600 6460 16652
rect 6512 16640 6518 16652
rect 6549 16643 6607 16649
rect 6549 16640 6561 16643
rect 6512 16612 6561 16640
rect 6512 16600 6518 16612
rect 6549 16609 6561 16612
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 6730 16600 6736 16652
rect 6788 16600 6794 16652
rect 9306 16600 9312 16652
rect 9364 16600 9370 16652
rect 4709 16575 4767 16581
rect 4709 16572 4721 16575
rect 4488 16544 4721 16572
rect 4488 16532 4494 16544
rect 4709 16541 4721 16544
rect 4755 16541 4767 16575
rect 4709 16535 4767 16541
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16541 5043 16575
rect 4985 16535 5043 16541
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16541 5503 16575
rect 5445 16535 5503 16541
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16541 5871 16575
rect 7098 16572 7104 16584
rect 5813 16535 5871 16541
rect 6380 16544 7104 16572
rect 3513 16507 3571 16513
rect 3513 16473 3525 16507
rect 3559 16504 3571 16507
rect 3694 16504 3700 16516
rect 3559 16476 3700 16504
rect 3559 16473 3571 16476
rect 3513 16467 3571 16473
rect 3694 16464 3700 16476
rect 3752 16464 3758 16516
rect 4522 16464 4528 16516
rect 4580 16464 4586 16516
rect 4614 16464 4620 16516
rect 4672 16504 4678 16516
rect 5460 16504 5488 16535
rect 4672 16476 5488 16504
rect 4672 16464 4678 16476
rect 5626 16464 5632 16516
rect 5684 16464 5690 16516
rect 5721 16507 5779 16513
rect 5721 16473 5733 16507
rect 5767 16504 5779 16507
rect 6380 16504 6408 16544
rect 7098 16532 7104 16544
rect 7156 16572 7162 16584
rect 7469 16575 7527 16581
rect 7469 16572 7481 16575
rect 7156 16544 7481 16572
rect 7156 16532 7162 16544
rect 7469 16541 7481 16544
rect 7515 16541 7527 16575
rect 7469 16535 7527 16541
rect 8478 16532 8484 16584
rect 8536 16532 8542 16584
rect 8938 16532 8944 16584
rect 8996 16532 9002 16584
rect 9033 16575 9091 16581
rect 9033 16541 9045 16575
rect 9079 16572 9091 16575
rect 9324 16572 9352 16600
rect 9416 16581 9444 16680
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 12710 16668 12716 16720
rect 12768 16668 12774 16720
rect 18874 16668 18880 16720
rect 18932 16708 18938 16720
rect 22002 16708 22008 16720
rect 18932 16680 22008 16708
rect 18932 16668 18938 16680
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 23198 16708 23204 16720
rect 22204 16680 23204 16708
rect 9490 16600 9496 16652
rect 9548 16600 9554 16652
rect 10781 16643 10839 16649
rect 10781 16609 10793 16643
rect 10827 16640 10839 16643
rect 12728 16640 12756 16668
rect 19334 16640 19340 16652
rect 10827 16612 12756 16640
rect 12820 16612 19340 16640
rect 10827 16609 10839 16612
rect 10781 16603 10839 16609
rect 9079 16544 9352 16572
rect 9401 16575 9459 16581
rect 9079 16541 9091 16544
rect 9033 16535 9091 16541
rect 9401 16541 9413 16575
rect 9447 16541 9459 16575
rect 10505 16575 10563 16581
rect 10505 16572 10517 16575
rect 9401 16535 9459 16541
rect 10428 16544 10517 16572
rect 5767 16476 6408 16504
rect 6457 16507 6515 16513
rect 5767 16473 5779 16476
rect 5721 16467 5779 16473
rect 6457 16473 6469 16507
rect 6503 16504 6515 16507
rect 6917 16507 6975 16513
rect 6917 16504 6929 16507
rect 6503 16476 6929 16504
rect 6503 16473 6515 16476
rect 6457 16467 6515 16473
rect 6917 16473 6929 16476
rect 6963 16473 6975 16507
rect 8570 16504 8576 16516
rect 6917 16467 6975 16473
rect 7484 16476 8576 16504
rect 3602 16396 3608 16448
rect 3660 16436 3666 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3660 16408 3801 16436
rect 3660 16396 3666 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 4893 16439 4951 16445
rect 4893 16436 4905 16439
rect 4856 16408 4905 16436
rect 4856 16396 4862 16408
rect 4893 16405 4905 16408
rect 4939 16405 4951 16439
rect 4893 16399 4951 16405
rect 5997 16439 6055 16445
rect 5997 16405 6009 16439
rect 6043 16436 6055 16439
rect 7484 16436 7512 16476
rect 8570 16464 8576 16476
rect 8628 16464 8634 16516
rect 9217 16507 9275 16513
rect 9217 16504 9229 16507
rect 8680 16476 9229 16504
rect 6043 16408 7512 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 7558 16396 7564 16448
rect 7616 16436 7622 16448
rect 7929 16439 7987 16445
rect 7929 16436 7941 16439
rect 7616 16408 7941 16436
rect 7616 16396 7622 16408
rect 7929 16405 7941 16408
rect 7975 16405 7987 16439
rect 7929 16399 7987 16405
rect 8294 16396 8300 16448
rect 8352 16436 8358 16448
rect 8680 16436 8708 16476
rect 9217 16473 9229 16476
rect 9263 16473 9275 16507
rect 9217 16467 9275 16473
rect 9309 16507 9367 16513
rect 9309 16473 9321 16507
rect 9355 16504 9367 16507
rect 9490 16504 9496 16516
rect 9355 16476 9496 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 9490 16464 9496 16476
rect 9548 16464 9554 16516
rect 9674 16464 9680 16516
rect 9732 16464 9738 16516
rect 8352 16408 8708 16436
rect 8352 16396 8358 16408
rect 8938 16396 8944 16448
rect 8996 16436 9002 16448
rect 10428 16436 10456 16544
rect 10505 16541 10517 16544
rect 10551 16572 10563 16575
rect 11054 16572 11060 16584
rect 10551 16544 11060 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 11606 16532 11612 16584
rect 11664 16532 11670 16584
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11808 16581 11836 16612
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 11756 16544 11805 16572
rect 11756 16532 11762 16544
rect 11793 16541 11805 16544
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 12710 16572 12716 16584
rect 12667 16544 12716 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 12820 16581 12848 16612
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 22204 16640 22232 16680
rect 23198 16668 23204 16680
rect 23256 16668 23262 16720
rect 24210 16668 24216 16720
rect 24268 16708 24274 16720
rect 25314 16708 25320 16720
rect 24268 16680 25320 16708
rect 24268 16668 24274 16680
rect 25314 16668 25320 16680
rect 25372 16668 25378 16720
rect 22112 16612 22232 16640
rect 12805 16575 12863 16581
rect 12805 16541 12817 16575
rect 12851 16541 12863 16575
rect 12805 16535 12863 16541
rect 18322 16532 18328 16584
rect 18380 16572 18386 16584
rect 22112 16572 22140 16612
rect 22646 16600 22652 16652
rect 22704 16640 22710 16652
rect 23382 16640 23388 16652
rect 22704 16612 23388 16640
rect 22704 16600 22710 16612
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 24412 16612 25084 16640
rect 18380 16544 22140 16572
rect 18380 16532 18386 16544
rect 22186 16532 22192 16584
rect 22244 16572 22250 16584
rect 23477 16575 23535 16581
rect 23477 16572 23489 16575
rect 22244 16544 23489 16572
rect 22244 16532 22250 16544
rect 23477 16541 23489 16544
rect 23523 16572 23535 16575
rect 23523 16544 23904 16572
rect 23523 16541 23535 16544
rect 23477 16535 23535 16541
rect 10594 16464 10600 16516
rect 10652 16504 10658 16516
rect 10873 16507 10931 16513
rect 10873 16504 10885 16507
rect 10652 16476 10885 16504
rect 10652 16464 10658 16476
rect 10873 16473 10885 16476
rect 10919 16473 10931 16507
rect 11624 16504 11652 16532
rect 13538 16504 13544 16516
rect 11624 16476 13544 16504
rect 10873 16467 10931 16473
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 14182 16464 14188 16516
rect 14240 16504 14246 16516
rect 15654 16504 15660 16516
rect 14240 16476 15660 16504
rect 14240 16464 14246 16476
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 18046 16464 18052 16516
rect 18104 16504 18110 16516
rect 21634 16504 21640 16516
rect 18104 16476 21640 16504
rect 18104 16464 18110 16476
rect 21634 16464 21640 16476
rect 21692 16464 21698 16516
rect 8996 16408 10456 16436
rect 8996 16396 9002 16408
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 23106 16436 23112 16448
rect 12124 16408 23112 16436
rect 12124 16396 12130 16408
rect 23106 16396 23112 16408
rect 23164 16396 23170 16448
rect 23876 16436 23904 16544
rect 23934 16532 23940 16584
rect 23992 16572 23998 16584
rect 24412 16572 24440 16612
rect 23992 16544 24440 16572
rect 23992 16532 23998 16544
rect 24486 16532 24492 16584
rect 24544 16581 24550 16584
rect 24544 16575 24593 16581
rect 24544 16541 24547 16575
rect 24581 16541 24593 16575
rect 24544 16535 24593 16541
rect 24544 16532 24550 16535
rect 24854 16532 24860 16584
rect 24912 16581 24918 16584
rect 25056 16581 25084 16612
rect 25130 16600 25136 16652
rect 25188 16640 25194 16652
rect 26329 16643 26387 16649
rect 26329 16640 26341 16643
rect 25188 16612 26341 16640
rect 25188 16600 25194 16612
rect 26329 16609 26341 16612
rect 26375 16609 26387 16643
rect 27080 16640 27108 16748
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 28810 16736 28816 16788
rect 28868 16776 28874 16788
rect 34054 16776 34060 16788
rect 28868 16748 34060 16776
rect 28868 16736 28874 16748
rect 27154 16708 27160 16720
rect 26329 16603 26387 16609
rect 26436 16612 27108 16640
rect 27148 16668 27160 16708
rect 27212 16668 27218 16720
rect 27430 16668 27436 16720
rect 27488 16668 27494 16720
rect 24912 16575 24951 16581
rect 24939 16541 24951 16575
rect 24912 16535 24951 16541
rect 25041 16575 25099 16581
rect 25041 16541 25053 16575
rect 25087 16541 25099 16575
rect 25041 16535 25099 16541
rect 24912 16532 24918 16535
rect 25222 16532 25228 16584
rect 25280 16572 25286 16584
rect 25501 16575 25559 16581
rect 25501 16572 25513 16575
rect 25280 16544 25513 16572
rect 25280 16532 25286 16544
rect 25501 16541 25513 16544
rect 25547 16541 25559 16575
rect 25501 16535 25559 16541
rect 25682 16532 25688 16584
rect 25740 16532 25746 16584
rect 25961 16575 26019 16581
rect 25961 16541 25973 16575
rect 26007 16572 26019 16575
rect 26436 16572 26464 16612
rect 26007 16544 26464 16572
rect 26007 16541 26019 16544
rect 25961 16535 26019 16541
rect 26510 16532 26516 16584
rect 26568 16532 26574 16584
rect 26602 16532 26608 16584
rect 26660 16532 26666 16584
rect 26786 16532 26792 16584
rect 26844 16532 26850 16584
rect 26881 16575 26939 16581
rect 26881 16541 26893 16575
rect 26927 16572 26939 16575
rect 26970 16572 26976 16584
rect 26927 16544 26976 16572
rect 26927 16541 26939 16544
rect 26881 16535 26939 16541
rect 26970 16532 26976 16544
rect 27028 16532 27034 16584
rect 27148 16582 27176 16668
rect 27448 16640 27476 16668
rect 27614 16640 27620 16652
rect 27264 16612 27620 16640
rect 27148 16581 27200 16582
rect 27264 16581 27292 16612
rect 27614 16600 27620 16612
rect 27672 16600 27678 16652
rect 32048 16649 32076 16748
rect 34054 16736 34060 16748
rect 34112 16736 34118 16788
rect 32033 16643 32091 16649
rect 32033 16609 32045 16643
rect 32079 16609 32091 16643
rect 32033 16603 32091 16609
rect 32306 16600 32312 16652
rect 32364 16600 32370 16652
rect 35161 16643 35219 16649
rect 35161 16609 35173 16643
rect 35207 16640 35219 16643
rect 35250 16640 35256 16652
rect 35207 16612 35256 16640
rect 35207 16609 35219 16612
rect 35161 16603 35219 16609
rect 35250 16600 35256 16612
rect 35308 16600 35314 16652
rect 27148 16575 27215 16581
rect 27148 16554 27169 16575
rect 27157 16541 27169 16554
rect 27203 16541 27215 16575
rect 27157 16535 27215 16541
rect 27249 16575 27307 16581
rect 27249 16541 27261 16575
rect 27295 16541 27307 16575
rect 27249 16535 27307 16541
rect 27430 16532 27436 16584
rect 27488 16572 27494 16584
rect 27525 16575 27583 16581
rect 27525 16572 27537 16575
rect 27488 16544 27537 16572
rect 27488 16532 27494 16544
rect 27525 16541 27537 16544
rect 27571 16541 27583 16575
rect 29178 16572 29184 16584
rect 27525 16535 27583 16541
rect 27632 16544 29184 16572
rect 24670 16464 24676 16516
rect 24728 16464 24734 16516
rect 24765 16507 24823 16513
rect 24765 16473 24777 16507
rect 24811 16504 24823 16507
rect 26326 16504 26332 16516
rect 24811 16476 26332 16504
rect 24811 16473 24823 16476
rect 24765 16467 24823 16473
rect 26326 16464 26332 16476
rect 26384 16464 26390 16516
rect 26528 16504 26556 16532
rect 27341 16507 27399 16513
rect 27341 16504 27353 16507
rect 26528 16476 27353 16504
rect 27341 16473 27353 16476
rect 27387 16504 27399 16507
rect 27632 16504 27660 16544
rect 29178 16532 29184 16544
rect 29236 16532 29242 16584
rect 33870 16532 33876 16584
rect 33928 16572 33934 16584
rect 34057 16575 34115 16581
rect 34057 16572 34069 16575
rect 33928 16544 34069 16572
rect 33928 16532 33934 16544
rect 34057 16541 34069 16544
rect 34103 16541 34115 16575
rect 34057 16535 34115 16541
rect 35529 16575 35587 16581
rect 35529 16541 35541 16575
rect 35575 16572 35587 16575
rect 36078 16572 36084 16584
rect 35575 16544 36084 16572
rect 35575 16541 35587 16544
rect 35529 16535 35587 16541
rect 36078 16532 36084 16544
rect 36136 16532 36142 16584
rect 27387 16476 27660 16504
rect 28169 16507 28227 16513
rect 27387 16473 27399 16476
rect 27341 16467 27399 16473
rect 28169 16473 28181 16507
rect 28215 16473 28227 16507
rect 28169 16467 28227 16473
rect 27982 16436 27988 16448
rect 23876 16408 27988 16436
rect 27982 16396 27988 16408
rect 28040 16436 28046 16448
rect 28184 16436 28212 16467
rect 28258 16464 28264 16516
rect 28316 16504 28322 16516
rect 28905 16507 28963 16513
rect 28905 16504 28917 16507
rect 28316 16476 28917 16504
rect 28316 16464 28322 16476
rect 28905 16473 28917 16476
rect 28951 16473 28963 16507
rect 28905 16467 28963 16473
rect 30374 16464 30380 16516
rect 30432 16504 30438 16516
rect 31294 16504 31300 16516
rect 30432 16476 31300 16504
rect 30432 16464 30438 16476
rect 31294 16464 31300 16476
rect 31352 16464 31358 16516
rect 33594 16504 33600 16516
rect 33534 16476 33600 16504
rect 33594 16464 33600 16476
rect 33652 16464 33658 16516
rect 28040 16408 28212 16436
rect 28040 16396 28046 16408
rect 1104 16346 36432 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 36432 16346
rect 1104 16272 36432 16294
rect 3145 16235 3203 16241
rect 3145 16201 3157 16235
rect 3191 16201 3203 16235
rect 3145 16195 3203 16201
rect 3160 16164 3188 16195
rect 3602 16192 3608 16244
rect 3660 16192 3666 16244
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 3878 16232 3884 16244
rect 3743 16204 3884 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 3878 16192 3884 16204
rect 3936 16192 3942 16244
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 4939 16204 5365 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 5353 16195 5411 16201
rect 8205 16235 8263 16241
rect 8205 16201 8217 16235
rect 8251 16232 8263 16235
rect 8478 16232 8484 16244
rect 8251 16204 8484 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 8662 16192 8668 16244
rect 8720 16232 8726 16244
rect 9030 16232 9036 16244
rect 8720 16204 9036 16232
rect 8720 16192 8726 16204
rect 9030 16192 9036 16204
rect 9088 16192 9094 16244
rect 9674 16192 9680 16244
rect 9732 16192 9738 16244
rect 11330 16192 11336 16244
rect 11388 16192 11394 16244
rect 12986 16192 12992 16244
rect 13044 16232 13050 16244
rect 13044 16204 15332 16232
rect 13044 16192 13050 16204
rect 4338 16164 4344 16176
rect 3160 16136 4344 16164
rect 4338 16124 4344 16136
rect 4396 16124 4402 16176
rect 6730 16164 6736 16176
rect 5184 16136 6736 16164
rect 1394 16056 1400 16108
rect 1452 16056 1458 16108
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 4890 16096 4896 16108
rect 2832 16068 4896 16096
rect 2832 16056 2838 16068
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 1719 16000 2774 16028
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 2746 15960 2774 16000
rect 3878 15988 3884 16040
rect 3936 15988 3942 16040
rect 4985 16031 5043 16037
rect 4985 16028 4997 16031
rect 3988 16000 4997 16028
rect 3237 15963 3295 15969
rect 3237 15960 3249 15963
rect 2746 15932 3249 15960
rect 3237 15929 3249 15932
rect 3283 15929 3295 15963
rect 3237 15923 3295 15929
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 3988 15892 4016 16000
rect 4985 15997 4997 16000
rect 5031 15997 5043 16031
rect 4985 15991 5043 15997
rect 5000 15960 5028 15991
rect 5074 15988 5080 16040
rect 5132 16028 5138 16040
rect 5184 16037 5212 16136
rect 6730 16124 6736 16136
rect 6788 16124 6794 16176
rect 9692 16164 9720 16192
rect 7958 16150 9720 16164
rect 7944 16136 9720 16150
rect 5350 16056 5356 16108
rect 5408 16096 5414 16108
rect 6457 16099 6515 16105
rect 6457 16096 6469 16099
rect 5408 16068 6469 16096
rect 5408 16056 5414 16068
rect 6457 16065 6469 16068
rect 6503 16065 6515 16099
rect 6457 16059 6515 16065
rect 5169 16031 5227 16037
rect 5169 16028 5181 16031
rect 5132 16000 5181 16028
rect 5132 15988 5138 16000
rect 5169 15997 5181 16000
rect 5215 15997 5227 16031
rect 5169 15991 5227 15997
rect 5534 15988 5540 16040
rect 5592 16028 5598 16040
rect 5810 16028 5816 16040
rect 5592 16000 5816 16028
rect 5592 15988 5598 16000
rect 5810 15988 5816 16000
rect 5868 16028 5874 16040
rect 5905 16031 5963 16037
rect 5905 16028 5917 16031
rect 5868 16000 5917 16028
rect 5868 15988 5874 16000
rect 5905 15997 5917 16000
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 6733 16031 6791 16037
rect 6733 15997 6745 16031
rect 6779 16028 6791 16031
rect 7190 16028 7196 16040
rect 6779 16000 7196 16028
rect 6779 15997 6791 16000
rect 6733 15991 6791 15997
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 5718 15960 5724 15972
rect 5000 15932 5724 15960
rect 5718 15920 5724 15932
rect 5776 15920 5782 15972
rect 2464 15864 4016 15892
rect 2464 15852 2470 15864
rect 4062 15852 4068 15904
rect 4120 15892 4126 15904
rect 4525 15895 4583 15901
rect 4525 15892 4537 15895
rect 4120 15864 4537 15892
rect 4120 15852 4126 15864
rect 4525 15861 4537 15864
rect 4571 15861 4583 15895
rect 4525 15855 4583 15861
rect 5442 15852 5448 15904
rect 5500 15892 5506 15904
rect 7944 15892 7972 16136
rect 12250 16124 12256 16176
rect 12308 16124 12314 16176
rect 13004 16164 13032 16192
rect 13814 16164 13820 16176
rect 13004 16136 13124 16164
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16096 8999 16099
rect 9306 16096 9312 16108
rect 8987 16068 9312 16096
rect 8987 16065 8999 16068
rect 8941 16059 8999 16065
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 10962 16056 10968 16108
rect 11020 16056 11026 16108
rect 11698 16056 11704 16108
rect 11756 16056 11762 16108
rect 12066 16056 12072 16108
rect 12124 16056 12130 16108
rect 12434 16056 12440 16108
rect 12492 16096 12498 16108
rect 12713 16099 12771 16105
rect 12713 16096 12725 16099
rect 12492 16068 12725 16096
rect 12492 16056 12498 16068
rect 12713 16065 12725 16068
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 12897 16099 12955 16105
rect 12897 16096 12909 16099
rect 12860 16068 12909 16096
rect 12860 16056 12866 16068
rect 12897 16065 12909 16068
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 13096 16094 13124 16136
rect 13372 16136 13820 16164
rect 13372 16105 13400 16136
rect 13814 16124 13820 16136
rect 13872 16124 13878 16176
rect 14829 16167 14887 16173
rect 14829 16164 14841 16167
rect 14108 16136 14841 16164
rect 13173 16099 13231 16105
rect 13173 16094 13185 16099
rect 13096 16066 13185 16094
rect 12989 16059 13047 16065
rect 13173 16065 13185 16066
rect 13219 16065 13231 16099
rect 13173 16059 13231 16065
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 9217 16031 9275 16037
rect 9217 15997 9229 16031
rect 9263 16028 9275 16031
rect 9263 16000 9339 16028
rect 9263 15997 9275 16000
rect 9217 15991 9275 15997
rect 5500 15864 7972 15892
rect 5500 15852 5506 15864
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 8573 15895 8631 15901
rect 8573 15892 8585 15895
rect 8168 15864 8585 15892
rect 8168 15852 8174 15864
rect 8573 15861 8585 15864
rect 8619 15861 8631 15895
rect 8573 15855 8631 15861
rect 8754 15852 8760 15904
rect 8812 15892 8818 15904
rect 9311 15892 9339 16000
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 9861 16031 9919 16037
rect 9861 15997 9873 16031
rect 9907 16028 9919 16031
rect 10594 16028 10600 16040
rect 9907 16000 10600 16028
rect 9907 15997 9919 16000
rect 9861 15991 9919 15997
rect 10594 15988 10600 16000
rect 10652 15988 10658 16040
rect 12802 15920 12808 15972
rect 12860 15920 12866 15972
rect 13004 15960 13032 16059
rect 13538 16056 13544 16108
rect 13596 16096 13602 16108
rect 14007 16099 14065 16105
rect 14007 16096 14019 16099
rect 13596 16068 14019 16096
rect 13596 16056 13602 16068
rect 14007 16065 14019 16068
rect 14053 16096 14065 16099
rect 14108 16096 14136 16136
rect 14829 16133 14841 16136
rect 14875 16133 14887 16167
rect 15304 16164 15332 16204
rect 17126 16192 17132 16244
rect 17184 16192 17190 16244
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 19610 16232 19616 16244
rect 19392 16204 19616 16232
rect 19392 16192 19398 16204
rect 19610 16192 19616 16204
rect 19668 16232 19674 16244
rect 24581 16235 24639 16241
rect 19668 16204 24348 16232
rect 19668 16192 19674 16204
rect 24320 16176 24348 16204
rect 24581 16201 24593 16235
rect 24627 16201 24639 16235
rect 24581 16195 24639 16201
rect 17218 16164 17224 16176
rect 15304 16136 17224 16164
rect 14829 16127 14887 16133
rect 17218 16124 17224 16136
rect 17276 16164 17282 16176
rect 21634 16164 21640 16176
rect 17276 16136 21640 16164
rect 17276 16124 17282 16136
rect 21634 16124 21640 16136
rect 21692 16124 21698 16176
rect 21836 16136 22554 16164
rect 14053 16068 14136 16096
rect 14053 16065 14065 16068
rect 14007 16059 14065 16065
rect 14182 16056 14188 16108
rect 14240 16056 14246 16108
rect 14461 16099 14519 16105
rect 14461 16065 14473 16099
rect 14507 16096 14519 16099
rect 14645 16099 14703 16105
rect 14507 16068 14596 16096
rect 14507 16065 14519 16068
rect 14461 16059 14519 16065
rect 13262 15988 13268 16040
rect 13320 15988 13326 16040
rect 14366 15960 14372 15972
rect 13004 15932 14372 15960
rect 14366 15920 14372 15932
rect 14424 15920 14430 15972
rect 11238 15892 11244 15904
rect 8812 15864 11244 15892
rect 8812 15852 8818 15864
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 12529 15895 12587 15901
rect 12529 15861 12541 15895
rect 12575 15892 12587 15895
rect 13630 15892 13636 15904
rect 12575 15864 13636 15892
rect 12575 15861 12587 15864
rect 12529 15855 12587 15861
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15892 14151 15895
rect 14182 15892 14188 15904
rect 14139 15864 14188 15892
rect 14139 15861 14151 15864
rect 14093 15855 14151 15861
rect 14182 15852 14188 15864
rect 14240 15852 14246 15904
rect 14277 15895 14335 15901
rect 14277 15861 14289 15895
rect 14323 15892 14335 15895
rect 14458 15892 14464 15904
rect 14323 15864 14464 15892
rect 14323 15861 14335 15864
rect 14277 15855 14335 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 14568 15892 14596 16068
rect 14645 16065 14657 16099
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 14660 15960 14688 16059
rect 14752 16028 14780 16059
rect 14918 16056 14924 16108
rect 14976 16056 14982 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15470 16096 15476 16108
rect 15243 16068 15476 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15212 16028 15240 16059
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 17313 16099 17371 16105
rect 17313 16096 17325 16099
rect 17236 16068 17325 16096
rect 17236 16040 17264 16068
rect 17313 16065 17325 16068
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 17586 16056 17592 16108
rect 17644 16056 17650 16108
rect 14752 16000 15240 16028
rect 17218 15988 17224 16040
rect 17276 15988 17282 16040
rect 18690 15988 18696 16040
rect 18748 16028 18754 16040
rect 19886 16028 19892 16040
rect 18748 16000 19892 16028
rect 18748 15988 18754 16000
rect 19886 15988 19892 16000
rect 19944 16028 19950 16040
rect 21542 16028 21548 16040
rect 19944 16000 21548 16028
rect 19944 15988 19950 16000
rect 21542 15988 21548 16000
rect 21600 15988 21606 16040
rect 16942 15960 16948 15972
rect 14660 15932 16948 15960
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 17405 15963 17463 15969
rect 17405 15929 17417 15963
rect 17451 15929 17463 15963
rect 17405 15923 17463 15929
rect 17497 15963 17555 15969
rect 17497 15929 17509 15963
rect 17543 15960 17555 15963
rect 19150 15960 19156 15972
rect 17543 15932 19156 15960
rect 17543 15929 17555 15932
rect 17497 15923 17555 15929
rect 15194 15892 15200 15904
rect 14568 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 15930 15852 15936 15904
rect 15988 15892 15994 15904
rect 17420 15892 17448 15923
rect 19150 15920 19156 15932
rect 19208 15920 19214 15972
rect 19058 15892 19064 15904
rect 15988 15864 19064 15892
rect 15988 15852 15994 15864
rect 19058 15852 19064 15864
rect 19116 15892 19122 15904
rect 20530 15892 20536 15904
rect 19116 15864 20536 15892
rect 19116 15852 19122 15864
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 21836 15901 21864 16136
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21968 16068 22017 16096
rect 21968 16056 21974 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 22278 16056 22284 16108
rect 22336 16056 22342 16108
rect 22526 16105 22554 16136
rect 23658 16124 23664 16176
rect 23716 16164 23722 16176
rect 24210 16164 24216 16176
rect 23716 16136 24216 16164
rect 23716 16124 23722 16136
rect 24210 16124 24216 16136
rect 24268 16124 24274 16176
rect 24302 16124 24308 16176
rect 24360 16124 24366 16176
rect 24596 16164 24624 16195
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 25682 16232 25688 16244
rect 25004 16204 25688 16232
rect 25004 16192 25010 16204
rect 25682 16192 25688 16204
rect 25740 16192 25746 16244
rect 29549 16235 29607 16241
rect 29549 16201 29561 16235
rect 29595 16232 29607 16235
rect 29730 16232 29736 16244
rect 29595 16204 29736 16232
rect 29595 16201 29607 16204
rect 29549 16195 29607 16201
rect 29730 16192 29736 16204
rect 29788 16192 29794 16244
rect 32030 16192 32036 16244
rect 32088 16232 32094 16244
rect 32582 16232 32588 16244
rect 32088 16204 32588 16232
rect 32088 16192 32094 16204
rect 32582 16192 32588 16204
rect 32640 16192 32646 16244
rect 33410 16192 33416 16244
rect 33468 16232 33474 16244
rect 33468 16204 34928 16232
rect 33468 16192 33474 16204
rect 25869 16167 25927 16173
rect 24596 16136 25176 16164
rect 22511 16099 22569 16105
rect 22511 16065 22523 16099
rect 22557 16065 22569 16099
rect 22511 16059 22569 16065
rect 22695 16099 22753 16105
rect 22695 16065 22707 16099
rect 22741 16096 22753 16099
rect 22741 16068 23904 16096
rect 22741 16065 22753 16068
rect 22695 16059 22753 16065
rect 22094 16028 22100 16040
rect 22020 16000 22100 16028
rect 22020 15901 22048 16000
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 22186 15988 22192 16040
rect 22244 15988 22250 16040
rect 22833 16031 22891 16037
rect 22833 16028 22845 16031
rect 22664 16000 22845 16028
rect 22664 15972 22692 16000
rect 22833 15997 22845 16000
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 16028 23443 16031
rect 23474 16028 23480 16040
rect 23431 16000 23480 16028
rect 23431 15997 23443 16000
rect 23385 15991 23443 15997
rect 23474 15988 23480 16000
rect 23532 15988 23538 16040
rect 23876 16028 23904 16068
rect 23934 16056 23940 16108
rect 23992 16056 23998 16108
rect 24026 16056 24032 16108
rect 24084 16096 24090 16108
rect 24443 16099 24501 16105
rect 24084 16068 24129 16096
rect 24084 16056 24090 16068
rect 24443 16065 24455 16099
rect 24489 16096 24501 16099
rect 24578 16096 24584 16108
rect 24489 16068 24584 16096
rect 24489 16065 24501 16068
rect 24443 16059 24501 16065
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 24762 16056 24768 16108
rect 24820 16096 24826 16108
rect 24857 16099 24915 16105
rect 24857 16096 24869 16099
rect 24820 16068 24869 16096
rect 24820 16056 24826 16068
rect 24857 16065 24869 16068
rect 24903 16065 24915 16099
rect 24857 16059 24915 16065
rect 24946 16056 24952 16108
rect 25004 16056 25010 16108
rect 25148 16105 25176 16136
rect 25869 16133 25881 16167
rect 25915 16164 25927 16167
rect 26326 16164 26332 16176
rect 25915 16136 26332 16164
rect 25915 16133 25927 16136
rect 25869 16127 25927 16133
rect 26326 16124 26332 16136
rect 26384 16124 26390 16176
rect 27985 16167 28043 16173
rect 27985 16133 27997 16167
rect 28031 16164 28043 16167
rect 29181 16167 29239 16173
rect 29181 16164 29193 16167
rect 28031 16136 29193 16164
rect 28031 16133 28043 16136
rect 27985 16127 28043 16133
rect 29181 16133 29193 16136
rect 29227 16164 29239 16167
rect 30466 16164 30472 16176
rect 29227 16136 30472 16164
rect 29227 16133 29239 16136
rect 29181 16127 29239 16133
rect 30466 16124 30472 16136
rect 30524 16124 30530 16176
rect 31478 16124 31484 16176
rect 31536 16164 31542 16176
rect 34900 16173 34928 16204
rect 34885 16167 34943 16173
rect 31536 16136 34652 16164
rect 31536 16124 31542 16136
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 25222 16056 25228 16108
rect 25280 16056 25286 16108
rect 26050 16056 26056 16108
rect 26108 16056 26114 16108
rect 27890 16056 27896 16108
rect 27948 16056 27954 16108
rect 28074 16056 28080 16108
rect 28132 16056 28138 16108
rect 28258 16056 28264 16108
rect 28316 16056 28322 16108
rect 28997 16099 29055 16105
rect 28997 16065 29009 16099
rect 29043 16065 29055 16099
rect 28997 16059 29055 16065
rect 26142 16028 26148 16040
rect 23876 16000 26148 16028
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 29012 16028 29040 16059
rect 29270 16056 29276 16108
rect 29328 16056 29334 16108
rect 29365 16099 29423 16105
rect 29365 16065 29377 16099
rect 29411 16096 29423 16099
rect 29454 16096 29460 16108
rect 29411 16068 29460 16096
rect 29411 16065 29423 16068
rect 29365 16059 29423 16065
rect 29454 16056 29460 16068
rect 29512 16056 29518 16108
rect 31018 16056 31024 16108
rect 31076 16096 31082 16108
rect 31205 16099 31263 16105
rect 31205 16096 31217 16099
rect 31076 16068 31217 16096
rect 31076 16056 31082 16068
rect 31205 16065 31217 16068
rect 31251 16065 31263 16099
rect 31205 16059 31263 16065
rect 31389 16099 31447 16105
rect 31389 16065 31401 16099
rect 31435 16096 31447 16099
rect 31754 16096 31760 16108
rect 31435 16068 31760 16096
rect 31435 16065 31447 16068
rect 31389 16059 31447 16065
rect 30098 16028 30104 16040
rect 29012 16000 30104 16028
rect 29380 15972 29408 16000
rect 30098 15988 30104 16000
rect 30156 15988 30162 16040
rect 31220 16028 31248 16059
rect 31754 16056 31760 16068
rect 31812 16056 31818 16108
rect 34624 16105 34652 16136
rect 34885 16133 34897 16167
rect 34931 16133 34943 16167
rect 34885 16127 34943 16133
rect 34609 16099 34667 16105
rect 34609 16065 34621 16099
rect 34655 16065 34667 16099
rect 34609 16059 34667 16065
rect 34793 16099 34851 16105
rect 34793 16065 34805 16099
rect 34839 16065 34851 16099
rect 34793 16059 34851 16065
rect 34977 16099 35035 16105
rect 34977 16065 34989 16099
rect 35023 16065 35035 16099
rect 34977 16059 35035 16065
rect 31478 16028 31484 16040
rect 31220 16000 31484 16028
rect 31478 15988 31484 16000
rect 31536 15988 31542 16040
rect 31570 15988 31576 16040
rect 31628 16028 31634 16040
rect 34808 16028 34836 16059
rect 31628 16000 34836 16028
rect 31628 15988 31634 16000
rect 22646 15920 22652 15972
rect 22704 15920 22710 15972
rect 29362 15920 29368 15972
rect 29420 15920 29426 15972
rect 31662 15960 31668 15972
rect 31588 15932 31668 15960
rect 21821 15895 21879 15901
rect 21821 15861 21833 15895
rect 21867 15861 21879 15895
rect 21821 15855 21879 15861
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15861 22063 15895
rect 22005 15855 22063 15861
rect 23014 15852 23020 15904
rect 23072 15892 23078 15904
rect 24673 15895 24731 15901
rect 24673 15892 24685 15895
rect 23072 15864 24685 15892
rect 23072 15852 23078 15864
rect 24673 15861 24685 15864
rect 24719 15861 24731 15895
rect 24673 15855 24731 15861
rect 25314 15852 25320 15904
rect 25372 15892 25378 15904
rect 25685 15895 25743 15901
rect 25685 15892 25697 15895
rect 25372 15864 25697 15892
rect 25372 15852 25378 15864
rect 25685 15861 25697 15864
rect 25731 15861 25743 15895
rect 25685 15855 25743 15861
rect 27614 15852 27620 15904
rect 27672 15892 27678 15904
rect 30742 15892 30748 15904
rect 27672 15864 30748 15892
rect 27672 15852 27678 15864
rect 30742 15852 30748 15864
rect 30800 15892 30806 15904
rect 30929 15895 30987 15901
rect 30929 15892 30941 15895
rect 30800 15864 30941 15892
rect 30800 15852 30806 15864
rect 30929 15861 30941 15864
rect 30975 15861 30987 15895
rect 30929 15855 30987 15861
rect 31018 15852 31024 15904
rect 31076 15892 31082 15904
rect 31588 15901 31616 15932
rect 31662 15920 31668 15932
rect 31720 15960 31726 15972
rect 34992 15960 35020 16059
rect 31720 15932 35020 15960
rect 31720 15920 31726 15932
rect 31573 15895 31631 15901
rect 31573 15892 31585 15895
rect 31076 15864 31585 15892
rect 31076 15852 31082 15864
rect 31573 15861 31585 15864
rect 31619 15861 31631 15895
rect 31573 15855 31631 15861
rect 34790 15852 34796 15904
rect 34848 15892 34854 15904
rect 35161 15895 35219 15901
rect 35161 15892 35173 15895
rect 34848 15864 35173 15892
rect 34848 15852 34854 15864
rect 35161 15861 35173 15864
rect 35207 15861 35219 15895
rect 35161 15855 35219 15861
rect 1104 15802 36432 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 36432 15802
rect 1104 15728 36432 15750
rect 3605 15691 3663 15697
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 4798 15688 4804 15700
rect 3651 15660 4804 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 4798 15648 4804 15660
rect 4856 15688 4862 15700
rect 4856 15660 5212 15688
rect 4856 15648 4862 15660
rect 3789 15623 3847 15629
rect 3789 15589 3801 15623
rect 3835 15589 3847 15623
rect 3789 15583 3847 15589
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 1854 15552 1860 15564
rect 1452 15524 1860 15552
rect 1452 15512 1458 15524
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 3804 15552 3832 15583
rect 2179 15524 3832 15552
rect 4433 15555 4491 15561
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 5074 15552 5080 15564
rect 4479 15524 5080 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 5184 15561 5212 15660
rect 5442 15648 5448 15700
rect 5500 15648 5506 15700
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 5684 15660 6679 15688
rect 5684 15648 5690 15660
rect 5460 15620 5488 15648
rect 5276 15592 5488 15620
rect 5169 15555 5227 15561
rect 5169 15521 5181 15555
rect 5215 15521 5227 15555
rect 5169 15515 5227 15521
rect 3234 15444 3240 15496
rect 3292 15484 3298 15496
rect 5276 15484 5304 15592
rect 5350 15512 5356 15564
rect 5408 15512 5414 15564
rect 5629 15555 5687 15561
rect 5629 15521 5641 15555
rect 5675 15552 5687 15555
rect 6086 15552 6092 15564
rect 5675 15524 6092 15552
rect 5675 15521 5687 15524
rect 5629 15515 5687 15521
rect 6086 15512 6092 15524
rect 6144 15512 6150 15564
rect 6651 15552 6679 15660
rect 7098 15648 7104 15700
rect 7156 15648 7162 15700
rect 7190 15648 7196 15700
rect 7248 15648 7254 15700
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8202 15688 8208 15700
rect 8067 15660 8208 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 9306 15648 9312 15700
rect 9364 15648 9370 15700
rect 10594 15648 10600 15700
rect 10652 15648 10658 15700
rect 16022 15648 16028 15700
rect 16080 15688 16086 15700
rect 16485 15691 16543 15697
rect 16485 15688 16497 15691
rect 16080 15660 16497 15688
rect 16080 15648 16086 15660
rect 16485 15657 16497 15660
rect 16531 15657 16543 15691
rect 19337 15691 19395 15697
rect 19337 15688 19349 15691
rect 16485 15651 16543 15657
rect 18340 15660 19349 15688
rect 6730 15580 6736 15632
rect 6788 15620 6794 15632
rect 8754 15620 8760 15632
rect 6788 15592 8760 15620
rect 6788 15580 6794 15592
rect 7852 15561 7880 15592
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9122 15580 9128 15632
rect 9180 15620 9186 15632
rect 12437 15623 12495 15629
rect 12437 15620 12449 15623
rect 9180 15592 12449 15620
rect 9180 15580 9186 15592
rect 12437 15589 12449 15592
rect 12483 15589 12495 15623
rect 12437 15583 12495 15589
rect 12802 15580 12808 15632
rect 12860 15620 12866 15632
rect 12860 15592 12940 15620
rect 12860 15580 12866 15592
rect 7837 15555 7895 15561
rect 6651 15524 6955 15552
rect 3292 15456 5304 15484
rect 3292 15444 3298 15456
rect 4157 15419 4215 15425
rect 4157 15385 4169 15419
rect 4203 15416 4215 15419
rect 4617 15419 4675 15425
rect 4617 15416 4629 15419
rect 4203 15388 4629 15416
rect 4203 15385 4215 15388
rect 4157 15379 4215 15385
rect 4617 15385 4629 15388
rect 4663 15385 4675 15419
rect 4617 15379 4675 15385
rect 4798 15376 4804 15428
rect 4856 15416 4862 15428
rect 4856 15388 6118 15416
rect 4856 15376 4862 15388
rect 2130 15308 2136 15360
rect 2188 15348 2194 15360
rect 4249 15351 4307 15357
rect 4249 15348 4261 15351
rect 2188 15320 4261 15348
rect 2188 15308 2194 15320
rect 4249 15317 4261 15320
rect 4295 15348 4307 15351
rect 5258 15348 5264 15360
rect 4295 15320 5264 15348
rect 4295 15317 4307 15320
rect 4249 15311 4307 15317
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 6028 15348 6056 15388
rect 6638 15348 6644 15360
rect 6028 15320 6644 15348
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 6927 15348 6955 15524
rect 7837 15521 7849 15555
rect 7883 15521 7895 15555
rect 8386 15552 8392 15564
rect 7837 15515 7895 15521
rect 8220 15524 8392 15552
rect 7558 15444 7564 15496
rect 7616 15444 7622 15496
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15484 7711 15487
rect 8018 15484 8024 15496
rect 7699 15456 8024 15484
rect 7699 15453 7711 15456
rect 7653 15447 7711 15453
rect 7466 15376 7472 15428
rect 7524 15416 7530 15428
rect 7668 15416 7696 15447
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 8220 15493 8248 15524
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 9490 15512 9496 15564
rect 9548 15552 9554 15564
rect 9861 15555 9919 15561
rect 9861 15552 9873 15555
rect 9548 15524 9873 15552
rect 9548 15512 9554 15524
rect 9861 15521 9873 15524
rect 9907 15521 9919 15555
rect 10226 15552 10232 15564
rect 9861 15515 9919 15521
rect 9968 15524 10232 15552
rect 8205 15487 8263 15493
rect 8205 15453 8217 15487
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15484 8355 15487
rect 8478 15484 8484 15496
rect 8343 15456 8484 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 8570 15444 8576 15496
rect 8628 15444 8634 15496
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9398 15484 9404 15496
rect 9171 15456 9404 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 8389 15419 8447 15425
rect 8389 15416 8401 15419
rect 7524 15388 7696 15416
rect 8266 15388 8401 15416
rect 7524 15376 7530 15388
rect 8266 15348 8294 15388
rect 8389 15385 8401 15388
rect 8435 15416 8447 15419
rect 9968 15416 9996 15524
rect 10226 15512 10232 15524
rect 10284 15512 10290 15564
rect 11238 15512 11244 15564
rect 11296 15512 11302 15564
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 12912 15561 12940 15592
rect 14826 15580 14832 15632
rect 14884 15620 14890 15632
rect 15102 15620 15108 15632
rect 14884 15592 15108 15620
rect 14884 15580 14890 15592
rect 15102 15580 15108 15592
rect 15160 15620 15166 15632
rect 15160 15592 15976 15620
rect 15160 15580 15166 15592
rect 11977 15555 12035 15561
rect 11977 15552 11989 15555
rect 11388 15524 11989 15552
rect 11388 15512 11394 15524
rect 11977 15521 11989 15524
rect 12023 15521 12035 15555
rect 11977 15515 12035 15521
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 14274 15552 14280 15564
rect 12943 15524 14280 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 14642 15512 14648 15564
rect 14700 15552 14706 15564
rect 14700 15524 15608 15552
rect 14700 15512 14706 15524
rect 10042 15444 10048 15496
rect 10100 15444 10106 15496
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 11256 15484 11284 15512
rect 12526 15484 12532 15496
rect 11256 15456 12532 15484
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 12618 15444 12624 15496
rect 12676 15444 12682 15496
rect 12802 15444 12808 15496
rect 12860 15444 12866 15496
rect 14752 15493 14780 15524
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14826 15444 14832 15496
rect 14884 15484 14890 15496
rect 14884 15456 14929 15484
rect 14884 15444 14890 15456
rect 15010 15444 15016 15496
rect 15068 15444 15074 15496
rect 15243 15487 15301 15493
rect 15243 15453 15255 15487
rect 15289 15484 15301 15487
rect 15470 15484 15476 15496
rect 15289 15456 15476 15484
rect 15289 15453 15301 15456
rect 15243 15447 15301 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 8435 15388 9996 15416
rect 10060 15416 10088 15444
rect 10870 15416 10876 15428
rect 10060 15388 10876 15416
rect 8435 15385 8447 15388
rect 8389 15379 8447 15385
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 10965 15419 11023 15425
rect 10965 15385 10977 15419
rect 11011 15416 11023 15419
rect 11425 15419 11483 15425
rect 11425 15416 11437 15419
rect 11011 15388 11437 15416
rect 11011 15385 11023 15388
rect 10965 15379 11023 15385
rect 11425 15385 11437 15388
rect 11471 15385 11483 15419
rect 15105 15419 15163 15425
rect 15105 15416 15117 15419
rect 11425 15379 11483 15385
rect 14936 15388 15117 15416
rect 14936 15360 14964 15388
rect 15105 15385 15117 15388
rect 15151 15385 15163 15419
rect 15105 15379 15163 15385
rect 6927 15320 8294 15348
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 10226 15308 10232 15360
rect 10284 15308 10290 15360
rect 10778 15308 10784 15360
rect 10836 15348 10842 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 10836 15320 11069 15348
rect 10836 15308 10842 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 12158 15308 12164 15360
rect 12216 15348 12222 15360
rect 13354 15348 13360 15360
rect 12216 15320 13360 15348
rect 12216 15308 12222 15320
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 14918 15308 14924 15360
rect 14976 15308 14982 15360
rect 15378 15308 15384 15360
rect 15436 15308 15442 15360
rect 15580 15348 15608 15524
rect 15838 15444 15844 15496
rect 15896 15444 15902 15496
rect 15948 15493 15976 15592
rect 15934 15487 15992 15493
rect 15934 15453 15946 15487
rect 15980 15453 15992 15487
rect 15934 15447 15992 15453
rect 16347 15487 16405 15493
rect 16347 15453 16359 15487
rect 16393 15484 16405 15487
rect 18340 15484 18368 15660
rect 19337 15657 19349 15660
rect 19383 15688 19395 15691
rect 19518 15688 19524 15700
rect 19383 15660 19524 15688
rect 19383 15657 19395 15660
rect 19337 15651 19395 15657
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 19794 15648 19800 15700
rect 19852 15688 19858 15700
rect 19889 15691 19947 15697
rect 19889 15688 19901 15691
rect 19852 15660 19901 15688
rect 19852 15648 19858 15660
rect 19889 15657 19901 15660
rect 19935 15657 19947 15691
rect 20257 15691 20315 15697
rect 20257 15688 20269 15691
rect 19889 15651 19947 15657
rect 19996 15660 20269 15688
rect 18601 15623 18659 15629
rect 18601 15589 18613 15623
rect 18647 15620 18659 15623
rect 18690 15620 18696 15632
rect 18647 15592 18696 15620
rect 18647 15589 18659 15592
rect 18601 15583 18659 15589
rect 18690 15580 18696 15592
rect 18748 15580 18754 15632
rect 18877 15623 18935 15629
rect 18877 15589 18889 15623
rect 18923 15620 18935 15623
rect 19996 15620 20024 15660
rect 20257 15657 20269 15660
rect 20303 15657 20315 15691
rect 20257 15651 20315 15657
rect 20625 15691 20683 15697
rect 20625 15657 20637 15691
rect 20671 15688 20683 15691
rect 20671 15660 21312 15688
rect 20671 15657 20683 15660
rect 20625 15651 20683 15657
rect 21177 15623 21235 15629
rect 21177 15620 21189 15623
rect 18923 15592 20024 15620
rect 20180 15592 21189 15620
rect 18923 15589 18935 15592
rect 18877 15583 18935 15589
rect 18414 15512 18420 15564
rect 18472 15552 18478 15564
rect 18472 15524 18920 15552
rect 18472 15512 18478 15524
rect 18892 15493 18920 15524
rect 16393 15456 18368 15484
rect 18877 15487 18935 15493
rect 16393 15453 16405 15456
rect 16347 15447 16405 15453
rect 18877 15453 18889 15487
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 19058 15444 19064 15496
rect 19116 15444 19122 15496
rect 19260 15493 19288 15592
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15552 19579 15555
rect 19610 15552 19616 15564
rect 19567 15524 19616 15552
rect 19567 15521 19579 15524
rect 19521 15515 19579 15521
rect 19610 15512 19616 15524
rect 19668 15552 19674 15564
rect 19797 15555 19855 15561
rect 19797 15552 19809 15555
rect 19668 15524 19809 15552
rect 19668 15512 19674 15524
rect 19797 15521 19809 15524
rect 19843 15521 19855 15555
rect 19797 15515 19855 15521
rect 19245 15487 19303 15493
rect 19245 15453 19257 15487
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 20180 15493 20208 15592
rect 21177 15589 21189 15592
rect 21223 15589 21235 15623
rect 21284 15620 21312 15660
rect 21358 15648 21364 15700
rect 21416 15648 21422 15700
rect 30558 15648 30564 15700
rect 30616 15688 30622 15700
rect 31113 15691 31171 15697
rect 31113 15688 31125 15691
rect 30616 15660 31125 15688
rect 30616 15648 30622 15660
rect 31113 15657 31125 15660
rect 31159 15688 31171 15691
rect 31202 15688 31208 15700
rect 31159 15660 31208 15688
rect 31159 15657 31171 15660
rect 31113 15651 31171 15657
rect 31202 15648 31208 15660
rect 31260 15648 31266 15700
rect 32766 15648 32772 15700
rect 32824 15688 32830 15700
rect 33137 15691 33195 15697
rect 33137 15688 33149 15691
rect 32824 15660 33149 15688
rect 32824 15648 32830 15660
rect 33137 15657 33149 15660
rect 33183 15657 33195 15691
rect 33137 15651 33195 15657
rect 33962 15648 33968 15700
rect 34020 15648 34026 15700
rect 34698 15648 34704 15700
rect 34756 15648 34762 15700
rect 34790 15648 34796 15700
rect 34848 15688 34854 15700
rect 34885 15691 34943 15697
rect 34885 15688 34897 15691
rect 34848 15660 34897 15688
rect 34848 15648 34854 15660
rect 34885 15657 34897 15660
rect 34931 15657 34943 15691
rect 34885 15651 34943 15657
rect 21910 15620 21916 15632
rect 21284 15592 21916 15620
rect 21177 15583 21235 15589
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 23106 15580 23112 15632
rect 23164 15580 23170 15632
rect 26234 15580 26240 15632
rect 26292 15620 26298 15632
rect 31849 15623 31907 15629
rect 26292 15592 31432 15620
rect 26292 15580 26298 15592
rect 21542 15512 21548 15564
rect 21600 15512 21606 15564
rect 23569 15555 23627 15561
rect 23569 15521 23581 15555
rect 23615 15552 23627 15555
rect 25130 15552 25136 15564
rect 23615 15524 25136 15552
rect 23615 15521 23627 15524
rect 23569 15515 23627 15521
rect 25130 15512 25136 15524
rect 25188 15512 25194 15564
rect 30466 15512 30472 15564
rect 30524 15552 30530 15564
rect 30524 15524 31340 15552
rect 30524 15512 30530 15524
rect 19981 15487 20039 15493
rect 19484 15456 19564 15484
rect 19484 15444 19490 15456
rect 15654 15376 15660 15428
rect 15712 15416 15718 15428
rect 16117 15419 16175 15425
rect 16117 15416 16129 15419
rect 15712 15388 16129 15416
rect 15712 15376 15718 15388
rect 16117 15385 16129 15388
rect 16163 15385 16175 15419
rect 16117 15379 16175 15385
rect 16209 15419 16267 15425
rect 16209 15385 16221 15419
rect 16255 15416 16267 15419
rect 16942 15416 16948 15428
rect 16255 15388 16948 15416
rect 16255 15385 16267 15388
rect 16209 15379 16267 15385
rect 16942 15376 16948 15388
rect 17000 15416 17006 15428
rect 17494 15416 17500 15428
rect 17000 15388 17500 15416
rect 17000 15376 17006 15388
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 19536 15425 19564 15456
rect 19981 15453 19993 15487
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20073 15487 20131 15493
rect 20073 15453 20085 15487
rect 20119 15484 20131 15487
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 20119 15456 20177 15484
rect 20119 15453 20131 15456
rect 20073 15447 20131 15453
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15484 20499 15487
rect 20622 15484 20628 15496
rect 20487 15456 20628 15484
rect 20487 15453 20499 15456
rect 20441 15447 20499 15453
rect 19521 15419 19579 15425
rect 19521 15385 19533 15419
rect 19567 15385 19579 15419
rect 19996 15416 20024 15447
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 20824 15456 21097 15484
rect 20346 15416 20352 15428
rect 19996 15388 20352 15416
rect 19521 15379 19579 15385
rect 20346 15376 20352 15388
rect 20404 15416 20410 15428
rect 20717 15419 20775 15425
rect 20717 15416 20729 15419
rect 20404 15388 20729 15416
rect 20404 15376 20410 15388
rect 20717 15385 20729 15388
rect 20763 15385 20775 15419
rect 20717 15379 20775 15385
rect 17310 15348 17316 15360
rect 15580 15320 17316 15348
rect 17310 15308 17316 15320
rect 17368 15308 17374 15360
rect 17862 15308 17868 15360
rect 17920 15348 17926 15360
rect 20824 15348 20852 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21560 15484 21588 15512
rect 21085 15447 21143 15453
rect 21192 15456 21588 15484
rect 20901 15419 20959 15425
rect 20901 15385 20913 15419
rect 20947 15416 20959 15419
rect 21192 15416 21220 15456
rect 23014 15444 23020 15496
rect 23072 15444 23078 15496
rect 23198 15444 23204 15496
rect 23256 15484 23262 15496
rect 30650 15493 30656 15496
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 23256 15456 23397 15484
rect 23256 15444 23262 15456
rect 23385 15453 23397 15456
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 30627 15487 30656 15493
rect 30627 15453 30639 15487
rect 30627 15447 30656 15453
rect 30650 15444 30656 15447
rect 30708 15444 30714 15496
rect 30742 15444 30748 15496
rect 30800 15444 30806 15496
rect 30929 15487 30987 15493
rect 30929 15453 30941 15487
rect 30975 15484 30987 15487
rect 31018 15484 31024 15496
rect 30975 15456 31024 15484
rect 30975 15453 30987 15456
rect 30929 15447 30987 15453
rect 31018 15444 31024 15456
rect 31076 15444 31082 15496
rect 31202 15444 31208 15496
rect 31260 15444 31266 15496
rect 31312 15493 31340 15524
rect 31298 15487 31356 15493
rect 31298 15453 31310 15487
rect 31344 15453 31356 15487
rect 31298 15447 31356 15453
rect 20947 15388 21220 15416
rect 20947 15385 20959 15388
rect 20901 15379 20959 15385
rect 21266 15376 21272 15428
rect 21324 15425 21330 15428
rect 21324 15419 21387 15425
rect 21324 15385 21341 15419
rect 21375 15385 21387 15419
rect 21324 15379 21387 15385
rect 21545 15419 21603 15425
rect 21545 15385 21557 15419
rect 21591 15416 21603 15419
rect 24946 15416 24952 15428
rect 21591 15388 24952 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 21324 15376 21330 15379
rect 17920 15320 20852 15348
rect 17920 15308 17926 15320
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 21560 15348 21588 15379
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 27338 15376 27344 15428
rect 27396 15416 27402 15428
rect 27396 15388 29960 15416
rect 27396 15376 27402 15388
rect 21232 15320 21588 15348
rect 21232 15308 21238 15320
rect 28074 15308 28080 15360
rect 28132 15348 28138 15360
rect 29822 15348 29828 15360
rect 28132 15320 29828 15348
rect 28132 15308 28138 15320
rect 29822 15308 29828 15320
rect 29880 15308 29886 15360
rect 29932 15348 29960 15388
rect 30374 15376 30380 15428
rect 30432 15416 30438 15428
rect 30837 15419 30895 15425
rect 30837 15416 30849 15419
rect 30432 15388 30849 15416
rect 30432 15376 30438 15388
rect 30760 15360 30788 15388
rect 30837 15385 30849 15388
rect 30883 15385 30895 15419
rect 30837 15379 30895 15385
rect 30558 15348 30564 15360
rect 29932 15320 30564 15348
rect 30558 15308 30564 15320
rect 30616 15308 30622 15360
rect 30742 15308 30748 15360
rect 30800 15308 30806 15360
rect 31312 15348 31340 15447
rect 31404 15416 31432 15592
rect 31849 15589 31861 15623
rect 31895 15620 31907 15623
rect 32858 15620 32864 15632
rect 31895 15592 32864 15620
rect 31895 15589 31907 15592
rect 31849 15583 31907 15589
rect 32858 15580 32864 15592
rect 32916 15580 32922 15632
rect 32950 15580 32956 15632
rect 33008 15620 33014 15632
rect 34238 15620 34244 15632
rect 33008 15592 33272 15620
rect 33008 15580 33014 15592
rect 31570 15552 31576 15564
rect 31496 15524 31576 15552
rect 31496 15493 31524 15524
rect 31570 15512 31576 15524
rect 31628 15512 31634 15564
rect 31754 15512 31760 15564
rect 31812 15552 31818 15564
rect 33045 15555 33103 15561
rect 33045 15552 33057 15555
rect 31812 15524 33057 15552
rect 31812 15512 31818 15524
rect 33045 15521 33057 15524
rect 33091 15521 33103 15555
rect 33045 15515 33103 15521
rect 33134 15512 33140 15564
rect 33192 15512 33198 15564
rect 33244 15561 33272 15592
rect 34164 15592 34244 15620
rect 34164 15561 34192 15592
rect 34238 15580 34244 15592
rect 34296 15580 34302 15632
rect 33229 15555 33287 15561
rect 33229 15521 33241 15555
rect 33275 15521 33287 15555
rect 33229 15515 33287 15521
rect 34149 15555 34207 15561
rect 34149 15521 34161 15555
rect 34195 15521 34207 15555
rect 34149 15515 34207 15521
rect 34606 15512 34612 15564
rect 34664 15552 34670 15564
rect 34977 15555 35035 15561
rect 34977 15552 34989 15555
rect 34664 15524 34989 15552
rect 34664 15512 34670 15524
rect 34977 15521 34989 15524
rect 35023 15521 35035 15555
rect 34977 15515 35035 15521
rect 31481 15487 31539 15493
rect 31481 15453 31493 15487
rect 31527 15453 31539 15487
rect 31481 15447 31539 15453
rect 31662 15444 31668 15496
rect 31720 15493 31726 15496
rect 31720 15484 31728 15493
rect 32769 15487 32827 15493
rect 31720 15456 31765 15484
rect 31720 15447 31728 15456
rect 32769 15453 32781 15487
rect 32815 15484 32827 15487
rect 32950 15484 32956 15496
rect 32815 15456 32956 15484
rect 32815 15453 32827 15456
rect 32769 15447 32827 15453
rect 31720 15444 31726 15447
rect 32950 15444 32956 15456
rect 33008 15444 33014 15496
rect 33152 15484 33180 15512
rect 33413 15487 33471 15493
rect 33413 15484 33425 15487
rect 33152 15456 33425 15484
rect 33413 15453 33425 15456
rect 33459 15453 33471 15487
rect 33413 15447 33471 15453
rect 34241 15487 34299 15493
rect 34241 15453 34253 15487
rect 34287 15484 34299 15487
rect 34514 15484 34520 15496
rect 34287 15456 34520 15484
rect 34287 15453 34299 15456
rect 34241 15447 34299 15453
rect 34514 15444 34520 15456
rect 34572 15444 34578 15496
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34624 15456 34897 15484
rect 31573 15419 31631 15425
rect 31573 15416 31585 15419
rect 31404 15388 31585 15416
rect 31573 15385 31585 15388
rect 31619 15385 31631 15419
rect 31573 15379 31631 15385
rect 33134 15376 33140 15428
rect 33192 15376 33198 15428
rect 33965 15419 34023 15425
rect 33965 15416 33977 15419
rect 33612 15388 33977 15416
rect 31754 15348 31760 15360
rect 31312 15320 31760 15348
rect 31754 15308 31760 15320
rect 31812 15308 31818 15360
rect 33612 15357 33640 15388
rect 33965 15385 33977 15388
rect 34011 15385 34023 15419
rect 33965 15379 34023 15385
rect 34624 15360 34652 15456
rect 34885 15453 34897 15456
rect 34931 15453 34943 15487
rect 34885 15447 34943 15453
rect 35161 15487 35219 15493
rect 35161 15453 35173 15487
rect 35207 15484 35219 15487
rect 35526 15484 35532 15496
rect 35207 15456 35532 15484
rect 35207 15453 35219 15456
rect 35161 15447 35219 15453
rect 35526 15444 35532 15456
rect 35584 15444 35590 15496
rect 33597 15351 33655 15357
rect 33597 15317 33609 15351
rect 33643 15317 33655 15351
rect 33597 15311 33655 15317
rect 34422 15308 34428 15360
rect 34480 15308 34486 15360
rect 34606 15308 34612 15360
rect 34664 15308 34670 15360
rect 1104 15258 36432 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 36432 15258
rect 1104 15184 36432 15206
rect 1964 15116 3832 15144
rect 1854 14968 1860 15020
rect 1912 15008 1918 15020
rect 1964 15017 1992 15116
rect 3234 15036 3240 15088
rect 3292 15036 3298 15088
rect 3804 15017 3832 15116
rect 5534 15104 5540 15156
rect 5592 15104 5598 15156
rect 9582 15144 9588 15156
rect 6196 15116 6868 15144
rect 4062 15036 4068 15088
rect 4120 15036 4126 15088
rect 4798 15036 4804 15088
rect 4856 15036 4862 15088
rect 1949 15011 2007 15017
rect 1949 15008 1961 15011
rect 1912 14980 1961 15008
rect 1912 14968 1918 14980
rect 1949 14977 1961 14980
rect 1995 14977 2007 15011
rect 1949 14971 2007 14977
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 14977 3847 15011
rect 3789 14971 3847 14977
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 5776 14980 5825 15008
rect 5776 14968 5782 14980
rect 5813 14977 5825 14980
rect 5859 14977 5871 15011
rect 6196 15008 6224 15116
rect 6270 15036 6276 15088
rect 6328 15076 6334 15088
rect 6328 15048 6684 15076
rect 6328 15036 6334 15048
rect 6656 15017 6684 15048
rect 6840 15020 6868 15116
rect 7852 15116 9588 15144
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 6196 14980 6377 15008
rect 5813 14971 5871 14977
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 2222 14900 2228 14952
rect 2280 14900 2286 14952
rect 3620 14912 5120 14940
rect 2038 14764 2044 14816
rect 2096 14804 2102 14816
rect 3620 14804 3648 14912
rect 3694 14832 3700 14884
rect 3752 14832 3758 14884
rect 5092 14872 5120 14912
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 5629 14943 5687 14949
rect 5629 14940 5641 14943
rect 5592 14912 5641 14940
rect 5592 14900 5598 14912
rect 5629 14909 5641 14912
rect 5675 14909 5687 14943
rect 5629 14903 5687 14909
rect 6564 14872 6592 14971
rect 6822 14968 6828 15020
rect 6880 14968 6886 15020
rect 7466 14968 7472 15020
rect 7524 14968 7530 15020
rect 7852 15017 7880 15116
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 10134 15104 10140 15156
rect 10192 15104 10198 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 15028 15116 15577 15144
rect 8110 15036 8116 15088
rect 8168 15036 8174 15088
rect 9766 15076 9772 15088
rect 9338 15048 9772 15076
rect 9766 15036 9772 15048
rect 9824 15036 9830 15088
rect 10152 15076 10180 15104
rect 10152 15048 10824 15076
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 14977 7711 15011
rect 7653 14971 7711 14977
rect 7837 15011 7895 15017
rect 7837 14977 7849 15011
rect 7883 14977 7895 15011
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 7837 14971 7895 14977
rect 9324 14980 9873 15008
rect 7668 14940 7696 14971
rect 9324 14952 9352 14980
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 15008 10195 15011
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 10183 14980 10333 15008
rect 10183 14977 10195 14980
rect 10137 14971 10195 14977
rect 10321 14977 10333 14980
rect 10367 14977 10379 15011
rect 10321 14971 10379 14977
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 9122 14940 9128 14952
rect 7668 14912 9128 14940
rect 9122 14900 9128 14912
rect 9180 14900 9186 14952
rect 9306 14900 9312 14952
rect 9364 14900 9370 14952
rect 9490 14900 9496 14952
rect 9548 14940 9554 14952
rect 9585 14943 9643 14949
rect 9585 14940 9597 14943
rect 9548 14912 9597 14940
rect 9548 14900 9554 14912
rect 9585 14909 9597 14912
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14940 10103 14943
rect 10226 14940 10232 14952
rect 10091 14912 10232 14940
rect 10091 14909 10103 14912
rect 10045 14903 10103 14909
rect 10226 14900 10232 14912
rect 10284 14900 10290 14952
rect 10520 14940 10548 14971
rect 10686 14968 10692 15020
rect 10744 14968 10750 15020
rect 10796 15017 10824 15048
rect 14918 15036 14924 15088
rect 14976 15076 14982 15088
rect 15028 15085 15056 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 17678 15104 17684 15156
rect 17736 15144 17742 15156
rect 17773 15147 17831 15153
rect 17773 15144 17785 15147
rect 17736 15116 17785 15144
rect 17736 15104 17742 15116
rect 17773 15113 17785 15116
rect 17819 15113 17831 15147
rect 18046 15144 18052 15156
rect 17773 15107 17831 15113
rect 17926 15116 18052 15144
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 14976 15048 15025 15076
rect 14976 15036 14982 15048
rect 15013 15045 15025 15048
rect 15059 15045 15071 15079
rect 17926 15076 17954 15116
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 19058 15104 19064 15156
rect 19116 15144 19122 15156
rect 19245 15147 19303 15153
rect 19245 15144 19257 15147
rect 19116 15116 19257 15144
rect 19116 15104 19122 15116
rect 19245 15113 19257 15116
rect 19291 15113 19303 15147
rect 19245 15107 19303 15113
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 21450 15144 21456 15156
rect 19576 15116 21456 15144
rect 19576 15104 19582 15116
rect 21450 15104 21456 15116
rect 21508 15104 21514 15156
rect 23014 15104 23020 15156
rect 23072 15144 23078 15156
rect 23753 15147 23811 15153
rect 23753 15144 23765 15147
rect 23072 15116 23765 15144
rect 23072 15104 23078 15116
rect 23753 15113 23765 15116
rect 23799 15113 23811 15147
rect 23753 15107 23811 15113
rect 24670 15104 24676 15156
rect 24728 15144 24734 15156
rect 24949 15147 25007 15153
rect 24949 15144 24961 15147
rect 24728 15116 24961 15144
rect 24728 15104 24734 15116
rect 24949 15113 24961 15116
rect 24995 15113 25007 15147
rect 24949 15107 25007 15113
rect 26970 15104 26976 15156
rect 27028 15144 27034 15156
rect 32122 15144 32128 15156
rect 27028 15116 32128 15144
rect 27028 15104 27034 15116
rect 32122 15104 32128 15116
rect 32180 15104 32186 15156
rect 32766 15104 32772 15156
rect 32824 15104 32830 15156
rect 15013 15039 15071 15045
rect 15304 15048 17954 15076
rect 20257 15079 20315 15085
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 15304 15017 15332 15048
rect 20257 15045 20269 15079
rect 20303 15076 20315 15079
rect 20346 15076 20352 15088
rect 20303 15048 20352 15076
rect 20303 15045 20315 15048
rect 20257 15039 20315 15045
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 20441 15079 20499 15085
rect 20441 15045 20453 15079
rect 20487 15076 20499 15079
rect 20806 15076 20812 15088
rect 20487 15048 20812 15076
rect 20487 15045 20499 15048
rect 20441 15039 20499 15045
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 23566 15036 23572 15088
rect 23624 15076 23630 15088
rect 24688 15076 24716 15104
rect 25498 15076 25504 15088
rect 23624 15048 24716 15076
rect 24780 15048 25504 15076
rect 23624 15036 23630 15048
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10928 14980 10977 15008
rect 10928 14968 10934 14980
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 10965 14971 11023 14977
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 10520 14912 10916 14940
rect 10888 14884 10916 14912
rect 15194 14900 15200 14952
rect 15252 14940 15258 14952
rect 15396 14940 15424 14971
rect 15470 14968 15476 15020
rect 15528 15008 15534 15020
rect 15654 15008 15660 15020
rect 15528 14980 15660 15008
rect 15528 14968 15534 14980
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 17402 14968 17408 15020
rect 17460 15008 17466 15020
rect 17926 15008 18276 15014
rect 18598 15008 18604 15020
rect 17460 14986 18604 15008
rect 17460 14980 17954 14986
rect 18248 14980 18604 14986
rect 17460 14968 17466 14980
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 19334 14968 19340 15020
rect 19392 14968 19398 15020
rect 20530 14968 20536 15020
rect 20588 14968 20594 15020
rect 23474 15008 23480 15020
rect 22066 14980 23480 15008
rect 16206 14940 16212 14952
rect 15252 14912 16212 14940
rect 15252 14900 15258 14912
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 17957 14943 18015 14949
rect 17957 14909 17969 14943
rect 18003 14909 18015 14943
rect 17957 14903 18015 14909
rect 5092 14844 6592 14872
rect 9398 14832 9404 14884
rect 9456 14872 9462 14884
rect 9953 14875 10011 14881
rect 9953 14872 9965 14875
rect 9456 14844 9965 14872
rect 9456 14832 9462 14844
rect 9953 14841 9965 14844
rect 9999 14841 10011 14875
rect 9953 14835 10011 14841
rect 10870 14832 10876 14884
rect 10928 14832 10934 14884
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 17972 14872 18000 14903
rect 18046 14900 18052 14952
rect 18104 14900 18110 14952
rect 18138 14900 18144 14952
rect 18196 14900 18202 14952
rect 18233 14943 18291 14949
rect 18233 14909 18245 14943
rect 18279 14940 18291 14943
rect 18322 14940 18328 14952
rect 18279 14912 18328 14940
rect 18279 14909 18291 14912
rect 18233 14903 18291 14909
rect 18322 14900 18328 14912
rect 18380 14940 18386 14952
rect 19242 14940 19248 14952
rect 18380 14912 19248 14940
rect 18380 14900 18386 14912
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 20990 14940 20996 14952
rect 19484 14912 20996 14940
rect 19484 14900 19490 14912
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 18966 14872 18972 14884
rect 12584 14844 15608 14872
rect 17972 14844 18972 14872
rect 12584 14832 12590 14844
rect 2096 14776 3648 14804
rect 5997 14807 6055 14813
rect 2096 14764 2102 14776
rect 5997 14773 6009 14807
rect 6043 14804 6055 14807
rect 6086 14804 6092 14816
rect 6043 14776 6092 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 6638 14764 6644 14816
rect 6696 14764 6702 14816
rect 7561 14807 7619 14813
rect 7561 14773 7573 14807
rect 7607 14804 7619 14807
rect 7650 14804 7656 14816
rect 7607 14776 7656 14804
rect 7607 14773 7619 14776
rect 7561 14767 7619 14773
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 11112 14776 11161 14804
rect 11112 14764 11118 14776
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 11149 14767 11207 14773
rect 15381 14807 15439 14813
rect 15381 14773 15393 14807
rect 15427 14804 15439 14807
rect 15470 14804 15476 14816
rect 15427 14776 15476 14804
rect 15427 14773 15439 14776
rect 15381 14767 15439 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15580 14804 15608 14844
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 20070 14832 20076 14884
rect 20128 14872 20134 14884
rect 20257 14875 20315 14881
rect 20257 14872 20269 14875
rect 20128 14844 20269 14872
rect 20128 14832 20134 14844
rect 20257 14841 20269 14844
rect 20303 14841 20315 14875
rect 20257 14835 20315 14841
rect 21358 14832 21364 14884
rect 21416 14872 21422 14884
rect 22066 14872 22094 14980
rect 23474 14968 23480 14980
rect 23532 15008 23538 15020
rect 23937 15011 23995 15017
rect 23937 15008 23949 15011
rect 23532 14980 23949 15008
rect 23532 14968 23538 14980
rect 23937 14977 23949 14980
rect 23983 15008 23995 15011
rect 24026 15008 24032 15020
rect 23983 14980 24032 15008
rect 23983 14977 23995 14980
rect 23937 14971 23995 14977
rect 24026 14968 24032 14980
rect 24084 15008 24090 15020
rect 24780 15008 24808 15048
rect 25498 15036 25504 15048
rect 25556 15036 25562 15088
rect 31846 15036 31852 15088
rect 31904 15076 31910 15088
rect 32401 15079 32459 15085
rect 32401 15076 32413 15079
rect 31904 15048 32413 15076
rect 31904 15036 31910 15048
rect 32401 15045 32413 15048
rect 32447 15045 32459 15079
rect 32401 15039 32459 15045
rect 32493 15079 32551 15085
rect 32493 15045 32505 15079
rect 32539 15076 32551 15079
rect 32674 15076 32680 15088
rect 32539 15048 32680 15076
rect 32539 15045 32551 15048
rect 32493 15039 32551 15045
rect 32674 15036 32680 15048
rect 32732 15036 32738 15088
rect 24084 14980 24808 15008
rect 25041 15011 25099 15017
rect 24084 14968 24090 14980
rect 25041 14977 25053 15011
rect 25087 15008 25099 15011
rect 26234 15008 26240 15020
rect 25087 14980 26240 15008
rect 25087 14977 25099 14980
rect 25041 14971 25099 14977
rect 26234 14968 26240 14980
rect 26292 14968 26298 15020
rect 27246 14968 27252 15020
rect 27304 15008 27310 15020
rect 27525 15011 27583 15017
rect 27525 15008 27537 15011
rect 27304 14980 27537 15008
rect 27304 14968 27310 14980
rect 27525 14977 27537 14980
rect 27571 14977 27583 15011
rect 27525 14971 27583 14977
rect 27706 14968 27712 15020
rect 27764 14968 27770 15020
rect 31754 14968 31760 15020
rect 31812 15008 31818 15020
rect 32306 15017 32312 15020
rect 32125 15011 32183 15017
rect 32125 15008 32137 15011
rect 31812 14980 32137 15008
rect 31812 14968 31818 14980
rect 32125 14977 32137 14980
rect 32171 14977 32183 15011
rect 32125 14971 32183 14977
rect 32283 15011 32312 15017
rect 32283 14977 32295 15011
rect 32283 14971 32312 14977
rect 32306 14968 32312 14971
rect 32364 14968 32370 15020
rect 32585 15011 32643 15017
rect 32585 14977 32597 15011
rect 32631 15008 32643 15011
rect 32950 15008 32956 15020
rect 32631 14980 32956 15008
rect 32631 14977 32643 14980
rect 32585 14971 32643 14977
rect 32950 14968 32956 14980
rect 33008 14968 33014 15020
rect 24210 14900 24216 14952
rect 24268 14900 24274 14952
rect 24765 14943 24823 14949
rect 24765 14909 24777 14943
rect 24811 14940 24823 14943
rect 25222 14940 25228 14952
rect 24811 14912 25228 14940
rect 24811 14909 24823 14912
rect 24765 14903 24823 14909
rect 25222 14900 25228 14912
rect 25280 14900 25286 14952
rect 25590 14900 25596 14952
rect 25648 14940 25654 14952
rect 25774 14940 25780 14952
rect 25648 14912 25780 14940
rect 25648 14900 25654 14912
rect 25774 14900 25780 14912
rect 25832 14940 25838 14952
rect 25832 14912 31754 14940
rect 25832 14900 25838 14912
rect 21416 14844 22094 14872
rect 21416 14832 21422 14844
rect 22738 14832 22744 14884
rect 22796 14872 22802 14884
rect 24121 14875 24179 14881
rect 22796 14844 23980 14872
rect 22796 14832 22802 14844
rect 21542 14804 21548 14816
rect 15580 14776 21548 14804
rect 21542 14764 21548 14776
rect 21600 14764 21606 14816
rect 23952 14804 23980 14844
rect 24121 14841 24133 14875
rect 24167 14872 24179 14875
rect 24167 14844 25268 14872
rect 24167 14841 24179 14844
rect 24121 14835 24179 14841
rect 24780 14816 24808 14844
rect 25240 14816 25268 14844
rect 30374 14832 30380 14884
rect 30432 14872 30438 14884
rect 31386 14872 31392 14884
rect 30432 14844 31392 14872
rect 30432 14832 30438 14844
rect 31386 14832 31392 14844
rect 31444 14832 31450 14884
rect 31726 14872 31754 14912
rect 33778 14872 33784 14884
rect 31726 14844 33784 14872
rect 33778 14832 33784 14844
rect 33836 14832 33842 14884
rect 24305 14807 24363 14813
rect 24305 14804 24317 14807
rect 23952 14776 24317 14804
rect 24305 14773 24317 14776
rect 24351 14773 24363 14807
rect 24305 14767 24363 14773
rect 24578 14764 24584 14816
rect 24636 14764 24642 14816
rect 24670 14764 24676 14816
rect 24728 14764 24734 14816
rect 24762 14764 24768 14816
rect 24820 14764 24826 14816
rect 25222 14764 25228 14816
rect 25280 14764 25286 14816
rect 27430 14764 27436 14816
rect 27488 14804 27494 14816
rect 27525 14807 27583 14813
rect 27525 14804 27537 14807
rect 27488 14776 27537 14804
rect 27488 14764 27494 14776
rect 27525 14773 27537 14776
rect 27571 14773 27583 14807
rect 27525 14767 27583 14773
rect 27893 14807 27951 14813
rect 27893 14773 27905 14807
rect 27939 14804 27951 14807
rect 34054 14804 34060 14816
rect 27939 14776 34060 14804
rect 27939 14773 27951 14776
rect 27893 14767 27951 14773
rect 34054 14764 34060 14776
rect 34112 14764 34118 14816
rect 1104 14714 36432 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 36432 14714
rect 1104 14640 36432 14662
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 2280 14572 3801 14600
rect 2280 14560 2286 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 3789 14563 3847 14569
rect 9217 14603 9275 14609
rect 9217 14569 9229 14603
rect 9263 14569 9275 14603
rect 9217 14563 9275 14569
rect 3605 14535 3663 14541
rect 3605 14501 3617 14535
rect 3651 14532 3663 14535
rect 4706 14532 4712 14544
rect 3651 14504 4712 14532
rect 3651 14501 3663 14504
rect 3605 14495 3663 14501
rect 4706 14492 4712 14504
rect 4764 14492 4770 14544
rect 7837 14535 7895 14541
rect 7837 14532 7849 14535
rect 6564 14504 7849 14532
rect 1854 14424 1860 14476
rect 1912 14424 1918 14476
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 4246 14464 4252 14476
rect 3844 14436 4252 14464
rect 3844 14424 3850 14436
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 5350 14464 5356 14476
rect 4488 14436 5356 14464
rect 4488 14424 4494 14436
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 6564 14473 6592 14504
rect 7837 14501 7849 14504
rect 7883 14532 7895 14535
rect 8478 14532 8484 14544
rect 7883 14504 8484 14532
rect 7883 14501 7895 14504
rect 7837 14495 7895 14501
rect 8478 14492 8484 14504
rect 8536 14492 8542 14544
rect 9232 14532 9260 14563
rect 9398 14560 9404 14612
rect 9456 14560 9462 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10502 14600 10508 14612
rect 9824 14572 10508 14600
rect 9824 14560 9830 14572
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 10686 14560 10692 14612
rect 10744 14600 10750 14612
rect 13262 14600 13268 14612
rect 10744 14572 13268 14600
rect 10744 14560 10750 14572
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 18414 14600 18420 14612
rect 14976 14572 18420 14600
rect 14976 14560 14982 14572
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 23014 14560 23020 14612
rect 23072 14600 23078 14612
rect 23293 14603 23351 14609
rect 23293 14600 23305 14603
rect 23072 14572 23305 14600
rect 23072 14560 23078 14572
rect 23293 14569 23305 14572
rect 23339 14569 23351 14603
rect 23293 14563 23351 14569
rect 24670 14560 24676 14612
rect 24728 14600 24734 14612
rect 25041 14603 25099 14609
rect 25041 14600 25053 14603
rect 24728 14572 25053 14600
rect 24728 14560 24734 14572
rect 25041 14569 25053 14572
rect 25087 14569 25099 14603
rect 25041 14563 25099 14569
rect 26142 14560 26148 14612
rect 26200 14600 26206 14612
rect 26237 14603 26295 14609
rect 26237 14600 26249 14603
rect 26200 14572 26249 14600
rect 26200 14560 26206 14572
rect 26237 14569 26249 14572
rect 26283 14569 26295 14603
rect 26237 14563 26295 14569
rect 27430 14560 27436 14612
rect 27488 14560 27494 14612
rect 30285 14603 30343 14609
rect 30285 14569 30297 14603
rect 30331 14600 30343 14603
rect 33781 14603 33839 14609
rect 33781 14600 33793 14603
rect 30331 14572 33793 14600
rect 30331 14569 30343 14572
rect 30285 14563 30343 14569
rect 33781 14569 33793 14572
rect 33827 14569 33839 14603
rect 33781 14563 33839 14569
rect 35250 14560 35256 14612
rect 35308 14600 35314 14612
rect 35434 14600 35440 14612
rect 35308 14572 35440 14600
rect 35308 14560 35314 14572
rect 35434 14560 35440 14572
rect 35492 14560 35498 14612
rect 10134 14532 10140 14544
rect 8588 14504 8800 14532
rect 9232 14504 10140 14532
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 7340 14436 7389 14464
rect 7340 14424 7346 14436
rect 7377 14433 7389 14436
rect 7423 14464 7435 14467
rect 8202 14464 8208 14476
rect 7423 14436 8208 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8588 14464 8616 14504
rect 8404 14436 8616 14464
rect 3234 14356 3240 14408
rect 3292 14356 3298 14408
rect 3694 14356 3700 14408
rect 3752 14396 3758 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 3752 14368 5181 14396
rect 3752 14356 3758 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14396 5779 14399
rect 5994 14396 6000 14408
rect 5767 14368 6000 14396
rect 5767 14365 5779 14368
rect 5721 14359 5779 14365
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 6822 14396 6828 14408
rect 6196 14368 6828 14396
rect 2133 14331 2191 14337
rect 2133 14297 2145 14331
rect 2179 14328 2191 14331
rect 2406 14328 2412 14340
rect 2179 14300 2412 14328
rect 2179 14297 2191 14300
rect 2133 14291 2191 14297
rect 2406 14288 2412 14300
rect 2464 14288 2470 14340
rect 4157 14331 4215 14337
rect 4157 14297 4169 14331
rect 4203 14328 4215 14331
rect 4617 14331 4675 14337
rect 4617 14328 4629 14331
rect 4203 14300 4629 14328
rect 4203 14297 4215 14300
rect 4157 14291 4215 14297
rect 4617 14297 4629 14300
rect 4663 14297 4675 14331
rect 4617 14291 4675 14297
rect 5537 14331 5595 14337
rect 5537 14297 5549 14331
rect 5583 14328 5595 14331
rect 6196 14328 6224 14368
rect 6822 14356 6828 14368
rect 6880 14396 6886 14408
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 6880 14368 7757 14396
rect 6880 14356 6886 14368
rect 7745 14365 7757 14368
rect 7791 14396 7803 14399
rect 8294 14396 8300 14408
rect 7791 14368 8300 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 8294 14356 8300 14368
rect 8352 14356 8358 14408
rect 8404 14405 8432 14436
rect 8662 14424 8668 14476
rect 8720 14424 8726 14476
rect 8772 14464 8800 14504
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 16206 14492 16212 14544
rect 16264 14532 16270 14544
rect 19426 14532 19432 14544
rect 16264 14504 19432 14532
rect 16264 14492 16270 14504
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 20714 14532 20720 14544
rect 19904 14504 20720 14532
rect 9766 14464 9772 14476
rect 8772 14436 9772 14464
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 9950 14424 9956 14476
rect 10008 14424 10014 14476
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 5583 14300 6224 14328
rect 6273 14331 6331 14337
rect 5583 14297 5595 14300
rect 5537 14291 5595 14297
rect 6273 14297 6285 14331
rect 6319 14328 6331 14331
rect 7193 14331 7251 14337
rect 6319 14300 6868 14328
rect 6319 14297 6331 14300
rect 6273 14291 6331 14297
rect 2498 14220 2504 14272
rect 2556 14260 2562 14272
rect 3694 14260 3700 14272
rect 2556 14232 3700 14260
rect 2556 14220 2562 14232
rect 3694 14220 3700 14232
rect 3752 14220 3758 14272
rect 5350 14220 5356 14272
rect 5408 14220 5414 14272
rect 5902 14220 5908 14272
rect 5960 14220 5966 14272
rect 6362 14220 6368 14272
rect 6420 14220 6426 14272
rect 6840 14269 6868 14300
rect 7193 14297 7205 14331
rect 7239 14328 7251 14331
rect 7466 14328 7472 14340
rect 7239 14300 7472 14328
rect 7239 14297 7251 14300
rect 7193 14291 7251 14297
rect 7466 14288 7472 14300
rect 7524 14328 7530 14340
rect 8404 14328 8432 14359
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 9306 14396 9312 14408
rect 8536 14368 9312 14396
rect 8536 14356 8542 14368
rect 9306 14356 9312 14368
rect 9364 14396 9370 14408
rect 10060 14396 10088 14427
rect 10502 14424 10508 14476
rect 10560 14464 10566 14476
rect 10781 14467 10839 14473
rect 10781 14464 10793 14467
rect 10560 14436 10793 14464
rect 10560 14424 10566 14436
rect 10781 14433 10793 14436
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 12342 14464 12348 14476
rect 11011 14436 12348 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 9364 14368 10088 14396
rect 10796 14396 10824 14427
rect 12342 14424 12348 14436
rect 12400 14464 12406 14476
rect 12894 14464 12900 14476
rect 12400 14436 12900 14464
rect 12400 14424 12406 14436
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 13228 14436 13400 14464
rect 13228 14424 13234 14436
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 10796 14368 11161 14396
rect 9364 14356 9370 14368
rect 11149 14365 11161 14368
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14396 11575 14399
rect 13081 14399 13139 14405
rect 13081 14396 13093 14399
rect 11563 14368 13093 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 13081 14365 13093 14368
rect 13127 14365 13139 14399
rect 13081 14359 13139 14365
rect 13262 14356 13268 14408
rect 13320 14356 13326 14408
rect 13372 14405 13400 14436
rect 18690 14424 18696 14476
rect 18748 14464 18754 14476
rect 19904 14464 19932 14504
rect 20714 14492 20720 14504
rect 20772 14492 20778 14544
rect 21634 14492 21640 14544
rect 21692 14532 21698 14544
rect 24486 14532 24492 14544
rect 21692 14504 24492 14532
rect 21692 14492 21698 14504
rect 24486 14492 24492 14504
rect 24544 14492 24550 14544
rect 25406 14492 25412 14544
rect 25464 14492 25470 14544
rect 25958 14492 25964 14544
rect 26016 14492 26022 14544
rect 27154 14492 27160 14544
rect 27212 14532 27218 14544
rect 34238 14532 34244 14544
rect 27212 14504 34244 14532
rect 27212 14492 27218 14504
rect 34238 14492 34244 14504
rect 34296 14492 34302 14544
rect 20533 14467 20591 14473
rect 20533 14464 20545 14467
rect 18748 14436 19932 14464
rect 19996 14436 20545 14464
rect 18748 14424 18754 14436
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13538 14356 13544 14408
rect 13596 14356 13602 14408
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14396 13691 14399
rect 13906 14396 13912 14408
rect 13679 14368 13912 14396
rect 13679 14365 13691 14368
rect 13633 14359 13691 14365
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 17678 14356 17684 14408
rect 17736 14396 17742 14408
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17736 14368 17785 14396
rect 17736 14356 17742 14368
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 17954 14356 17960 14408
rect 18012 14356 18018 14408
rect 19996 14405 20024 14436
rect 20533 14433 20545 14436
rect 20579 14433 20591 14467
rect 22554 14464 22560 14476
rect 20533 14427 20591 14433
rect 20824 14436 22560 14464
rect 20824 14408 20852 14436
rect 22554 14424 22560 14436
rect 22612 14424 22618 14476
rect 23198 14424 23204 14476
rect 23256 14464 23262 14476
rect 23477 14467 23535 14473
rect 23477 14464 23489 14467
rect 23256 14436 23489 14464
rect 23256 14424 23262 14436
rect 23477 14433 23489 14436
rect 23523 14433 23535 14467
rect 23477 14427 23535 14433
rect 25317 14467 25375 14473
rect 25317 14433 25329 14467
rect 25363 14464 25375 14467
rect 25363 14436 26096 14464
rect 25363 14433 25375 14436
rect 25317 14427 25375 14433
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 19889 14399 19947 14405
rect 18095 14368 19748 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 8846 14328 8852 14340
rect 7524 14300 8432 14328
rect 8496 14300 8852 14328
rect 7524 14288 7530 14300
rect 6825 14263 6883 14269
rect 6825 14229 6837 14263
rect 6871 14229 6883 14263
rect 6825 14223 6883 14229
rect 7282 14220 7288 14272
rect 7340 14220 7346 14272
rect 8021 14263 8079 14269
rect 8021 14229 8033 14263
rect 8067 14260 8079 14263
rect 8294 14260 8300 14272
rect 8067 14232 8300 14260
rect 8067 14229 8079 14232
rect 8021 14223 8079 14229
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 8496 14269 8524 14300
rect 8846 14288 8852 14300
rect 8904 14328 8910 14340
rect 9033 14331 9091 14337
rect 9033 14328 9045 14331
rect 8904 14300 9045 14328
rect 8904 14288 8910 14300
rect 9033 14297 9045 14300
rect 9079 14297 9091 14331
rect 9861 14331 9919 14337
rect 9033 14291 9091 14297
rect 9253 14300 9812 14328
rect 9253 14269 9281 14300
rect 8481 14263 8539 14269
rect 8481 14229 8493 14263
rect 8527 14229 8539 14263
rect 8481 14223 8539 14229
rect 9238 14263 9296 14269
rect 9238 14229 9250 14263
rect 9284 14229 9296 14263
rect 9238 14223 9296 14229
rect 9398 14220 9404 14272
rect 9456 14260 9462 14272
rect 9493 14263 9551 14269
rect 9493 14260 9505 14263
rect 9456 14232 9505 14260
rect 9456 14220 9462 14232
rect 9493 14229 9505 14232
rect 9539 14229 9551 14263
rect 9784 14260 9812 14300
rect 9861 14297 9873 14331
rect 9907 14328 9919 14331
rect 9907 14300 10364 14328
rect 9907 14297 9919 14300
rect 9861 14291 9919 14297
rect 10042 14260 10048 14272
rect 9784 14232 10048 14260
rect 9493 14223 9551 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 10336 14269 10364 14300
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 19245 14331 19303 14337
rect 19245 14328 19257 14331
rect 13780 14300 19257 14328
rect 13780 14288 13786 14300
rect 19245 14297 19257 14300
rect 19291 14297 19303 14331
rect 19245 14291 19303 14297
rect 10321 14263 10379 14269
rect 10321 14229 10333 14263
rect 10367 14229 10379 14263
rect 10321 14223 10379 14229
rect 10410 14220 10416 14272
rect 10468 14260 10474 14272
rect 10689 14263 10747 14269
rect 10689 14260 10701 14263
rect 10468 14232 10701 14260
rect 10468 14220 10474 14232
rect 10689 14229 10701 14232
rect 10735 14229 10747 14263
rect 10689 14223 10747 14229
rect 14734 14220 14740 14272
rect 14792 14260 14798 14272
rect 17589 14263 17647 14269
rect 17589 14260 17601 14263
rect 14792 14232 17601 14260
rect 14792 14220 14798 14232
rect 17589 14229 17601 14232
rect 17635 14229 17647 14263
rect 17589 14223 17647 14229
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18690 14260 18696 14272
rect 18104 14232 18696 14260
rect 18104 14220 18110 14232
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 19720 14260 19748 14368
rect 19889 14365 19901 14399
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 19904 14328 19932 14359
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 20128 14368 20269 14396
rect 20128 14356 20134 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20438 14356 20444 14408
rect 20496 14356 20502 14408
rect 20714 14356 20720 14408
rect 20772 14356 20778 14408
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 20990 14356 20996 14408
rect 21048 14356 21054 14408
rect 21082 14356 21088 14408
rect 21140 14356 21146 14408
rect 23382 14356 23388 14408
rect 23440 14356 23446 14408
rect 23566 14356 23572 14408
rect 23624 14356 23630 14408
rect 23750 14356 23756 14408
rect 23808 14356 23814 14408
rect 25225 14399 25283 14405
rect 25225 14365 25237 14399
rect 25271 14365 25283 14399
rect 25225 14359 25283 14365
rect 20898 14328 20904 14340
rect 19904 14300 20904 14328
rect 20898 14288 20904 14300
rect 20956 14328 20962 14340
rect 22646 14328 22652 14340
rect 20956 14300 22652 14328
rect 20956 14288 20962 14300
rect 22646 14288 22652 14300
rect 22704 14288 22710 14340
rect 22922 14288 22928 14340
rect 22980 14328 22986 14340
rect 23017 14331 23075 14337
rect 23017 14328 23029 14331
rect 22980 14300 23029 14328
rect 22980 14288 22986 14300
rect 23017 14297 23029 14300
rect 23063 14297 23075 14331
rect 25240 14328 25268 14359
rect 25498 14356 25504 14408
rect 25556 14396 25562 14408
rect 25777 14399 25835 14405
rect 25777 14396 25789 14399
rect 25556 14368 25789 14396
rect 25556 14356 25562 14368
rect 25777 14365 25789 14368
rect 25823 14365 25835 14399
rect 25777 14359 25835 14365
rect 25866 14356 25872 14408
rect 25924 14356 25930 14408
rect 26068 14405 26096 14436
rect 26878 14424 26884 14476
rect 26936 14464 26942 14476
rect 27801 14467 27859 14473
rect 27801 14464 27813 14467
rect 26936 14436 27813 14464
rect 26936 14424 26942 14436
rect 27801 14433 27813 14436
rect 27847 14464 27859 14467
rect 28169 14467 28227 14473
rect 28169 14464 28181 14467
rect 27847 14436 28181 14464
rect 27847 14433 27859 14436
rect 27801 14427 27859 14433
rect 28169 14433 28181 14436
rect 28215 14433 28227 14467
rect 30834 14464 30840 14476
rect 28169 14427 28227 14433
rect 29804 14436 30840 14464
rect 26053 14399 26111 14405
rect 26053 14365 26065 14399
rect 26099 14396 26111 14399
rect 26513 14399 26571 14405
rect 26513 14396 26525 14399
rect 26099 14368 26525 14396
rect 26099 14365 26111 14368
rect 26053 14359 26111 14365
rect 26513 14365 26525 14368
rect 26559 14365 26571 14399
rect 26513 14359 26571 14365
rect 26697 14399 26755 14405
rect 26697 14365 26709 14399
rect 26743 14365 26755 14399
rect 26697 14359 26755 14365
rect 25590 14328 25596 14340
rect 25240 14300 25596 14328
rect 23017 14291 23075 14297
rect 25590 14288 25596 14300
rect 25648 14288 25654 14340
rect 26712 14328 26740 14359
rect 26970 14356 26976 14408
rect 27028 14356 27034 14408
rect 27246 14356 27252 14408
rect 27304 14396 27310 14408
rect 27341 14399 27399 14405
rect 27341 14396 27353 14399
rect 27304 14368 27353 14396
rect 27304 14356 27310 14368
rect 27341 14365 27353 14368
rect 27387 14365 27399 14399
rect 27341 14359 27399 14365
rect 27617 14399 27675 14405
rect 27617 14365 27629 14399
rect 27663 14365 27675 14399
rect 27617 14359 27675 14365
rect 27062 14328 27068 14340
rect 26712 14300 27068 14328
rect 27062 14288 27068 14300
rect 27120 14328 27126 14340
rect 27522 14328 27528 14340
rect 27120 14300 27528 14328
rect 27120 14288 27126 14300
rect 27522 14288 27528 14300
rect 27580 14288 27586 14340
rect 26142 14260 26148 14272
rect 19720 14232 26148 14260
rect 26142 14220 26148 14232
rect 26200 14220 26206 14272
rect 26602 14220 26608 14272
rect 26660 14260 26666 14272
rect 26881 14263 26939 14269
rect 26881 14260 26893 14263
rect 26660 14232 26893 14260
rect 26660 14220 26666 14232
rect 26881 14229 26893 14232
rect 26927 14260 26939 14263
rect 27157 14263 27215 14269
rect 27157 14260 27169 14263
rect 26927 14232 27169 14260
rect 26927 14229 26939 14232
rect 26881 14223 26939 14229
rect 27157 14229 27169 14232
rect 27203 14229 27215 14263
rect 27632 14260 27660 14359
rect 27706 14356 27712 14408
rect 27764 14356 27770 14408
rect 27890 14356 27896 14408
rect 27948 14356 27954 14408
rect 29638 14356 29644 14408
rect 29696 14356 29702 14408
rect 29804 14405 29832 14436
rect 30834 14424 30840 14436
rect 30892 14424 30898 14476
rect 33502 14424 33508 14476
rect 33560 14464 33566 14476
rect 33873 14467 33931 14473
rect 33873 14464 33885 14467
rect 33560 14436 33885 14464
rect 33560 14424 33566 14436
rect 33873 14433 33885 14436
rect 33919 14433 33931 14467
rect 33873 14427 33931 14433
rect 29789 14399 29847 14405
rect 29789 14365 29801 14399
rect 29835 14365 29847 14399
rect 29789 14359 29847 14365
rect 30147 14399 30205 14405
rect 30147 14365 30159 14399
rect 30193 14396 30205 14399
rect 31662 14396 31668 14408
rect 30193 14368 31668 14396
rect 30193 14365 30205 14368
rect 30147 14359 30205 14365
rect 31662 14356 31668 14368
rect 31720 14356 31726 14408
rect 34054 14356 34060 14408
rect 34112 14356 34118 14408
rect 27724 14328 27752 14356
rect 28350 14328 28356 14340
rect 27724 14300 28356 14328
rect 28350 14288 28356 14300
rect 28408 14288 28414 14340
rect 28445 14331 28503 14337
rect 28445 14297 28457 14331
rect 28491 14328 28503 14331
rect 29086 14328 29092 14340
rect 28491 14300 29092 14328
rect 28491 14297 28503 14300
rect 28445 14291 28503 14297
rect 29086 14288 29092 14300
rect 29144 14288 29150 14340
rect 29917 14331 29975 14337
rect 29917 14297 29929 14331
rect 29963 14297 29975 14331
rect 29917 14291 29975 14297
rect 28810 14260 28816 14272
rect 27632 14232 28816 14260
rect 27157 14223 27215 14229
rect 28810 14220 28816 14232
rect 28868 14260 28874 14272
rect 29932 14260 29960 14291
rect 30006 14288 30012 14340
rect 30064 14288 30070 14340
rect 30374 14328 30380 14340
rect 30116 14300 30380 14328
rect 30116 14260 30144 14300
rect 30374 14288 30380 14300
rect 30432 14288 30438 14340
rect 30466 14288 30472 14340
rect 30524 14328 30530 14340
rect 30650 14328 30656 14340
rect 30524 14300 30656 14328
rect 30524 14288 30530 14300
rect 30650 14288 30656 14300
rect 30708 14328 30714 14340
rect 31202 14328 31208 14340
rect 30708 14300 31208 14328
rect 30708 14288 30714 14300
rect 31202 14288 31208 14300
rect 31260 14288 31266 14340
rect 31386 14288 31392 14340
rect 31444 14328 31450 14340
rect 32306 14328 32312 14340
rect 31444 14300 32312 14328
rect 31444 14288 31450 14300
rect 32306 14288 32312 14300
rect 32364 14288 32370 14340
rect 33502 14288 33508 14340
rect 33560 14328 33566 14340
rect 33686 14328 33692 14340
rect 33560 14300 33692 14328
rect 33560 14288 33566 14300
rect 33686 14288 33692 14300
rect 33744 14288 33750 14340
rect 33781 14331 33839 14337
rect 33781 14297 33793 14331
rect 33827 14328 33839 14331
rect 34606 14328 34612 14340
rect 33827 14300 34612 14328
rect 33827 14297 33839 14300
rect 33781 14291 33839 14297
rect 34606 14288 34612 14300
rect 34664 14288 34670 14340
rect 28868 14232 30144 14260
rect 28868 14220 28874 14232
rect 30190 14220 30196 14272
rect 30248 14260 30254 14272
rect 33318 14260 33324 14272
rect 30248 14232 33324 14260
rect 30248 14220 30254 14232
rect 33318 14220 33324 14232
rect 33376 14220 33382 14272
rect 34241 14263 34299 14269
rect 34241 14229 34253 14263
rect 34287 14260 34299 14263
rect 34514 14260 34520 14272
rect 34287 14232 34520 14260
rect 34287 14229 34299 14232
rect 34241 14223 34299 14229
rect 34514 14220 34520 14232
rect 34572 14260 34578 14272
rect 34974 14260 34980 14272
rect 34572 14232 34980 14260
rect 34572 14220 34578 14232
rect 34974 14220 34980 14232
rect 35032 14220 35038 14272
rect 1104 14170 36432 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 36432 14170
rect 1104 14096 36432 14118
rect 1854 14016 1860 14068
rect 1912 14016 1918 14068
rect 2406 14016 2412 14068
rect 2464 14056 2470 14068
rect 3237 14059 3295 14065
rect 3237 14056 3249 14059
rect 2464 14028 3249 14056
rect 2464 14016 2470 14028
rect 3237 14025 3249 14028
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 3694 14016 3700 14068
rect 3752 14016 3758 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5552 14028 5917 14056
rect 1872 13988 1900 14016
rect 5552 13988 5580 14028
rect 5905 14025 5917 14028
rect 5951 14056 5963 14059
rect 6362 14056 6368 14068
rect 5951 14028 6368 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6733 14059 6791 14065
rect 6733 14025 6745 14059
rect 6779 14056 6791 14059
rect 6822 14056 6828 14068
rect 6779 14028 6828 14056
rect 6779 14025 6791 14028
rect 6733 14019 6791 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 6917 14059 6975 14065
rect 6917 14025 6929 14059
rect 6963 14025 6975 14059
rect 6917 14019 6975 14025
rect 7377 14059 7435 14065
rect 7377 14025 7389 14059
rect 7423 14056 7435 14059
rect 7466 14056 7472 14068
rect 7423 14028 7472 14056
rect 7423 14025 7435 14028
rect 7377 14019 7435 14025
rect 6638 13988 6644 14000
rect 1412 13960 1900 13988
rect 3436 13960 5580 13988
rect 5828 13960 6644 13988
rect 1412 13929 1440 13960
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 3234 13920 3240 13932
rect 2832 13892 3240 13920
rect 2832 13880 2838 13892
rect 3234 13880 3240 13892
rect 3292 13880 3298 13932
rect 1670 13812 1676 13864
rect 1728 13812 1734 13864
rect 2038 13812 2044 13864
rect 2096 13852 2102 13864
rect 3436 13852 3464 13960
rect 5828 13932 5856 13960
rect 6638 13948 6644 13960
rect 6696 13948 6702 14000
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 4065 13923 4123 13929
rect 4065 13920 4077 13923
rect 3651 13892 4077 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 4065 13889 4077 13892
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 4246 13880 4252 13932
rect 4304 13920 4310 13932
rect 4304 13892 4660 13920
rect 4304 13880 4310 13892
rect 2096 13824 3464 13852
rect 3881 13855 3939 13861
rect 2096 13812 2102 13824
rect 3881 13821 3893 13855
rect 3927 13852 3939 13855
rect 4430 13852 4436 13864
rect 3927 13824 4436 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 4430 13812 4436 13824
rect 4488 13812 4494 13864
rect 4632 13852 4660 13892
rect 4706 13880 4712 13932
rect 4764 13880 4770 13932
rect 4801 13923 4859 13929
rect 4801 13889 4813 13923
rect 4847 13920 4859 13923
rect 4890 13920 4896 13932
rect 4847 13892 4896 13920
rect 4847 13889 4859 13892
rect 4801 13883 4859 13889
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13920 5227 13923
rect 5534 13920 5540 13932
rect 5215 13892 5540 13920
rect 5215 13889 5227 13892
rect 5169 13883 5227 13889
rect 5000 13852 5028 13883
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5626 13880 5632 13932
rect 5684 13880 5690 13932
rect 5810 13880 5816 13932
rect 5868 13880 5874 13932
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 6932 13920 6960 14019
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 7892 14028 7941 14056
rect 7892 14016 7898 14028
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 7929 14019 7987 14025
rect 8294 14016 8300 14068
rect 8352 14016 8358 14068
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 9030 14056 9036 14068
rect 8435 14028 9036 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 9030 14016 9036 14028
rect 9088 14016 9094 14068
rect 10778 14056 10784 14068
rect 9508 14028 10784 14056
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 9398 13988 9404 14000
rect 8260 13960 9404 13988
rect 8260 13948 8266 13960
rect 9398 13948 9404 13960
rect 9456 13948 9462 14000
rect 6871 13892 6960 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 7282 13880 7288 13932
rect 7340 13920 7346 13932
rect 8018 13920 8024 13932
rect 7340 13892 8024 13920
rect 7340 13880 7346 13892
rect 8018 13880 8024 13892
rect 8076 13920 8082 13932
rect 8076 13892 8616 13920
rect 8076 13880 8082 13892
rect 4632 13824 5028 13852
rect 5092 13824 5947 13852
rect 4816 13796 4844 13824
rect 2866 13744 2872 13796
rect 2924 13784 2930 13796
rect 3145 13787 3203 13793
rect 3145 13784 3157 13787
rect 2924 13756 3157 13784
rect 2924 13744 2930 13756
rect 3145 13753 3157 13756
rect 3191 13784 3203 13787
rect 3970 13784 3976 13796
rect 3191 13756 3976 13784
rect 3191 13753 3203 13756
rect 3145 13747 3203 13753
rect 3970 13744 3976 13756
rect 4028 13744 4034 13796
rect 4798 13744 4804 13796
rect 4856 13744 4862 13796
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 5092 13716 5120 13824
rect 5442 13744 5448 13796
rect 5500 13744 5506 13796
rect 5718 13744 5724 13796
rect 5776 13784 5782 13796
rect 5776 13756 5856 13784
rect 5776 13744 5782 13756
rect 5828 13725 5856 13756
rect 3108 13688 5120 13716
rect 5813 13719 5871 13725
rect 3108 13676 3114 13688
rect 5813 13685 5825 13719
rect 5859 13685 5871 13719
rect 5919 13716 5947 13824
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 6328 13824 6377 13852
rect 6328 13812 6334 13824
rect 6365 13821 6377 13824
rect 6411 13821 6423 13855
rect 6365 13815 6423 13821
rect 7469 13855 7527 13861
rect 7469 13821 7481 13855
rect 7515 13821 7527 13855
rect 7469 13815 7527 13821
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 7484 13784 7512 13815
rect 8478 13812 8484 13864
rect 8536 13812 8542 13864
rect 8588 13852 8616 13892
rect 8754 13880 8760 13932
rect 8812 13880 8818 13932
rect 8938 13880 8944 13932
rect 8996 13880 9002 13932
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 9508 13929 9536 14028
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11514 14056 11520 14068
rect 11379 14028 11520 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 13906 14016 13912 14068
rect 13964 14016 13970 14068
rect 15746 14016 15752 14068
rect 15804 14056 15810 14068
rect 15841 14059 15899 14065
rect 15841 14056 15853 14059
rect 15804 14028 15853 14056
rect 15804 14016 15810 14028
rect 15841 14025 15853 14028
rect 15887 14025 15899 14059
rect 15841 14019 15899 14025
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17678 14056 17684 14068
rect 17000 14028 17684 14056
rect 17000 14016 17006 14028
rect 17678 14016 17684 14028
rect 17736 14016 17742 14068
rect 21358 14016 21364 14068
rect 21416 14016 21422 14068
rect 21542 14016 21548 14068
rect 21600 14056 21606 14068
rect 25593 14059 25651 14065
rect 21600 14028 22140 14056
rect 21600 14016 21606 14028
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 9180 13892 9229 13920
rect 9180 13880 9186 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 9582 13880 9588 13932
rect 9640 13880 9646 13932
rect 10962 13880 10968 13932
rect 11020 13880 11026 13932
rect 11532 13920 11560 14016
rect 12253 13991 12311 13997
rect 12253 13957 12265 13991
rect 12299 13988 12311 13991
rect 12894 13988 12900 14000
rect 12299 13960 12900 13988
rect 12299 13957 12311 13960
rect 12253 13951 12311 13957
rect 12894 13948 12900 13960
rect 12952 13948 12958 14000
rect 14369 13991 14427 13997
rect 14369 13957 14381 13991
rect 14415 13988 14427 13991
rect 16669 13991 16727 13997
rect 16669 13988 16681 13991
rect 14415 13960 16681 13988
rect 14415 13957 14427 13960
rect 14369 13951 14427 13957
rect 16669 13957 16681 13960
rect 16715 13957 16727 13991
rect 17862 13988 17868 14000
rect 16669 13951 16727 13957
rect 16868 13960 17868 13988
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11532 13892 12081 13920
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12710 13920 12716 13932
rect 12483 13892 12716 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 12710 13880 12716 13892
rect 12768 13920 12774 13932
rect 13998 13920 14004 13932
rect 12768 13892 14004 13920
rect 12768 13880 12774 13892
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13920 14151 13923
rect 14734 13920 14740 13932
rect 14139 13892 14740 13920
rect 14139 13889 14151 13892
rect 14093 13883 14151 13889
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16071 13892 16252 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 8846 13852 8852 13864
rect 8588 13824 8852 13852
rect 8846 13812 8852 13824
rect 8904 13852 8910 13864
rect 8904 13824 8984 13852
rect 8904 13812 8910 13824
rect 6788 13756 7512 13784
rect 8956 13784 8984 13824
rect 9030 13812 9036 13864
rect 9088 13852 9094 13864
rect 9600 13852 9628 13880
rect 9088 13824 9628 13852
rect 9088 13812 9094 13824
rect 9858 13812 9864 13864
rect 9916 13812 9922 13864
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13852 12679 13855
rect 13078 13852 13084 13864
rect 12667 13824 13084 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 13078 13812 13084 13824
rect 13136 13852 13142 13864
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 13136 13824 14197 13852
rect 13136 13812 13142 13824
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 14185 13815 14243 13821
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15068 13824 16129 13852
rect 15068 13812 15074 13824
rect 16117 13821 16129 13824
rect 16163 13821 16175 13855
rect 16224 13852 16252 13892
rect 16298 13880 16304 13932
rect 16356 13880 16362 13932
rect 16868 13929 16896 13960
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 21818 13988 21824 14000
rect 21192 13960 21824 13988
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 16942 13880 16948 13932
rect 17000 13880 17006 13932
rect 17126 13880 17132 13932
rect 17184 13880 17190 13932
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13920 17279 13923
rect 17310 13920 17316 13932
rect 17267 13892 17316 13920
rect 17267 13889 17279 13892
rect 17221 13883 17279 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 21192 13929 21220 13960
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 22112 13997 22140 14028
rect 25593 14025 25605 14059
rect 25639 14056 25651 14059
rect 25866 14056 25872 14068
rect 25639 14028 25872 14056
rect 25639 14025 25651 14028
rect 25593 14019 25651 14025
rect 25866 14016 25872 14028
rect 25924 14016 25930 14068
rect 26142 14016 26148 14068
rect 26200 14016 26206 14068
rect 27617 14059 27675 14065
rect 27617 14025 27629 14059
rect 27663 14056 27675 14059
rect 27890 14056 27896 14068
rect 27663 14028 27896 14056
rect 27663 14025 27675 14028
rect 27617 14019 27675 14025
rect 27890 14016 27896 14028
rect 27948 14016 27954 14068
rect 28353 14059 28411 14065
rect 28353 14025 28365 14059
rect 28399 14056 28411 14059
rect 30650 14056 30656 14068
rect 28399 14028 30656 14056
rect 28399 14025 28411 14028
rect 28353 14019 28411 14025
rect 30650 14016 30656 14028
rect 30708 14016 30714 14068
rect 30834 14016 30840 14068
rect 30892 14056 30898 14068
rect 31665 14059 31723 14065
rect 30892 14028 31157 14056
rect 30892 14016 30898 14028
rect 22097 13991 22155 13997
rect 22097 13957 22109 13991
rect 22143 13957 22155 13991
rect 25133 13991 25191 13997
rect 25133 13988 25145 13991
rect 22097 13951 22155 13957
rect 22480 13960 22876 13988
rect 21177 13923 21235 13929
rect 19208 13892 21128 13920
rect 19208 13880 19214 13892
rect 17144 13852 17172 13880
rect 16224 13824 17172 13852
rect 16117 13815 16175 13821
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 17644 13824 18460 13852
rect 17644 13812 17650 13824
rect 8956 13756 9720 13784
rect 6788 13744 6794 13756
rect 8662 13716 8668 13728
rect 5919 13688 8668 13716
rect 5813 13679 5871 13685
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 8846 13676 8852 13728
rect 8904 13676 8910 13728
rect 9401 13719 9459 13725
rect 9401 13685 9413 13719
rect 9447 13716 9459 13719
rect 9490 13716 9496 13728
rect 9447 13688 9496 13716
rect 9447 13685 9459 13688
rect 9401 13679 9459 13685
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 9692 13716 9720 13756
rect 12434 13744 12440 13796
rect 12492 13784 12498 13796
rect 12710 13784 12716 13796
rect 12492 13756 12716 13784
rect 12492 13744 12498 13756
rect 12710 13744 12716 13756
rect 12768 13784 12774 13796
rect 18432 13784 18460 13824
rect 19794 13812 19800 13864
rect 19852 13852 19858 13864
rect 20530 13852 20536 13864
rect 19852 13824 20536 13852
rect 19852 13812 19858 13824
rect 20530 13812 20536 13824
rect 20588 13852 20594 13864
rect 20993 13855 21051 13861
rect 20993 13852 21005 13855
rect 20588 13824 21005 13852
rect 20588 13812 20594 13824
rect 20993 13821 21005 13824
rect 21039 13821 21051 13855
rect 21100 13852 21128 13892
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 21453 13923 21511 13929
rect 21453 13889 21465 13923
rect 21499 13920 21511 13923
rect 21634 13920 21640 13932
rect 21499 13892 21640 13920
rect 21499 13889 21511 13892
rect 21453 13883 21511 13889
rect 21634 13880 21640 13892
rect 21692 13880 21698 13932
rect 21836 13920 21864 13948
rect 22480 13920 22508 13960
rect 21836 13892 22508 13920
rect 22554 13880 22560 13932
rect 22612 13880 22618 13932
rect 22646 13880 22652 13932
rect 22704 13920 22710 13932
rect 22848 13929 22876 13960
rect 24412 13960 25145 13988
rect 22741 13923 22799 13929
rect 22741 13920 22753 13923
rect 22704 13892 22753 13920
rect 22704 13880 22710 13892
rect 22741 13889 22753 13892
rect 22787 13889 22799 13923
rect 22741 13883 22799 13889
rect 22833 13923 22891 13929
rect 22833 13889 22845 13923
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 23017 13923 23075 13929
rect 23017 13889 23029 13923
rect 23063 13920 23075 13923
rect 23198 13920 23204 13932
rect 23063 13892 23204 13920
rect 23063 13889 23075 13892
rect 23017 13883 23075 13889
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 24210 13880 24216 13932
rect 24268 13880 24274 13932
rect 24412 13929 24440 13960
rect 25133 13957 25145 13960
rect 25179 13988 25191 13991
rect 26329 13991 26387 13997
rect 25179 13960 26280 13988
rect 25179 13957 25191 13960
rect 25133 13951 25191 13957
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 24486 13880 24492 13932
rect 24544 13880 24550 13932
rect 24946 13880 24952 13932
rect 25004 13920 25010 13932
rect 25409 13923 25467 13929
rect 25409 13920 25421 13923
rect 25004 13892 25421 13920
rect 25004 13880 25010 13892
rect 25409 13889 25421 13892
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 21100 13824 25237 13852
rect 20993 13815 21051 13821
rect 25225 13821 25237 13824
rect 25271 13852 25283 13855
rect 25314 13852 25320 13864
rect 25271 13824 25320 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 25314 13812 25320 13824
rect 25372 13812 25378 13864
rect 26252 13852 26280 13960
rect 26329 13957 26341 13991
rect 26375 13988 26387 13991
rect 27154 13988 27160 14000
rect 26375 13960 27160 13988
rect 26375 13957 26387 13960
rect 26329 13951 26387 13957
rect 27154 13948 27160 13960
rect 27212 13948 27218 14000
rect 27249 13991 27307 13997
rect 27249 13957 27261 13991
rect 27295 13957 27307 13991
rect 27249 13951 27307 13957
rect 27465 13991 27523 13997
rect 27465 13957 27477 13991
rect 27511 13988 27523 13991
rect 27798 13988 27804 14000
rect 27511 13960 27804 13988
rect 27511 13957 27523 13960
rect 27465 13951 27523 13957
rect 26513 13923 26571 13929
rect 26513 13889 26525 13923
rect 26559 13920 26571 13923
rect 26694 13920 26700 13932
rect 26559 13892 26700 13920
rect 26559 13889 26571 13892
rect 26513 13883 26571 13889
rect 26694 13880 26700 13892
rect 26752 13880 26758 13932
rect 27264 13920 27292 13951
rect 27798 13948 27804 13960
rect 27856 13948 27862 14000
rect 28721 13991 28779 13997
rect 28721 13957 28733 13991
rect 28767 13988 28779 13991
rect 29086 13988 29092 14000
rect 28767 13960 29092 13988
rect 28767 13957 28779 13960
rect 28721 13951 28779 13957
rect 29086 13948 29092 13960
rect 29144 13988 29150 14000
rect 29822 13988 29828 14000
rect 29144 13960 29828 13988
rect 29144 13948 29150 13960
rect 29822 13948 29828 13960
rect 29880 13948 29886 14000
rect 28537 13923 28595 13929
rect 27264 13892 27568 13920
rect 27540 13864 27568 13892
rect 28537 13889 28549 13923
rect 28583 13889 28595 13923
rect 28537 13883 28595 13889
rect 28629 13923 28687 13929
rect 28629 13889 28641 13923
rect 28675 13920 28687 13923
rect 28810 13920 28816 13932
rect 28675 13892 28816 13920
rect 28675 13889 28687 13892
rect 28629 13883 28687 13889
rect 26326 13852 26332 13864
rect 26252 13824 26332 13852
rect 26326 13812 26332 13824
rect 26384 13812 26390 13864
rect 27522 13812 27528 13864
rect 27580 13812 27586 13864
rect 28552 13852 28580 13883
rect 28810 13880 28816 13892
rect 28868 13880 28874 13932
rect 28902 13880 28908 13932
rect 28960 13880 28966 13932
rect 28994 13880 29000 13932
rect 29052 13880 29058 13932
rect 30926 13880 30932 13932
rect 30984 13920 30990 13932
rect 31129 13929 31157 14028
rect 31665 14025 31677 14059
rect 31711 14056 31723 14059
rect 32490 14056 32496 14068
rect 31711 14028 32496 14056
rect 31711 14025 31723 14028
rect 31665 14019 31723 14025
rect 32490 14016 32496 14028
rect 32548 14016 32554 14068
rect 32861 14059 32919 14065
rect 32861 14025 32873 14059
rect 32907 14056 32919 14059
rect 33226 14056 33232 14068
rect 32907 14028 33232 14056
rect 32907 14025 32919 14028
rect 32861 14019 32919 14025
rect 33226 14016 33232 14028
rect 33284 14016 33290 14068
rect 33597 14059 33655 14065
rect 33597 14025 33609 14059
rect 33643 14056 33655 14059
rect 33778 14056 33784 14068
rect 33643 14028 33784 14056
rect 33643 14025 33655 14028
rect 33597 14019 33655 14025
rect 33778 14016 33784 14028
rect 33836 14016 33842 14068
rect 34330 14016 34336 14068
rect 34388 14056 34394 14068
rect 34514 14056 34520 14068
rect 34388 14028 34520 14056
rect 34388 14016 34394 14028
rect 34514 14016 34520 14028
rect 34572 14016 34578 14068
rect 35345 14059 35403 14065
rect 35345 14025 35357 14059
rect 35391 14025 35403 14059
rect 35345 14019 35403 14025
rect 31202 13948 31208 14000
rect 31260 13988 31266 14000
rect 31297 13991 31355 13997
rect 31297 13988 31309 13991
rect 31260 13960 31309 13988
rect 31260 13948 31266 13960
rect 31297 13957 31309 13960
rect 31343 13957 31355 13991
rect 31297 13951 31355 13957
rect 33318 13948 33324 14000
rect 33376 13988 33382 14000
rect 34885 13991 34943 13997
rect 34885 13988 34897 13991
rect 33376 13960 34897 13988
rect 33376 13948 33382 13960
rect 34885 13957 34897 13960
rect 34931 13957 34943 13991
rect 34885 13951 34943 13957
rect 31021 13923 31079 13929
rect 31021 13920 31033 13923
rect 30984 13892 31033 13920
rect 30984 13880 30990 13892
rect 31021 13889 31033 13892
rect 31067 13889 31079 13923
rect 31021 13883 31079 13889
rect 31114 13923 31172 13929
rect 31114 13889 31126 13923
rect 31160 13889 31172 13923
rect 31114 13883 31172 13889
rect 31389 13923 31447 13929
rect 31389 13889 31401 13923
rect 31435 13889 31447 13923
rect 31389 13883 31447 13889
rect 31527 13923 31585 13929
rect 31527 13889 31539 13923
rect 31573 13920 31585 13923
rect 31573 13889 31600 13920
rect 31527 13883 31600 13889
rect 29914 13852 29920 13864
rect 28552 13824 29920 13852
rect 29914 13812 29920 13824
rect 29972 13812 29978 13864
rect 31404 13852 31432 13883
rect 30944 13824 31432 13852
rect 31572 13852 31600 13883
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 32401 13923 32459 13929
rect 32401 13920 32413 13923
rect 31720 13892 32413 13920
rect 31720 13880 31726 13892
rect 32401 13889 32413 13892
rect 32447 13889 32459 13923
rect 32401 13883 32459 13889
rect 32677 13923 32735 13929
rect 32677 13889 32689 13923
rect 32723 13920 32735 13923
rect 32766 13920 32772 13932
rect 32723 13892 32772 13920
rect 32723 13889 32735 13892
rect 32677 13883 32735 13889
rect 32766 13880 32772 13892
rect 32824 13880 32830 13932
rect 33781 13923 33839 13929
rect 33781 13889 33793 13923
rect 33827 13920 33839 13923
rect 33962 13920 33968 13932
rect 33827 13892 33968 13920
rect 33827 13889 33839 13892
rect 33781 13883 33839 13889
rect 33962 13880 33968 13892
rect 34020 13880 34026 13932
rect 34057 13923 34115 13929
rect 34057 13889 34069 13923
rect 34103 13920 34115 13923
rect 34146 13920 34152 13932
rect 34103 13892 34152 13920
rect 34103 13889 34115 13892
rect 34057 13883 34115 13889
rect 34146 13880 34152 13892
rect 34204 13880 34210 13932
rect 35066 13880 35072 13932
rect 35124 13880 35130 13932
rect 35161 13923 35219 13929
rect 35161 13889 35173 13923
rect 35207 13889 35219 13923
rect 35360 13920 35388 14019
rect 35434 14016 35440 14068
rect 35492 14056 35498 14068
rect 35805 14059 35863 14065
rect 35805 14056 35817 14059
rect 35492 14028 35817 14056
rect 35492 14016 35498 14028
rect 35805 14025 35817 14028
rect 35851 14025 35863 14059
rect 35805 14019 35863 14025
rect 35437 13923 35495 13929
rect 35437 13920 35449 13923
rect 35360 13892 35449 13920
rect 35161 13883 35219 13889
rect 35437 13889 35449 13892
rect 35483 13889 35495 13923
rect 35437 13883 35495 13889
rect 31754 13852 31760 13864
rect 31572 13824 31760 13852
rect 30944 13796 30972 13824
rect 31754 13812 31760 13824
rect 31812 13812 31818 13864
rect 32490 13812 32496 13864
rect 32548 13812 32554 13864
rect 33226 13812 33232 13864
rect 33284 13852 33290 13864
rect 33873 13855 33931 13861
rect 33873 13852 33885 13855
rect 33284 13824 33885 13852
rect 33284 13812 33290 13824
rect 33873 13821 33885 13824
rect 33919 13821 33931 13855
rect 33873 13815 33931 13821
rect 19886 13784 19892 13796
rect 12768 13756 18368 13784
rect 18432 13756 19892 13784
rect 12768 13744 12774 13756
rect 18340 13728 18368 13756
rect 19886 13744 19892 13756
rect 19944 13784 19950 13796
rect 21358 13784 21364 13796
rect 19944 13756 21364 13784
rect 19944 13744 19950 13756
rect 21358 13744 21364 13756
rect 21416 13744 21422 13796
rect 22370 13744 22376 13796
rect 22428 13784 22434 13796
rect 22922 13784 22928 13796
rect 22428 13756 22928 13784
rect 22428 13744 22434 13756
rect 22922 13744 22928 13756
rect 22980 13744 22986 13796
rect 23382 13744 23388 13796
rect 23440 13784 23446 13796
rect 24029 13787 24087 13793
rect 24029 13784 24041 13787
rect 23440 13756 24041 13784
rect 23440 13744 23446 13756
rect 24029 13753 24041 13756
rect 24075 13753 24087 13787
rect 24029 13747 24087 13753
rect 25682 13744 25688 13796
rect 25740 13784 25746 13796
rect 29454 13784 29460 13796
rect 25740 13756 29460 13784
rect 25740 13744 25746 13756
rect 29454 13744 29460 13756
rect 29512 13744 29518 13796
rect 30926 13744 30932 13796
rect 30984 13744 30990 13796
rect 33244 13784 33272 13812
rect 35176 13784 35204 13883
rect 35250 13812 35256 13864
rect 35308 13852 35314 13864
rect 35529 13855 35587 13861
rect 35529 13852 35541 13855
rect 35308 13824 35541 13852
rect 35308 13812 35314 13824
rect 35529 13821 35541 13824
rect 35575 13821 35587 13855
rect 35529 13815 35587 13821
rect 32692 13756 33272 13784
rect 33796 13756 35204 13784
rect 10410 13716 10416 13728
rect 9692 13688 10416 13716
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 11514 13676 11520 13728
rect 11572 13676 11578 13728
rect 14369 13719 14427 13725
rect 14369 13685 14381 13719
rect 14415 13716 14427 13719
rect 15010 13716 15016 13728
rect 14415 13688 15016 13716
rect 14415 13685 14427 13688
rect 14369 13679 14427 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 16301 13719 16359 13725
rect 16301 13716 16313 13719
rect 15344 13688 16313 13716
rect 15344 13676 15350 13688
rect 16301 13685 16313 13688
rect 16347 13716 16359 13719
rect 18230 13716 18236 13728
rect 16347 13688 18236 13716
rect 16347 13685 16359 13688
rect 16301 13679 16359 13685
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 18322 13676 18328 13728
rect 18380 13716 18386 13728
rect 22462 13716 22468 13728
rect 18380 13688 22468 13716
rect 18380 13676 18386 13688
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 25406 13676 25412 13728
rect 25464 13676 25470 13728
rect 26418 13676 26424 13728
rect 26476 13716 26482 13728
rect 27433 13719 27491 13725
rect 27433 13716 27445 13719
rect 26476 13688 27445 13716
rect 26476 13676 26482 13688
rect 27433 13685 27445 13688
rect 27479 13685 27491 13719
rect 27433 13679 27491 13685
rect 31110 13676 31116 13728
rect 31168 13716 31174 13728
rect 31478 13716 31484 13728
rect 31168 13688 31484 13716
rect 31168 13676 31174 13688
rect 31478 13676 31484 13688
rect 31536 13676 31542 13728
rect 32692 13725 32720 13756
rect 32677 13719 32735 13725
rect 32677 13685 32689 13719
rect 32723 13685 32735 13719
rect 32677 13679 32735 13685
rect 33686 13676 33692 13728
rect 33744 13716 33750 13728
rect 33796 13725 33824 13756
rect 33781 13719 33839 13725
rect 33781 13716 33793 13719
rect 33744 13688 33793 13716
rect 33744 13676 33750 13688
rect 33781 13685 33793 13688
rect 33827 13685 33839 13719
rect 33781 13679 33839 13685
rect 34790 13676 34796 13728
rect 34848 13716 34854 13728
rect 34885 13719 34943 13725
rect 34885 13716 34897 13719
rect 34848 13688 34897 13716
rect 34848 13676 34854 13688
rect 34885 13685 34897 13688
rect 34931 13685 34943 13719
rect 34885 13679 34943 13685
rect 34974 13676 34980 13728
rect 35032 13716 35038 13728
rect 35437 13719 35495 13725
rect 35437 13716 35449 13719
rect 35032 13688 35449 13716
rect 35032 13676 35038 13688
rect 35437 13685 35449 13688
rect 35483 13685 35495 13719
rect 35437 13679 35495 13685
rect 1104 13626 36432 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 36432 13626
rect 1104 13552 36432 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 1728 13484 2421 13512
rect 1728 13472 1734 13484
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 2409 13475 2467 13481
rect 4430 13472 4436 13524
rect 4488 13472 4494 13524
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 4985 13515 5043 13521
rect 4985 13512 4997 13515
rect 4764 13484 4997 13512
rect 4764 13472 4770 13484
rect 4985 13481 4997 13484
rect 5031 13512 5043 13515
rect 5350 13512 5356 13524
rect 5031 13484 5356 13512
rect 5031 13481 5043 13484
rect 4985 13475 5043 13481
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 5537 13515 5595 13521
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 5810 13512 5816 13524
rect 5583 13484 5816 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 9766 13512 9772 13524
rect 6788 13484 9772 13512
rect 6788 13472 6794 13484
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 9953 13515 10011 13521
rect 9953 13512 9965 13515
rect 9916 13484 9965 13512
rect 9916 13472 9922 13484
rect 9953 13481 9965 13484
rect 9999 13481 10011 13515
rect 9953 13475 10011 13481
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 12584 13484 12725 13512
rect 12584 13472 12590 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 12713 13475 12771 13481
rect 14734 13472 14740 13524
rect 14792 13472 14798 13524
rect 16577 13515 16635 13521
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 17126 13512 17132 13524
rect 16623 13484 17132 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 4801 13447 4859 13453
rect 4801 13413 4813 13447
rect 4847 13444 4859 13447
rect 5258 13444 5264 13456
rect 4847 13416 5264 13444
rect 4847 13413 4859 13416
rect 4801 13407 4859 13413
rect 5258 13404 5264 13416
rect 5316 13444 5322 13456
rect 6546 13444 6552 13456
rect 5316 13416 6552 13444
rect 5316 13404 5322 13416
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 6825 13447 6883 13453
rect 6825 13413 6837 13447
rect 6871 13413 6883 13447
rect 6825 13407 6883 13413
rect 2866 13336 2872 13388
rect 2924 13336 2930 13388
rect 3050 13336 3056 13388
rect 3108 13336 3114 13388
rect 4982 13376 4988 13388
rect 4448 13348 4988 13376
rect 4448 13317 4476 13348
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 5810 13376 5816 13388
rect 5399 13348 5816 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 6840 13376 6868 13407
rect 7742 13404 7748 13456
rect 7800 13444 7806 13456
rect 7800 13416 8616 13444
rect 7800 13404 7806 13416
rect 6196 13348 6868 13376
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 5629 13311 5687 13317
rect 4755 13280 5304 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 2777 13243 2835 13249
rect 2777 13209 2789 13243
rect 2823 13240 2835 13243
rect 3234 13240 3240 13252
rect 2823 13212 3240 13240
rect 2823 13209 2835 13212
rect 2777 13203 2835 13209
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 3973 13243 4031 13249
rect 3973 13209 3985 13243
rect 4019 13209 4031 13243
rect 3973 13203 4031 13209
rect 3786 13132 3792 13184
rect 3844 13132 3850 13184
rect 3988 13172 4016 13203
rect 4154 13200 4160 13252
rect 4212 13200 4218 13252
rect 4448 13240 4476 13271
rect 5169 13243 5227 13249
rect 5169 13240 5181 13243
rect 4448 13212 5181 13240
rect 5169 13209 5181 13212
rect 5215 13209 5227 13243
rect 5169 13203 5227 13209
rect 5276 13240 5304 13280
rect 5629 13277 5641 13311
rect 5675 13308 5687 13311
rect 5718 13308 5724 13320
rect 5675 13280 5724 13308
rect 5675 13277 5687 13280
rect 5629 13271 5687 13277
rect 5718 13268 5724 13280
rect 5776 13308 5782 13320
rect 5905 13311 5963 13317
rect 5905 13308 5917 13311
rect 5776 13280 5917 13308
rect 5776 13268 5782 13280
rect 5905 13277 5917 13280
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 6196 13308 6224 13348
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7374 13376 7380 13388
rect 7156 13348 7380 13376
rect 7156 13336 7162 13348
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 6135 13280 6224 13308
rect 6273 13311 6331 13317
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 6273 13277 6285 13311
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 5994 13240 6000 13252
rect 5276 13212 6000 13240
rect 4522 13172 4528 13184
rect 3988 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 4706 13172 4712 13184
rect 4663 13144 4712 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4969 13175 5027 13181
rect 4969 13141 4981 13175
rect 5015 13172 5027 13175
rect 5276 13172 5304 13212
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 6178 13200 6184 13252
rect 6236 13240 6242 13252
rect 6288 13240 6316 13271
rect 6362 13268 6368 13320
rect 6420 13268 6426 13320
rect 6546 13268 6552 13320
rect 6604 13268 6610 13320
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 7285 13311 7343 13317
rect 7285 13308 7297 13311
rect 7064 13280 7297 13308
rect 7064 13268 7070 13280
rect 7285 13277 7297 13280
rect 7331 13308 7343 13311
rect 7466 13308 7472 13320
rect 7331 13280 7472 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 7466 13268 7472 13280
rect 7524 13308 7530 13320
rect 8021 13311 8079 13317
rect 8021 13308 8033 13311
rect 7524 13280 8033 13308
rect 7524 13268 7530 13280
rect 8021 13277 8033 13280
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 8294 13268 8300 13320
rect 8352 13268 8358 13320
rect 8478 13268 8484 13320
rect 8536 13268 8542 13320
rect 6822 13240 6828 13252
rect 6236 13212 6828 13240
rect 6236 13200 6242 13212
rect 6822 13200 6828 13212
rect 6880 13200 6886 13252
rect 7742 13200 7748 13252
rect 7800 13240 7806 13252
rect 7837 13243 7895 13249
rect 7837 13240 7849 13243
rect 7800 13212 7849 13240
rect 7800 13200 7806 13212
rect 7837 13209 7849 13212
rect 7883 13209 7895 13243
rect 7837 13203 7895 13209
rect 7926 13200 7932 13252
rect 7984 13240 7990 13252
rect 8389 13243 8447 13249
rect 8389 13240 8401 13243
rect 7984 13212 8401 13240
rect 7984 13200 7990 13212
rect 8389 13209 8401 13212
rect 8435 13209 8447 13243
rect 8389 13203 8447 13209
rect 5015 13144 5304 13172
rect 5015 13141 5027 13144
rect 4969 13135 5027 13141
rect 5350 13132 5356 13184
rect 5408 13132 5414 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 6457 13175 6515 13181
rect 6457 13172 6469 13175
rect 5500 13144 6469 13172
rect 5500 13132 5506 13144
rect 6457 13141 6469 13144
rect 6503 13141 6515 13175
rect 6457 13135 6515 13141
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 8018 13172 8024 13184
rect 7248 13144 8024 13172
rect 7248 13132 7254 13144
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8202 13132 8208 13184
rect 8260 13132 8266 13184
rect 8588 13172 8616 13416
rect 9214 13404 9220 13456
rect 9272 13444 9278 13456
rect 10686 13444 10692 13456
rect 9272 13416 10692 13444
rect 9272 13404 9278 13416
rect 9324 13385 9352 13416
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 9309 13379 9367 13385
rect 9309 13345 9321 13379
rect 9355 13345 9367 13379
rect 9309 13339 9367 13345
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 9631 13348 10824 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 8662 13268 8668 13320
rect 8720 13268 8726 13320
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9398 13308 9404 13320
rect 9263 13280 9404 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 10134 13268 10140 13320
rect 10192 13268 10198 13320
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13308 10287 13311
rect 10505 13311 10563 13317
rect 10275 13280 10456 13308
rect 10275 13277 10287 13280
rect 10229 13271 10287 13277
rect 8680 13240 8708 13268
rect 10318 13240 10324 13252
rect 8680 13212 10324 13240
rect 10318 13200 10324 13212
rect 10376 13200 10382 13252
rect 9950 13172 9956 13184
rect 8588 13144 9956 13172
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 10428 13172 10456 13280
rect 10505 13277 10517 13311
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 10520 13240 10548 13271
rect 10594 13268 10600 13320
rect 10652 13268 10658 13320
rect 10796 13317 10824 13348
rect 14642 13336 14648 13388
rect 14700 13376 14706 13388
rect 16025 13379 16083 13385
rect 16025 13376 16037 13379
rect 14700 13348 16037 13376
rect 14700 13336 14706 13348
rect 16025 13345 16037 13348
rect 16071 13345 16083 13379
rect 16592 13376 16620 13475
rect 17126 13472 17132 13484
rect 17184 13512 17190 13524
rect 19334 13512 19340 13524
rect 17184 13484 19340 13512
rect 17184 13472 17190 13484
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 20162 13472 20168 13524
rect 20220 13512 20226 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 20220 13484 20269 13512
rect 20220 13472 20226 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 20257 13475 20315 13481
rect 22738 13472 22744 13524
rect 22796 13512 22802 13524
rect 24486 13512 24492 13524
rect 22796 13484 24492 13512
rect 22796 13472 22802 13484
rect 24486 13472 24492 13484
rect 24544 13472 24550 13524
rect 26418 13472 26424 13524
rect 26476 13472 26482 13524
rect 28994 13472 29000 13524
rect 29052 13512 29058 13524
rect 29549 13515 29607 13521
rect 29549 13512 29561 13515
rect 29052 13484 29561 13512
rect 29052 13472 29058 13484
rect 29549 13481 29561 13484
rect 29595 13481 29607 13515
rect 29549 13475 29607 13481
rect 30282 13472 30288 13524
rect 30340 13472 30346 13524
rect 30558 13472 30564 13524
rect 30616 13512 30622 13524
rect 31386 13512 31392 13524
rect 30616 13484 31392 13512
rect 30616 13472 30622 13484
rect 31386 13472 31392 13484
rect 31444 13472 31450 13524
rect 33137 13515 33195 13521
rect 33137 13481 33149 13515
rect 33183 13512 33195 13515
rect 33226 13512 33232 13524
rect 33183 13484 33232 13512
rect 33183 13481 33195 13484
rect 33137 13475 33195 13481
rect 33226 13472 33232 13484
rect 33284 13472 33290 13524
rect 34606 13472 34612 13524
rect 34664 13512 34670 13524
rect 34790 13512 34796 13524
rect 34664 13484 34796 13512
rect 34664 13472 34670 13484
rect 34790 13472 34796 13484
rect 34848 13472 34854 13524
rect 35250 13472 35256 13524
rect 35308 13512 35314 13524
rect 35802 13512 35808 13524
rect 35308 13484 35808 13512
rect 35308 13472 35314 13484
rect 35802 13472 35808 13484
rect 35860 13472 35866 13524
rect 16945 13447 17003 13453
rect 16945 13413 16957 13447
rect 16991 13444 17003 13447
rect 17586 13444 17592 13456
rect 16991 13416 17592 13444
rect 16991 13413 17003 13416
rect 16945 13407 17003 13413
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 19518 13404 19524 13456
rect 19576 13404 19582 13456
rect 19613 13447 19671 13453
rect 19613 13413 19625 13447
rect 19659 13444 19671 13447
rect 19886 13444 19892 13456
rect 19659 13416 19892 13444
rect 19659 13413 19671 13416
rect 19613 13407 19671 13413
rect 19886 13404 19892 13416
rect 19944 13404 19950 13456
rect 20073 13447 20131 13453
rect 20073 13413 20085 13447
rect 20119 13444 20131 13447
rect 20119 13416 20208 13444
rect 20119 13413 20131 13416
rect 20073 13407 20131 13413
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 16025 13339 16083 13345
rect 16224 13348 16620 13376
rect 16960 13348 17785 13376
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 12894 13308 12900 13320
rect 12851 13280 12900 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 12894 13268 12900 13280
rect 12952 13308 12958 13320
rect 13630 13308 13636 13320
rect 12952 13280 13636 13308
rect 12952 13268 12958 13280
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14056 13280 14412 13308
rect 14056 13268 14062 13280
rect 11514 13240 11520 13252
rect 10520 13212 11520 13240
rect 11514 13200 11520 13212
rect 11572 13200 11578 13252
rect 12989 13243 13047 13249
rect 12989 13209 13001 13243
rect 13035 13240 13047 13243
rect 14274 13240 14280 13252
rect 13035 13212 14280 13240
rect 13035 13209 13047 13212
rect 12989 13203 13047 13209
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 14384 13240 14412 13280
rect 14458 13268 14464 13320
rect 14516 13268 14522 13320
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13308 14795 13311
rect 15746 13308 15752 13320
rect 14783 13280 15752 13308
rect 14783 13277 14795 13280
rect 14737 13271 14795 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16224 13317 16252 13348
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 16482 13268 16488 13320
rect 16540 13268 16546 13320
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 16761 13311 16819 13317
rect 16761 13308 16773 13311
rect 16632 13280 16773 13308
rect 16632 13268 16638 13280
rect 16761 13277 16773 13280
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 16393 13243 16451 13249
rect 14384 13212 15056 13240
rect 15028 13184 15056 13212
rect 16393 13209 16405 13243
rect 16439 13240 16451 13243
rect 16960 13240 16988 13348
rect 17773 13345 17785 13348
rect 17819 13376 17831 13379
rect 17954 13376 17960 13388
rect 17819 13348 17960 13376
rect 17819 13345 17831 13348
rect 17773 13339 17831 13345
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13376 19763 13379
rect 19751 13348 19840 13376
rect 19751 13345 19763 13348
rect 19705 13339 19763 13345
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13308 17095 13311
rect 17402 13308 17408 13320
rect 17083 13280 17408 13308
rect 17083 13277 17095 13280
rect 17037 13271 17095 13277
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 17586 13268 17592 13320
rect 17644 13268 17650 13320
rect 17681 13311 17739 13317
rect 17681 13277 17693 13311
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13308 17923 13311
rect 18322 13308 18328 13320
rect 17911 13280 18328 13308
rect 17911 13277 17923 13280
rect 17865 13271 17923 13277
rect 16439 13212 16988 13240
rect 16439 13209 16451 13212
rect 16393 13203 16451 13209
rect 17494 13200 17500 13252
rect 17552 13240 17558 13252
rect 17696 13240 17724 13271
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 17552 13212 17724 13240
rect 17552 13200 17558 13212
rect 19150 13200 19156 13252
rect 19208 13240 19214 13252
rect 19334 13240 19340 13252
rect 19208 13212 19340 13240
rect 19208 13200 19214 13212
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 19812 13240 19840 13348
rect 20180 13320 20208 13416
rect 21542 13404 21548 13456
rect 21600 13444 21606 13456
rect 26237 13447 26295 13453
rect 26237 13444 26249 13447
rect 21600 13416 26249 13444
rect 21600 13404 21606 13416
rect 26237 13413 26249 13416
rect 26283 13413 26295 13447
rect 31846 13444 31852 13456
rect 26237 13407 26295 13413
rect 29840 13416 31852 13444
rect 20530 13336 20536 13388
rect 20588 13336 20594 13388
rect 29638 13336 29644 13388
rect 29696 13376 29702 13388
rect 29840 13385 29868 13416
rect 31846 13404 31852 13416
rect 31904 13404 31910 13456
rect 34054 13444 34060 13456
rect 32416 13416 34060 13444
rect 29733 13379 29791 13385
rect 29733 13376 29745 13379
rect 29696 13348 29745 13376
rect 29696 13336 29702 13348
rect 29733 13345 29745 13348
rect 29779 13345 29791 13379
rect 29733 13339 29791 13345
rect 29825 13379 29883 13385
rect 29825 13345 29837 13379
rect 29871 13345 29883 13379
rect 29825 13339 29883 13345
rect 30009 13379 30067 13385
rect 30009 13345 30021 13379
rect 30055 13376 30067 13379
rect 30282 13376 30288 13388
rect 30055 13348 30288 13376
rect 30055 13345 30067 13348
rect 30009 13339 30067 13345
rect 30282 13336 30288 13348
rect 30340 13336 30346 13388
rect 30650 13336 30656 13388
rect 30708 13376 30714 13388
rect 31570 13376 31576 13388
rect 30708 13348 31576 13376
rect 30708 13336 30714 13348
rect 31570 13336 31576 13348
rect 31628 13376 31634 13388
rect 32416 13376 32444 13416
rect 34054 13404 34060 13416
rect 34112 13404 34118 13456
rect 31628 13348 32444 13376
rect 31628 13336 31634 13348
rect 32490 13336 32496 13388
rect 32548 13336 32554 13388
rect 19886 13268 19892 13320
rect 19944 13308 19950 13320
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 19944 13280 19993 13308
rect 19944 13268 19950 13280
rect 19981 13277 19993 13280
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 20162 13268 20168 13320
rect 20220 13268 20226 13320
rect 20257 13311 20315 13317
rect 20257 13277 20269 13311
rect 20303 13277 20315 13311
rect 20257 13271 20315 13277
rect 19720 13212 19840 13240
rect 20272 13240 20300 13271
rect 20346 13268 20352 13320
rect 20404 13268 20410 13320
rect 20438 13240 20444 13252
rect 20272 13212 20444 13240
rect 19720 13184 19748 13212
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 20548 13249 20576 13336
rect 29917 13311 29975 13317
rect 29917 13308 29929 13311
rect 28966 13280 29929 13308
rect 20533 13243 20591 13249
rect 20533 13209 20545 13243
rect 20579 13209 20591 13243
rect 26605 13243 26663 13249
rect 26605 13240 26617 13243
rect 20533 13203 20591 13209
rect 20916 13212 26617 13240
rect 10597 13175 10655 13181
rect 10597 13172 10609 13175
rect 10428 13144 10609 13172
rect 10597 13141 10609 13144
rect 10643 13141 10655 13175
rect 10597 13135 10655 13141
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12802 13172 12808 13184
rect 12575 13144 12808 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13170 13132 13176 13184
rect 13228 13172 13234 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 13228 13144 14933 13172
rect 13228 13132 13234 13144
rect 14921 13141 14933 13144
rect 14967 13141 14979 13175
rect 14921 13135 14979 13141
rect 15010 13132 15016 13184
rect 15068 13172 15074 13184
rect 17405 13175 17463 13181
rect 17405 13172 17417 13175
rect 15068 13144 17417 13172
rect 15068 13132 15074 13144
rect 17405 13141 17417 13144
rect 17451 13141 17463 13175
rect 17405 13135 17463 13141
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 18932 13144 19257 13172
rect 18932 13132 18938 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 19702 13132 19708 13184
rect 19760 13132 19766 13184
rect 19889 13175 19947 13181
rect 19889 13141 19901 13175
rect 19935 13172 19947 13175
rect 20806 13172 20812 13184
rect 19935 13144 20812 13172
rect 19935 13141 19947 13144
rect 19889 13135 19947 13141
rect 20806 13132 20812 13144
rect 20864 13172 20870 13184
rect 20916 13172 20944 13212
rect 26605 13209 26617 13212
rect 26651 13209 26663 13243
rect 26605 13203 26663 13209
rect 28810 13200 28816 13252
rect 28868 13240 28874 13252
rect 28966 13240 28994 13280
rect 29917 13277 29929 13280
rect 29963 13277 29975 13311
rect 30469 13311 30527 13317
rect 30469 13308 30481 13311
rect 29917 13271 29975 13277
rect 30024 13280 30481 13308
rect 28868 13212 28994 13240
rect 28868 13200 28874 13212
rect 29638 13200 29644 13252
rect 29696 13240 29702 13252
rect 30024 13240 30052 13280
rect 30469 13277 30481 13280
rect 30515 13308 30527 13311
rect 30515 13280 30788 13308
rect 30515 13277 30527 13280
rect 30469 13271 30527 13277
rect 29696 13212 30052 13240
rect 29696 13200 29702 13212
rect 30098 13200 30104 13252
rect 30156 13240 30162 13252
rect 30282 13240 30288 13252
rect 30156 13212 30288 13240
rect 30156 13200 30162 13212
rect 30282 13200 30288 13212
rect 30340 13200 30346 13252
rect 30561 13243 30619 13249
rect 30561 13209 30573 13243
rect 30607 13209 30619 13243
rect 30561 13203 30619 13209
rect 20864 13144 20944 13172
rect 26421 13175 26479 13181
rect 20864 13132 20870 13144
rect 26421 13141 26433 13175
rect 26467 13172 26479 13175
rect 26970 13172 26976 13184
rect 26467 13144 26976 13172
rect 26467 13141 26479 13144
rect 26421 13135 26479 13141
rect 26970 13132 26976 13144
rect 27028 13172 27034 13184
rect 27338 13172 27344 13184
rect 27028 13144 27344 13172
rect 27028 13132 27034 13144
rect 27338 13132 27344 13144
rect 27396 13132 27402 13184
rect 30576 13172 30604 13203
rect 30650 13200 30656 13252
rect 30708 13200 30714 13252
rect 30760 13240 30788 13280
rect 30834 13268 30840 13320
rect 30892 13268 30898 13320
rect 32306 13268 32312 13320
rect 32364 13308 32370 13320
rect 32631 13311 32689 13317
rect 32631 13308 32643 13311
rect 32364 13280 32643 13308
rect 32364 13268 32370 13280
rect 32631 13277 32643 13280
rect 32677 13277 32689 13311
rect 32631 13271 32689 13277
rect 32950 13268 32956 13320
rect 33008 13268 33014 13320
rect 33594 13268 33600 13320
rect 33652 13308 33658 13320
rect 34514 13308 34520 13320
rect 33652 13280 34520 13308
rect 33652 13268 33658 13280
rect 34514 13268 34520 13280
rect 34572 13268 34578 13320
rect 31018 13240 31024 13252
rect 30760 13212 31024 13240
rect 31018 13200 31024 13212
rect 31076 13240 31082 13252
rect 31754 13240 31760 13252
rect 31076 13212 31760 13240
rect 31076 13200 31082 13212
rect 31754 13200 31760 13212
rect 31812 13200 31818 13252
rect 32766 13200 32772 13252
rect 32824 13200 32830 13252
rect 32858 13200 32864 13252
rect 32916 13200 32922 13252
rect 31478 13172 31484 13184
rect 30576 13144 31484 13172
rect 31478 13132 31484 13144
rect 31536 13132 31542 13184
rect 1104 13082 36432 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 36432 13082
rect 1104 13008 36432 13030
rect 3142 12928 3148 12980
rect 3200 12928 3206 12980
rect 3234 12928 3240 12980
rect 3292 12928 3298 12980
rect 5258 12968 5264 12980
rect 4356 12940 5264 12968
rect 4356 12909 4384 12940
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 5810 12968 5816 12980
rect 5644 12940 5816 12968
rect 4341 12903 4399 12909
rect 4341 12869 4353 12903
rect 4387 12869 4399 12903
rect 4341 12863 4399 12869
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 4525 12903 4583 12909
rect 4525 12900 4537 12903
rect 4488 12872 4537 12900
rect 4488 12860 4494 12872
rect 4525 12869 4537 12872
rect 4571 12900 4583 12903
rect 4571 12872 5580 12900
rect 4571 12869 4583 12872
rect 4525 12863 4583 12869
rect 2774 12792 2780 12844
rect 2832 12792 2838 12844
rect 3602 12792 3608 12844
rect 3660 12792 3666 12844
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4798 12841 4804 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 4120 12804 4169 12832
rect 4120 12792 4126 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 4796 12795 4804 12841
rect 4798 12792 4804 12795
rect 4856 12792 4862 12844
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 1394 12724 1400 12776
rect 1452 12724 1458 12776
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 3694 12724 3700 12776
rect 3752 12724 3758 12776
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 4706 12764 4712 12776
rect 3927 12736 4712 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 3050 12656 3056 12708
rect 3108 12696 3114 12708
rect 3896 12696 3924 12727
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 3108 12668 3924 12696
rect 3108 12656 3114 12668
rect 4522 12656 4528 12708
rect 4580 12696 4586 12708
rect 4908 12696 4936 12795
rect 4982 12792 4988 12844
rect 5040 12792 5046 12844
rect 5166 12832 5172 12844
rect 5127 12804 5172 12832
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 5423 12835 5481 12841
rect 5423 12832 5435 12835
rect 5307 12804 5435 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5423 12801 5435 12804
rect 5469 12801 5481 12835
rect 5423 12795 5481 12801
rect 5552 12773 5580 12872
rect 5644 12832 5672 12940
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 6914 12928 6920 12980
rect 6972 12928 6978 12980
rect 7009 12971 7067 12977
rect 7009 12937 7021 12971
rect 7055 12968 7067 12971
rect 7190 12968 7196 12980
rect 7055 12940 7196 12968
rect 7055 12937 7067 12940
rect 7009 12931 7067 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 8202 12928 8208 12980
rect 8260 12928 8266 12980
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 8849 12971 8907 12977
rect 8849 12968 8861 12971
rect 8628 12940 8861 12968
rect 8628 12928 8634 12940
rect 8849 12937 8861 12940
rect 8895 12968 8907 12971
rect 8938 12968 8944 12980
rect 8895 12940 8944 12968
rect 8895 12937 8907 12940
rect 8849 12931 8907 12937
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 9674 12928 9680 12980
rect 9732 12928 9738 12980
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 11422 12968 11428 12980
rect 10376 12940 11428 12968
rect 10376 12928 10382 12940
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 14274 12928 14280 12980
rect 14332 12928 14338 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19521 12971 19579 12977
rect 19521 12968 19533 12971
rect 19392 12940 19533 12968
rect 19392 12928 19398 12940
rect 19521 12937 19533 12940
rect 19567 12937 19579 12971
rect 19521 12931 19579 12937
rect 21928 12940 22232 12968
rect 6638 12900 6644 12912
rect 5828 12872 6644 12900
rect 5828 12844 5856 12872
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 6932 12900 6960 12928
rect 6932 12872 7144 12900
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5644 12804 5733 12832
rect 5721 12801 5733 12804
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 5810 12792 5816 12844
rect 5868 12792 5874 12844
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 6454 12832 6460 12844
rect 6043 12804 6460 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12764 5595 12767
rect 6362 12764 6368 12776
rect 5583 12736 6368 12764
rect 5583 12733 5595 12736
rect 5537 12727 5595 12733
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 7116 12773 7144 12872
rect 8018 12860 8024 12912
rect 8076 12900 8082 12912
rect 8220 12900 8248 12928
rect 8076 12872 8156 12900
rect 8220 12872 8432 12900
rect 8076 12860 8082 12872
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 7561 12835 7619 12841
rect 7561 12832 7573 12835
rect 7340 12804 7573 12832
rect 7340 12792 7346 12804
rect 7561 12801 7573 12804
rect 7607 12801 7619 12835
rect 8128 12832 8156 12872
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 8128 12804 8217 12832
rect 7561 12795 7619 12801
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 7190 12764 7196 12776
rect 7147 12736 7196 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 4580 12668 4936 12696
rect 4580 12656 4586 12668
rect 3878 12588 3884 12640
rect 3936 12628 3942 12640
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 3936 12600 4629 12628
rect 3936 12588 3942 12600
rect 4617 12597 4629 12600
rect 4663 12597 4675 12631
rect 4908 12628 4936 12668
rect 5353 12699 5411 12705
rect 5353 12665 5365 12699
rect 5399 12696 5411 12699
rect 6914 12696 6920 12708
rect 5399 12668 6920 12696
rect 5399 12665 5411 12668
rect 5353 12659 5411 12665
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 7576 12696 7604 12795
rect 8294 12792 8300 12844
rect 8352 12792 8358 12844
rect 8404 12841 8432 12872
rect 8478 12860 8484 12912
rect 8536 12860 8542 12912
rect 9033 12903 9091 12909
rect 9033 12869 9045 12903
rect 9079 12900 9091 12903
rect 9582 12900 9588 12912
rect 9079 12872 9588 12900
rect 9079 12869 9091 12872
rect 9033 12863 9091 12869
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 10137 12903 10195 12909
rect 10137 12900 10149 12903
rect 9640 12872 10149 12900
rect 9640 12860 9646 12872
rect 10137 12869 10149 12872
rect 10183 12900 10195 12903
rect 10502 12900 10508 12912
rect 10183 12872 10508 12900
rect 10183 12869 10195 12872
rect 10137 12863 10195 12869
rect 10502 12860 10508 12872
rect 10560 12860 10566 12912
rect 14182 12860 14188 12912
rect 14240 12900 14246 12912
rect 14737 12903 14795 12909
rect 14737 12900 14749 12903
rect 14240 12872 14749 12900
rect 14240 12860 14246 12872
rect 14737 12869 14749 12872
rect 14783 12869 14795 12903
rect 14737 12863 14795 12869
rect 16482 12860 16488 12912
rect 16540 12900 16546 12912
rect 21928 12900 21956 12940
rect 16540 12872 21956 12900
rect 16540 12860 16546 12872
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12801 8447 12835
rect 8496 12832 8524 12860
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 8496 12804 8585 12832
rect 8389 12795 8447 12801
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12832 8723 12835
rect 9122 12832 9128 12844
rect 8711 12804 9128 12832
rect 8711 12801 8723 12804
rect 8665 12795 8723 12801
rect 9122 12792 9128 12804
rect 9180 12832 9186 12844
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 9180 12804 9321 12832
rect 9180 12792 9186 12804
rect 9309 12801 9321 12804
rect 9355 12801 9367 12835
rect 9309 12795 9367 12801
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10042 12832 10048 12844
rect 9999 12804 10048 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12832 10287 12835
rect 10686 12832 10692 12844
rect 10275 12804 10692 12832
rect 10275 12801 10287 12804
rect 10229 12795 10287 12801
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12832 14519 12835
rect 14507 12804 14780 12832
rect 14507 12801 14519 12804
rect 14461 12795 14519 12801
rect 7742 12724 7748 12776
rect 7800 12764 7806 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7800 12736 7849 12764
rect 7800 12724 7806 12736
rect 7837 12733 7849 12736
rect 7883 12764 7895 12767
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7883 12736 7941 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 7929 12733 7941 12736
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 8812 12736 9229 12764
rect 8812 12724 8818 12736
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 10318 12724 10324 12776
rect 10376 12724 10382 12776
rect 10594 12724 10600 12776
rect 10652 12724 10658 12776
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 14424 12736 14565 12764
rect 14424 12724 14430 12736
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 14752 12764 14780 12804
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 14884 12804 15025 12832
rect 14884 12792 14890 12804
rect 15013 12801 15025 12804
rect 15059 12801 15071 12835
rect 15013 12795 15071 12801
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 15838 12832 15844 12844
rect 15611 12804 15844 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 19702 12792 19708 12844
rect 19760 12792 19766 12844
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 20162 12832 20168 12844
rect 19935 12804 20168 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 21726 12792 21732 12844
rect 21784 12832 21790 12844
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 21784 12804 21833 12832
rect 21784 12792 21790 12804
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21968 12804 22017 12832
rect 21968 12792 21974 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22094 12792 22100 12844
rect 22152 12792 22158 12844
rect 14918 12764 14924 12776
rect 14752 12736 14924 12764
rect 14553 12727 14611 12733
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 15746 12724 15752 12776
rect 15804 12724 15810 12776
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 22204 12764 22232 12940
rect 22278 12928 22284 12980
rect 22336 12928 22342 12980
rect 24394 12968 24400 12980
rect 22848 12940 23152 12968
rect 22848 12909 22876 12940
rect 22833 12903 22891 12909
rect 22833 12869 22845 12903
rect 22879 12869 22891 12903
rect 22833 12863 22891 12869
rect 23014 12860 23020 12912
rect 23072 12909 23078 12912
rect 23072 12903 23091 12909
rect 23079 12869 23091 12903
rect 23124 12900 23152 12940
rect 23492 12940 24400 12968
rect 23492 12912 23520 12940
rect 24394 12928 24400 12940
rect 24452 12928 24458 12980
rect 29454 12928 29460 12980
rect 29512 12968 29518 12980
rect 32858 12968 32864 12980
rect 29512 12940 32864 12968
rect 29512 12928 29518 12940
rect 32858 12928 32864 12940
rect 32916 12928 32922 12980
rect 23474 12900 23480 12912
rect 23124 12872 23480 12900
rect 23072 12863 23091 12869
rect 23072 12860 23078 12863
rect 23474 12860 23480 12872
rect 23532 12860 23538 12912
rect 22922 12792 22928 12844
rect 22980 12832 22986 12844
rect 24029 12835 24087 12841
rect 24029 12832 24041 12835
rect 22980 12804 24041 12832
rect 22980 12792 22986 12804
rect 24029 12801 24041 12804
rect 24075 12801 24087 12835
rect 24029 12795 24087 12801
rect 32674 12792 32680 12844
rect 32732 12832 32738 12844
rect 32858 12832 32864 12844
rect 32732 12804 32864 12832
rect 32732 12792 32738 12804
rect 32858 12792 32864 12804
rect 32916 12792 32922 12844
rect 25038 12764 25044 12776
rect 17552 12736 22140 12764
rect 22204 12736 25044 12764
rect 17552 12724 17558 12736
rect 8294 12696 8300 12708
rect 7576 12668 8300 12696
rect 8294 12656 8300 12668
rect 8352 12696 8358 12708
rect 8846 12696 8852 12708
rect 8352 12668 8852 12696
rect 8352 12656 8358 12668
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 9674 12696 9680 12708
rect 8956 12668 9680 12696
rect 5442 12628 5448 12640
rect 4908 12600 5448 12628
rect 4617 12591 4675 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 5626 12588 5632 12640
rect 5684 12588 5690 12640
rect 6178 12588 6184 12640
rect 6236 12628 6242 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6236 12600 6561 12628
rect 6236 12588 6242 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 7374 12588 7380 12640
rect 7432 12588 7438 12640
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 7926 12628 7932 12640
rect 7791 12600 7932 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 8956 12628 8984 12668
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 10410 12656 10416 12708
rect 10468 12696 10474 12708
rect 15013 12699 15071 12705
rect 15013 12696 15025 12699
rect 10468 12668 15025 12696
rect 10468 12656 10474 12668
rect 15013 12665 15025 12668
rect 15059 12665 15071 12699
rect 15013 12659 15071 12665
rect 17402 12656 17408 12708
rect 17460 12696 17466 12708
rect 19334 12696 19340 12708
rect 17460 12668 19340 12696
rect 17460 12656 17466 12668
rect 19334 12656 19340 12668
rect 19392 12656 19398 12708
rect 22112 12696 22140 12736
rect 25038 12724 25044 12736
rect 25096 12724 25102 12776
rect 22462 12696 22468 12708
rect 22112 12668 22468 12696
rect 22462 12656 22468 12668
rect 22520 12656 22526 12708
rect 26602 12696 26608 12708
rect 23032 12668 26608 12696
rect 8260 12600 8984 12628
rect 8260 12588 8266 12600
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 9769 12631 9827 12637
rect 9769 12628 9781 12631
rect 9180 12600 9781 12628
rect 9180 12588 9186 12600
rect 9769 12597 9781 12600
rect 9815 12597 9827 12631
rect 9769 12591 9827 12597
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10778 12628 10784 12640
rect 10008 12600 10784 12628
rect 10008 12588 10014 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 14642 12588 14648 12640
rect 14700 12588 14706 12640
rect 19889 12631 19947 12637
rect 19889 12597 19901 12631
rect 19935 12628 19947 12631
rect 20070 12628 20076 12640
rect 19935 12600 20076 12628
rect 19935 12597 19947 12600
rect 19889 12591 19947 12597
rect 20070 12588 20076 12600
rect 20128 12628 20134 12640
rect 20346 12628 20352 12640
rect 20128 12600 20352 12628
rect 20128 12588 20134 12600
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 21818 12628 21824 12640
rect 20588 12600 21824 12628
rect 20588 12588 20594 12600
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22370 12628 22376 12640
rect 22152 12600 22376 12628
rect 22152 12588 22158 12600
rect 22370 12588 22376 12600
rect 22428 12628 22434 12640
rect 23032 12637 23060 12668
rect 26602 12656 26608 12668
rect 26660 12656 26666 12708
rect 23017 12631 23075 12637
rect 23017 12628 23029 12631
rect 22428 12600 23029 12628
rect 22428 12588 22434 12600
rect 23017 12597 23029 12600
rect 23063 12597 23075 12631
rect 23017 12591 23075 12597
rect 23198 12588 23204 12640
rect 23256 12588 23262 12640
rect 23566 12588 23572 12640
rect 23624 12628 23630 12640
rect 23937 12631 23995 12637
rect 23937 12628 23949 12631
rect 23624 12600 23949 12628
rect 23624 12588 23630 12600
rect 23937 12597 23949 12600
rect 23983 12628 23995 12631
rect 24302 12628 24308 12640
rect 23983 12600 24308 12628
rect 23983 12597 23995 12600
rect 23937 12591 23995 12597
rect 24302 12588 24308 12600
rect 24360 12588 24366 12640
rect 26418 12588 26424 12640
rect 26476 12628 26482 12640
rect 28810 12628 28816 12640
rect 26476 12600 28816 12628
rect 26476 12588 26482 12600
rect 28810 12588 28816 12600
rect 28868 12588 28874 12640
rect 29822 12588 29828 12640
rect 29880 12628 29886 12640
rect 32674 12628 32680 12640
rect 29880 12600 32680 12628
rect 29880 12588 29886 12600
rect 32674 12588 32680 12600
rect 32732 12588 32738 12640
rect 1104 12538 36432 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 36432 12538
rect 1104 12464 36432 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 2501 12427 2559 12433
rect 2501 12424 2513 12427
rect 1728 12396 2513 12424
rect 1728 12384 1734 12396
rect 2501 12393 2513 12396
rect 2547 12393 2559 12427
rect 2501 12387 2559 12393
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3660 12396 3801 12424
rect 3660 12384 3666 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 4246 12424 4252 12436
rect 3936 12396 4252 12424
rect 3936 12384 3942 12396
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 5902 12424 5908 12436
rect 5276 12396 5908 12424
rect 2958 12356 2964 12368
rect 2695 12328 2964 12356
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2406 12288 2412 12300
rect 2179 12260 2412 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 2038 12180 2044 12232
rect 2096 12180 2102 12232
rect 2222 12180 2228 12232
rect 2280 12220 2286 12232
rect 2695 12229 2723 12328
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 3142 12316 3148 12368
rect 3200 12316 3206 12368
rect 4706 12316 4712 12368
rect 4764 12316 4770 12368
rect 3160 12288 3188 12316
rect 3694 12288 3700 12300
rect 2792 12260 3188 12288
rect 3252 12260 3700 12288
rect 2792 12229 2820 12260
rect 2680 12223 2738 12229
rect 2680 12220 2692 12223
rect 2280 12192 2692 12220
rect 2280 12180 2286 12192
rect 2680 12189 2692 12192
rect 2726 12189 2738 12223
rect 2680 12183 2738 12189
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12189 2835 12223
rect 3050 12220 3056 12232
rect 3011 12192 3056 12220
rect 2777 12183 2835 12189
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 3142 12180 3148 12232
rect 3200 12180 3206 12232
rect 2866 12112 2872 12164
rect 2924 12112 2930 12164
rect 2409 12087 2467 12093
rect 2409 12053 2421 12087
rect 2455 12084 2467 12087
rect 3252 12084 3280 12260
rect 3694 12248 3700 12260
rect 3752 12248 3758 12300
rect 3786 12248 3792 12300
rect 3844 12288 3850 12300
rect 3973 12291 4031 12297
rect 3973 12288 3985 12291
rect 3844 12260 3985 12288
rect 3844 12248 3850 12260
rect 3973 12257 3985 12260
rect 4019 12257 4031 12291
rect 3973 12251 4031 12257
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12257 4215 12291
rect 4157 12251 4215 12257
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 3421 12223 3479 12229
rect 3421 12220 3433 12223
rect 3384 12192 3433 12220
rect 3384 12180 3390 12192
rect 3421 12189 3433 12192
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3602 12180 3608 12232
rect 3660 12180 3666 12232
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12189 4123 12223
rect 4172 12220 4200 12251
rect 4246 12248 4252 12300
rect 4304 12248 4310 12300
rect 4614 12288 4620 12300
rect 4540 12260 4620 12288
rect 4338 12220 4344 12232
rect 4172 12192 4344 12220
rect 4065 12183 4123 12189
rect 3513 12155 3571 12161
rect 3513 12121 3525 12155
rect 3559 12152 3571 12155
rect 4080 12152 4108 12183
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 4540 12229 4568 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12288 5227 12291
rect 5276 12288 5304 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7190 12424 7196 12436
rect 6972 12396 7196 12424
rect 6972 12384 6978 12396
rect 7190 12384 7196 12396
rect 7248 12424 7254 12436
rect 8018 12424 8024 12436
rect 7248 12396 8024 12424
rect 7248 12384 7254 12396
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8128 12396 8585 12424
rect 5442 12316 5448 12368
rect 5500 12356 5506 12368
rect 7377 12359 7435 12365
rect 5500 12328 5948 12356
rect 5500 12316 5506 12328
rect 5215 12260 5304 12288
rect 5215 12257 5227 12260
rect 5169 12251 5227 12257
rect 5718 12248 5724 12300
rect 5776 12248 5782 12300
rect 5920 12297 5948 12328
rect 6012 12328 6960 12356
rect 6012 12297 6040 12328
rect 6932 12300 6960 12328
rect 7377 12325 7389 12359
rect 7423 12356 7435 12359
rect 7558 12356 7564 12368
rect 7423 12328 7564 12356
rect 7423 12325 7435 12328
rect 7377 12319 7435 12325
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 7926 12356 7932 12368
rect 7668 12328 7932 12356
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12257 6055 12291
rect 5997 12251 6055 12257
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 6227 12260 6469 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 6914 12248 6920 12300
rect 6972 12248 6978 12300
rect 7193 12291 7251 12297
rect 7193 12257 7205 12291
rect 7239 12288 7251 12291
rect 7282 12288 7288 12300
rect 7239 12260 7288 12288
rect 7239 12257 7251 12260
rect 7193 12251 7251 12257
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 7668 12288 7696 12328
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 8128 12288 8156 12396
rect 8573 12393 8585 12396
rect 8619 12424 8631 12427
rect 8662 12424 8668 12436
rect 8619 12396 8668 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 10042 12424 10048 12436
rect 8812 12396 10048 12424
rect 8812 12384 8818 12396
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 10321 12427 10379 12433
rect 10321 12393 10333 12427
rect 10367 12424 10379 12427
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 10367 12396 10609 12424
rect 10367 12393 10379 12396
rect 10321 12387 10379 12393
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 10597 12387 10655 12393
rect 13078 12384 13084 12436
rect 13136 12384 13142 12436
rect 15378 12384 15384 12436
rect 15436 12384 15442 12436
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 15930 12424 15936 12436
rect 15620 12396 15936 12424
rect 15620 12384 15626 12396
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 17494 12384 17500 12436
rect 17552 12384 17558 12436
rect 18230 12384 18236 12436
rect 18288 12424 18294 12436
rect 18601 12427 18659 12433
rect 18601 12424 18613 12427
rect 18288 12396 18613 12424
rect 18288 12384 18294 12396
rect 18601 12393 18613 12396
rect 18647 12393 18659 12427
rect 18601 12387 18659 12393
rect 18785 12427 18843 12433
rect 18785 12393 18797 12427
rect 18831 12424 18843 12427
rect 18966 12424 18972 12436
rect 18831 12396 18972 12424
rect 18831 12393 18843 12396
rect 18785 12387 18843 12393
rect 18966 12384 18972 12396
rect 19024 12424 19030 12436
rect 21637 12427 21695 12433
rect 19024 12396 20300 12424
rect 19024 12384 19030 12396
rect 20272 12368 20300 12396
rect 21637 12393 21649 12427
rect 21683 12424 21695 12427
rect 21726 12424 21732 12436
rect 21683 12396 21732 12424
rect 21683 12393 21695 12396
rect 21637 12387 21695 12393
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 22462 12384 22468 12436
rect 22520 12424 22526 12436
rect 23845 12427 23903 12433
rect 23845 12424 23857 12427
rect 22520 12396 23857 12424
rect 22520 12384 22526 12396
rect 23845 12393 23857 12396
rect 23891 12393 23903 12427
rect 23845 12387 23903 12393
rect 23934 12384 23940 12436
rect 23992 12424 23998 12436
rect 24029 12427 24087 12433
rect 24029 12424 24041 12427
rect 23992 12396 24041 12424
rect 23992 12384 23998 12396
rect 24029 12393 24041 12396
rect 24075 12393 24087 12427
rect 24029 12387 24087 12393
rect 24578 12384 24584 12436
rect 24636 12424 24642 12436
rect 24765 12427 24823 12433
rect 24765 12424 24777 12427
rect 24636 12396 24777 12424
rect 24636 12384 24642 12396
rect 24765 12393 24777 12396
rect 24811 12393 24823 12427
rect 24765 12387 24823 12393
rect 25777 12427 25835 12433
rect 25777 12393 25789 12427
rect 25823 12424 25835 12427
rect 25958 12424 25964 12436
rect 25823 12396 25964 12424
rect 25823 12393 25835 12396
rect 25777 12387 25835 12393
rect 25958 12384 25964 12396
rect 26016 12384 26022 12436
rect 27614 12384 27620 12436
rect 27672 12384 27678 12436
rect 28074 12384 28080 12436
rect 28132 12384 28138 12436
rect 28350 12384 28356 12436
rect 28408 12424 28414 12436
rect 28408 12396 29960 12424
rect 28408 12384 28414 12396
rect 8202 12316 8208 12368
rect 8260 12316 8266 12368
rect 8478 12316 8484 12368
rect 8536 12356 8542 12368
rect 8536 12328 9444 12356
rect 8536 12316 8542 12328
rect 7576 12260 7696 12288
rect 7852 12260 8156 12288
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4890 12220 4896 12232
rect 4755 12192 4896 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 3559 12124 4108 12152
rect 3559 12121 3571 12124
rect 3513 12115 3571 12121
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4448 12152 4476 12183
rect 4212 12124 4476 12152
rect 4212 12112 4218 12124
rect 2455 12056 3280 12084
rect 2455 12053 2467 12056
rect 2409 12047 2467 12053
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 4540 12084 4568 12183
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 5442 12220 5448 12232
rect 5399 12192 5448 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 5276 12152 5304 12183
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 4672 12124 5304 12152
rect 4672 12112 4678 12124
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 5828 12152 5856 12183
rect 6546 12180 6552 12232
rect 6604 12180 6610 12232
rect 6730 12180 6736 12232
rect 6788 12220 6794 12232
rect 7469 12223 7527 12229
rect 6788 12192 6960 12220
rect 6788 12180 6794 12192
rect 5684 12124 6408 12152
rect 5684 12112 5690 12124
rect 3660 12056 4568 12084
rect 3660 12044 3666 12056
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 4985 12087 5043 12093
rect 4985 12084 4997 12087
rect 4856 12056 4997 12084
rect 4856 12044 4862 12056
rect 4985 12053 4997 12056
rect 5031 12053 5043 12087
rect 4985 12047 5043 12053
rect 6270 12044 6276 12096
rect 6328 12044 6334 12096
rect 6380 12084 6408 12124
rect 6454 12112 6460 12164
rect 6512 12152 6518 12164
rect 6932 12161 6960 12192
rect 7469 12189 7481 12223
rect 7515 12219 7527 12223
rect 7576 12219 7604 12260
rect 7515 12191 7604 12219
rect 7515 12189 7527 12191
rect 7469 12183 7527 12189
rect 7742 12180 7748 12232
rect 7800 12180 7806 12232
rect 7852 12229 7880 12260
rect 8662 12248 8668 12300
rect 8720 12288 8726 12300
rect 9416 12288 9444 12328
rect 9490 12316 9496 12368
rect 9548 12356 9554 12368
rect 9548 12328 9720 12356
rect 9548 12316 9554 12328
rect 8720 12260 9352 12288
rect 9416 12260 9536 12288
rect 8720 12248 8726 12260
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 6825 12155 6883 12161
rect 6825 12152 6837 12155
rect 6512 12124 6837 12152
rect 6512 12112 6518 12124
rect 6825 12121 6837 12124
rect 6871 12121 6883 12155
rect 6825 12115 6883 12121
rect 6917 12155 6975 12161
rect 6917 12121 6929 12155
rect 6963 12121 6975 12155
rect 7944 12152 7972 12183
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 9324 12229 9352 12260
rect 9125 12223 9183 12229
rect 8260 12192 8708 12220
rect 9125 12219 9137 12223
rect 8260 12180 8266 12192
rect 8570 12152 8576 12164
rect 6917 12115 6975 12121
rect 7024 12124 8576 12152
rect 6638 12084 6644 12096
rect 6380 12056 6644 12084
rect 6638 12044 6644 12056
rect 6696 12084 6702 12096
rect 7024 12084 7052 12124
rect 8570 12112 8576 12124
rect 8628 12112 8634 12164
rect 6696 12056 7052 12084
rect 6696 12044 6702 12056
rect 7466 12044 7472 12096
rect 7524 12044 7530 12096
rect 7558 12044 7564 12096
rect 7616 12044 7622 12096
rect 8680 12084 8708 12192
rect 9048 12191 9137 12219
rect 9048 12152 9076 12191
rect 9125 12189 9137 12191
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 9508 12229 9536 12260
rect 9692 12229 9720 12328
rect 10134 12316 10140 12368
rect 10192 12356 10198 12368
rect 10505 12359 10563 12365
rect 10505 12356 10517 12359
rect 10192 12328 10517 12356
rect 10192 12316 10198 12328
rect 10505 12325 10517 12328
rect 10551 12325 10563 12359
rect 10505 12319 10563 12325
rect 10870 12316 10876 12368
rect 10928 12356 10934 12368
rect 14093 12359 14151 12365
rect 14093 12356 14105 12359
rect 10928 12328 14105 12356
rect 10928 12316 10934 12328
rect 14093 12325 14105 12328
rect 14139 12325 14151 12359
rect 14093 12319 14151 12325
rect 14366 12316 14372 12368
rect 14424 12356 14430 12368
rect 14424 12328 15332 12356
rect 14424 12316 14430 12328
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 10100 12260 10977 12288
rect 10100 12248 10106 12260
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 15304 12297 15332 12328
rect 15746 12316 15752 12368
rect 15804 12356 15810 12368
rect 17681 12359 17739 12365
rect 17681 12356 17693 12359
rect 15804 12328 17693 12356
rect 15804 12316 15810 12328
rect 17681 12325 17693 12328
rect 17727 12356 17739 12359
rect 17770 12356 17776 12368
rect 17727 12328 17776 12356
rect 17727 12325 17739 12328
rect 17681 12319 17739 12325
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 18141 12359 18199 12365
rect 18141 12325 18153 12359
rect 18187 12356 18199 12359
rect 19150 12356 19156 12368
rect 18187 12328 19156 12356
rect 18187 12325 18199 12328
rect 18141 12319 18199 12325
rect 19150 12316 19156 12328
rect 19208 12316 19214 12368
rect 20254 12316 20260 12368
rect 20312 12356 20318 12368
rect 22094 12356 22100 12368
rect 20312 12328 22100 12356
rect 20312 12316 20318 12328
rect 22094 12316 22100 12328
rect 22152 12316 22158 12368
rect 22554 12316 22560 12368
rect 22612 12356 22618 12368
rect 22741 12359 22799 12365
rect 22741 12356 22753 12359
rect 22612 12328 22753 12356
rect 22612 12316 22618 12328
rect 22741 12325 22753 12328
rect 22787 12325 22799 12359
rect 22741 12319 22799 12325
rect 23293 12359 23351 12365
rect 23293 12325 23305 12359
rect 23339 12356 23351 12359
rect 23382 12356 23388 12368
rect 23339 12328 23388 12356
rect 23339 12325 23351 12328
rect 23293 12319 23351 12325
rect 23382 12316 23388 12328
rect 23440 12316 23446 12368
rect 25133 12359 25191 12365
rect 25133 12325 25145 12359
rect 25179 12356 25191 12359
rect 25179 12328 25452 12356
rect 25179 12325 25191 12328
rect 25133 12319 25191 12325
rect 15289 12291 15347 12297
rect 11756 12260 14688 12288
rect 11756 12248 11762 12260
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 9953 12223 10011 12229
rect 9953 12220 9965 12223
rect 9907 12192 9965 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 9953 12189 9965 12192
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 10192 12192 10333 12220
rect 10192 12180 10198 12192
rect 10321 12189 10333 12192
rect 10367 12220 10379 12223
rect 10594 12220 10600 12232
rect 10367 12192 10600 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12220 10839 12223
rect 10870 12220 10876 12232
rect 10827 12192 10876 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11606 12180 11612 12232
rect 11664 12180 11670 12232
rect 11803 12223 11861 12229
rect 11803 12189 11815 12223
rect 11849 12220 11861 12223
rect 12250 12220 12256 12232
rect 11849 12192 12256 12220
rect 11849 12189 11861 12192
rect 11803 12183 11861 12189
rect 12250 12180 12256 12192
rect 12308 12220 12314 12232
rect 12308 12192 12940 12220
rect 12308 12180 12314 12192
rect 10042 12152 10048 12164
rect 9048 12124 10048 12152
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 11701 12155 11759 12161
rect 11701 12152 11713 12155
rect 10152 12124 11713 12152
rect 10152 12084 10180 12124
rect 11701 12121 11713 12124
rect 11747 12121 11759 12155
rect 12912 12152 12940 12192
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 14660 12229 14688 12260
rect 15289 12257 15301 12291
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 17276 12260 18184 12288
rect 17276 12248 17282 12260
rect 18156 12232 18184 12260
rect 18322 12248 18328 12300
rect 18380 12248 18386 12300
rect 21082 12248 21088 12300
rect 21140 12288 21146 12300
rect 21177 12291 21235 12297
rect 21177 12288 21189 12291
rect 21140 12260 21189 12288
rect 21140 12248 21146 12260
rect 21177 12257 21189 12260
rect 21223 12257 21235 12291
rect 21177 12251 21235 12257
rect 21266 12248 21272 12300
rect 21324 12248 21330 12300
rect 23014 12288 23020 12300
rect 21376 12260 23020 12288
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 14645 12223 14703 12229
rect 13127 12192 14412 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13630 12152 13636 12164
rect 12912 12124 13636 12152
rect 11701 12115 11759 12121
rect 13630 12112 13636 12124
rect 13688 12112 13694 12164
rect 14274 12112 14280 12164
rect 14332 12112 14338 12164
rect 14384 12152 14412 12192
rect 14645 12189 14657 12223
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 15194 12180 15200 12232
rect 15252 12180 15258 12232
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 15519 12192 17785 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 18046 12180 18052 12232
rect 18104 12180 18110 12232
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 18196 12192 18245 12220
rect 18196 12180 18202 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12220 18567 12223
rect 19058 12220 19064 12232
rect 18555 12192 19064 12220
rect 18555 12189 18567 12192
rect 18509 12183 18567 12189
rect 19058 12180 19064 12192
rect 19116 12180 19122 12232
rect 21376 12220 21404 12260
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 19260 12192 21404 12220
rect 14384 12124 15056 12152
rect 8680 12056 10180 12084
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11330 12084 11336 12096
rect 11112 12056 11336 12084
rect 11112 12044 11118 12056
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 12713 12087 12771 12093
rect 12713 12053 12725 12087
rect 12759 12084 12771 12087
rect 12894 12084 12900 12096
rect 12759 12056 12900 12084
rect 12759 12053 12771 12056
rect 12713 12047 12771 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 14240 12056 14381 12084
rect 14240 12044 14246 12056
rect 14369 12053 14381 12056
rect 14415 12053 14427 12087
rect 14369 12047 14427 12053
rect 14461 12087 14519 12093
rect 14461 12053 14473 12087
rect 14507 12084 14519 12087
rect 14550 12084 14556 12096
rect 14507 12056 14556 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 15028 12093 15056 12124
rect 16482 12112 16488 12164
rect 16540 12152 16546 12164
rect 17313 12155 17371 12161
rect 17313 12152 17325 12155
rect 16540 12124 17325 12152
rect 16540 12112 16546 12124
rect 17313 12121 17325 12124
rect 17359 12152 17371 12155
rect 18064 12152 18092 12180
rect 18969 12155 19027 12161
rect 18969 12152 18981 12155
rect 17359 12124 18981 12152
rect 17359 12121 17371 12124
rect 17313 12115 17371 12121
rect 18969 12121 18981 12124
rect 19015 12121 19027 12155
rect 19260 12152 19288 12192
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 21726 12220 21732 12232
rect 21508 12192 21732 12220
rect 21508 12180 21514 12192
rect 21726 12180 21732 12192
rect 21784 12180 21790 12232
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22278 12220 22284 12232
rect 22143 12192 22284 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 22373 12223 22431 12229
rect 22373 12189 22385 12223
rect 22419 12220 22431 12223
rect 22738 12220 22744 12232
rect 22419 12192 22744 12220
rect 22419 12189 22431 12192
rect 22373 12183 22431 12189
rect 18969 12115 19027 12121
rect 19076 12124 19288 12152
rect 15013 12087 15071 12093
rect 15013 12053 15025 12087
rect 15059 12053 15071 12087
rect 15013 12047 15071 12053
rect 16666 12044 16672 12096
rect 16724 12084 16730 12096
rect 17402 12084 17408 12096
rect 16724 12056 17408 12084
rect 16724 12044 16730 12056
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 17523 12087 17581 12093
rect 17523 12053 17535 12087
rect 17569 12084 17581 12087
rect 18322 12084 18328 12096
rect 17569 12056 18328 12084
rect 17569 12053 17581 12056
rect 17523 12047 17581 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 18598 12044 18604 12096
rect 18656 12084 18662 12096
rect 18769 12087 18827 12093
rect 18769 12084 18781 12087
rect 18656 12056 18781 12084
rect 18656 12044 18662 12056
rect 18769 12053 18781 12056
rect 18815 12084 18827 12087
rect 19076 12084 19104 12124
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 22388 12152 22416 12183
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 22925 12223 22983 12229
rect 22925 12189 22937 12223
rect 22971 12220 22983 12223
rect 23566 12220 23572 12232
rect 22971 12192 23572 12220
rect 22971 12189 22983 12192
rect 22925 12183 22983 12189
rect 23566 12180 23572 12192
rect 23624 12180 23630 12232
rect 23891 12189 23949 12195
rect 23891 12186 23903 12189
rect 19760 12124 22416 12152
rect 23661 12155 23719 12161
rect 19760 12112 19766 12124
rect 23661 12121 23673 12155
rect 23707 12121 23719 12155
rect 23876 12155 23903 12186
rect 23937 12164 23949 12189
rect 24302 12180 24308 12232
rect 24360 12220 24366 12232
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 24360 12192 24409 12220
rect 24360 12180 24366 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 24946 12180 24952 12232
rect 25004 12180 25010 12232
rect 25038 12180 25044 12232
rect 25096 12180 25102 12232
rect 25424 12229 25452 12328
rect 26602 12316 26608 12368
rect 26660 12356 26666 12368
rect 27522 12356 27528 12368
rect 26660 12328 27528 12356
rect 26660 12316 26666 12328
rect 27522 12316 27528 12328
rect 27580 12316 27586 12368
rect 25682 12248 25688 12300
rect 25740 12288 25746 12300
rect 26973 12291 27031 12297
rect 26973 12288 26985 12291
rect 25740 12260 26985 12288
rect 25740 12248 25746 12260
rect 26973 12257 26985 12260
rect 27019 12257 27031 12291
rect 26973 12251 27031 12257
rect 27062 12248 27068 12300
rect 27120 12248 27126 12300
rect 28092 12288 28120 12384
rect 29178 12316 29184 12368
rect 29236 12356 29242 12368
rect 29730 12356 29736 12368
rect 29236 12328 29736 12356
rect 29236 12316 29242 12328
rect 29730 12316 29736 12328
rect 29788 12316 29794 12368
rect 27540 12260 28120 12288
rect 29549 12291 29607 12297
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12220 25467 12223
rect 25866 12220 25872 12232
rect 25455 12192 25872 12220
rect 25455 12189 25467 12192
rect 25409 12183 25467 12189
rect 23937 12155 23940 12164
rect 23876 12124 23940 12155
rect 23661 12115 23719 12121
rect 18815 12056 19104 12084
rect 18815 12053 18827 12056
rect 18769 12047 18827 12053
rect 20806 12044 20812 12096
rect 20864 12084 20870 12096
rect 21082 12084 21088 12096
rect 20864 12056 21088 12084
rect 20864 12044 20870 12056
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 21174 12044 21180 12096
rect 21232 12084 21238 12096
rect 21913 12087 21971 12093
rect 21913 12084 21925 12087
rect 21232 12056 21925 12084
rect 21232 12044 21238 12056
rect 21913 12053 21925 12056
rect 21959 12053 21971 12087
rect 21913 12047 21971 12053
rect 22278 12044 22284 12096
rect 22336 12044 22342 12096
rect 22462 12044 22468 12096
rect 22520 12084 22526 12096
rect 23014 12084 23020 12096
rect 22520 12056 23020 12084
rect 22520 12044 22526 12056
rect 23014 12044 23020 12056
rect 23072 12044 23078 12096
rect 23109 12087 23167 12093
rect 23109 12053 23121 12087
rect 23155 12084 23167 12087
rect 23198 12084 23204 12096
rect 23155 12056 23204 12084
rect 23155 12053 23167 12056
rect 23109 12047 23167 12053
rect 23198 12044 23204 12056
rect 23256 12084 23262 12096
rect 23676 12084 23704 12115
rect 23934 12112 23940 12124
rect 23992 12112 23998 12164
rect 24854 12112 24860 12164
rect 24912 12152 24918 12164
rect 25240 12152 25268 12183
rect 25866 12180 25872 12192
rect 25924 12180 25930 12232
rect 26789 12223 26847 12229
rect 26789 12189 26801 12223
rect 26835 12220 26847 12223
rect 26878 12220 26884 12232
rect 26835 12192 26884 12220
rect 26835 12189 26847 12192
rect 26789 12183 26847 12189
rect 26878 12180 26884 12192
rect 26936 12180 26942 12232
rect 27080 12220 27108 12248
rect 27540 12229 27568 12260
rect 29549 12257 29561 12291
rect 29595 12288 29607 12291
rect 29638 12288 29644 12300
rect 29595 12260 29644 12288
rect 29595 12257 29607 12260
rect 29549 12251 29607 12257
rect 29638 12248 29644 12260
rect 29696 12248 29702 12300
rect 27157 12223 27215 12229
rect 27157 12220 27169 12223
rect 27080 12192 27169 12220
rect 27157 12189 27169 12192
rect 27203 12189 27215 12223
rect 27157 12183 27215 12189
rect 27525 12223 27583 12229
rect 27525 12189 27537 12223
rect 27571 12189 27583 12223
rect 27525 12183 27583 12189
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 27801 12223 27859 12229
rect 27801 12220 27813 12223
rect 27672 12192 27813 12220
rect 27672 12180 27678 12192
rect 27801 12189 27813 12192
rect 27847 12189 27859 12223
rect 27801 12183 27859 12189
rect 27893 12223 27951 12229
rect 27893 12189 27905 12223
rect 27939 12189 27951 12223
rect 27893 12183 27951 12189
rect 24912 12124 25268 12152
rect 24912 12112 24918 12124
rect 25590 12112 25596 12164
rect 25648 12112 25654 12164
rect 25958 12112 25964 12164
rect 26016 12152 26022 12164
rect 27908 12152 27936 12183
rect 27982 12180 27988 12232
rect 28040 12220 28046 12232
rect 28166 12220 28172 12232
rect 28040 12192 28172 12220
rect 28040 12180 28046 12192
rect 28166 12180 28172 12192
rect 28224 12220 28230 12232
rect 28261 12223 28319 12229
rect 28261 12220 28273 12223
rect 28224 12192 28273 12220
rect 28224 12180 28230 12192
rect 28261 12189 28273 12192
rect 28307 12189 28319 12223
rect 28261 12183 28319 12189
rect 28445 12223 28503 12229
rect 28445 12189 28457 12223
rect 28491 12220 28503 12223
rect 29178 12220 29184 12232
rect 28491 12192 29184 12220
rect 28491 12189 28503 12192
rect 28445 12183 28503 12189
rect 26016 12124 27936 12152
rect 26016 12112 26022 12124
rect 24394 12084 24400 12096
rect 23256 12056 24400 12084
rect 23256 12044 23262 12056
rect 24394 12044 24400 12056
rect 24452 12084 24458 12096
rect 24581 12087 24639 12093
rect 24581 12084 24593 12087
rect 24452 12056 24593 12084
rect 24452 12044 24458 12056
rect 24581 12053 24593 12056
rect 24627 12053 24639 12087
rect 24581 12047 24639 12053
rect 25314 12044 25320 12096
rect 25372 12084 25378 12096
rect 28460 12084 28488 12183
rect 29178 12180 29184 12192
rect 29236 12180 29242 12232
rect 29932 12229 29960 12396
rect 30190 12384 30196 12436
rect 30248 12384 30254 12436
rect 31205 12427 31263 12433
rect 30760 12396 31064 12424
rect 29917 12223 29975 12229
rect 29917 12189 29929 12223
rect 29963 12189 29975 12223
rect 29917 12183 29975 12189
rect 30009 12223 30067 12229
rect 30009 12189 30021 12223
rect 30055 12220 30067 12223
rect 30466 12220 30472 12232
rect 30055 12192 30472 12220
rect 30055 12189 30067 12192
rect 30009 12183 30067 12189
rect 29086 12112 29092 12164
rect 29144 12152 29150 12164
rect 29454 12152 29460 12164
rect 29144 12124 29460 12152
rect 29144 12112 29150 12124
rect 29454 12112 29460 12124
rect 29512 12112 29518 12164
rect 29546 12112 29552 12164
rect 29604 12152 29610 12164
rect 29687 12155 29745 12161
rect 29687 12152 29699 12155
rect 29604 12124 29699 12152
rect 29604 12112 29610 12124
rect 29687 12121 29699 12124
rect 29733 12121 29745 12155
rect 29687 12115 29745 12121
rect 29822 12112 29828 12164
rect 29880 12112 29886 12164
rect 29932 12152 29960 12183
rect 30466 12180 30472 12192
rect 30524 12180 30530 12232
rect 30558 12180 30564 12232
rect 30616 12180 30622 12232
rect 30760 12229 30788 12396
rect 31036 12356 31064 12396
rect 31205 12393 31217 12427
rect 31251 12424 31263 12427
rect 31662 12424 31668 12436
rect 31251 12396 31668 12424
rect 31251 12393 31263 12396
rect 31205 12387 31263 12393
rect 31662 12384 31668 12396
rect 31720 12384 31726 12436
rect 32769 12427 32827 12433
rect 32769 12393 32781 12427
rect 32815 12424 32827 12427
rect 33502 12424 33508 12436
rect 32815 12396 33508 12424
rect 32815 12393 32827 12396
rect 32769 12387 32827 12393
rect 33502 12384 33508 12396
rect 33560 12384 33566 12436
rect 34517 12427 34575 12433
rect 34517 12393 34529 12427
rect 34563 12424 34575 12427
rect 34698 12424 34704 12436
rect 34563 12396 34704 12424
rect 34563 12393 34575 12396
rect 34517 12387 34575 12393
rect 34698 12384 34704 12396
rect 34756 12384 34762 12436
rect 34790 12384 34796 12436
rect 34848 12424 34854 12436
rect 35345 12427 35403 12433
rect 35345 12424 35357 12427
rect 34848 12396 35357 12424
rect 34848 12384 34854 12396
rect 35345 12393 35357 12396
rect 35391 12393 35403 12427
rect 35345 12387 35403 12393
rect 31036 12328 31984 12356
rect 30709 12223 30788 12229
rect 30709 12189 30721 12223
rect 30755 12192 30788 12223
rect 30755 12189 30767 12192
rect 30834 12190 30840 12242
rect 30892 12220 30898 12242
rect 30929 12223 30987 12229
rect 30929 12220 30941 12223
rect 30892 12192 30941 12220
rect 30892 12190 30898 12192
rect 30709 12183 30767 12189
rect 30929 12189 30941 12192
rect 30975 12189 30987 12223
rect 30929 12183 30987 12189
rect 31018 12180 31024 12232
rect 31076 12229 31082 12232
rect 31076 12220 31084 12229
rect 31076 12192 31121 12220
rect 31076 12183 31084 12192
rect 31076 12180 31082 12183
rect 30484 12152 30512 12180
rect 31956 12164 31984 12328
rect 34054 12316 34060 12368
rect 34112 12356 34118 12368
rect 34112 12328 35204 12356
rect 34112 12316 34118 12328
rect 32306 12248 32312 12300
rect 32364 12288 32370 12300
rect 32858 12288 32864 12300
rect 32364 12260 32864 12288
rect 32364 12248 32370 12260
rect 32122 12180 32128 12232
rect 32180 12220 32186 12232
rect 32600 12229 32628 12260
rect 32858 12248 32864 12260
rect 32916 12248 32922 12300
rect 33686 12248 33692 12300
rect 33744 12288 33750 12300
rect 34146 12288 34152 12300
rect 33744 12260 34152 12288
rect 33744 12248 33750 12260
rect 34146 12248 34152 12260
rect 34204 12248 34210 12300
rect 32401 12223 32459 12229
rect 32401 12220 32413 12223
rect 32180 12192 32413 12220
rect 32180 12180 32186 12192
rect 32401 12189 32413 12192
rect 32447 12189 32459 12223
rect 32401 12183 32459 12189
rect 32585 12223 32643 12229
rect 32585 12189 32597 12223
rect 32631 12189 32643 12223
rect 32585 12183 32643 12189
rect 33042 12180 33048 12232
rect 33100 12220 33106 12232
rect 33965 12223 34023 12229
rect 33965 12220 33977 12223
rect 33100 12192 33977 12220
rect 33100 12180 33106 12192
rect 33965 12189 33977 12192
rect 34011 12189 34023 12223
rect 34164 12220 34192 12248
rect 34241 12223 34299 12229
rect 34241 12220 34253 12223
rect 34164 12192 34253 12220
rect 33965 12183 34023 12189
rect 34241 12189 34253 12192
rect 34287 12189 34299 12223
rect 34241 12183 34299 12189
rect 34330 12180 34336 12232
rect 34388 12220 34394 12232
rect 34701 12223 34759 12229
rect 34701 12220 34713 12223
rect 34388 12192 34713 12220
rect 34388 12180 34394 12192
rect 34701 12189 34713 12192
rect 34747 12189 34759 12223
rect 34701 12183 34759 12189
rect 34790 12180 34796 12232
rect 34848 12229 34854 12232
rect 35176 12229 35204 12328
rect 34848 12223 34897 12229
rect 34848 12189 34851 12223
rect 34885 12189 34897 12223
rect 34848 12183 34897 12189
rect 35161 12223 35219 12229
rect 35161 12189 35173 12223
rect 35207 12189 35219 12223
rect 35161 12183 35219 12189
rect 34848 12180 34854 12183
rect 30837 12155 30895 12161
rect 30837 12152 30849 12155
rect 29932 12124 30420 12152
rect 30484 12124 30849 12152
rect 25372 12056 28488 12084
rect 30392 12084 30420 12124
rect 30837 12121 30849 12124
rect 30883 12121 30895 12155
rect 30837 12115 30895 12121
rect 30944 12124 31600 12152
rect 30944 12084 30972 12124
rect 30392 12056 30972 12084
rect 25372 12044 25378 12056
rect 31202 12044 31208 12096
rect 31260 12084 31266 12096
rect 31478 12084 31484 12096
rect 31260 12056 31484 12084
rect 31260 12044 31266 12056
rect 31478 12044 31484 12056
rect 31536 12044 31542 12096
rect 31572 12084 31600 12124
rect 31938 12112 31944 12164
rect 31996 12152 32002 12164
rect 33060 12152 33088 12180
rect 31996 12124 33088 12152
rect 31996 12112 32002 12124
rect 34054 12112 34060 12164
rect 34112 12152 34118 12164
rect 34149 12155 34207 12161
rect 34149 12152 34161 12155
rect 34112 12124 34161 12152
rect 34112 12112 34118 12124
rect 34149 12121 34161 12124
rect 34195 12121 34207 12155
rect 34149 12115 34207 12121
rect 34974 12112 34980 12164
rect 35032 12112 35038 12164
rect 35069 12155 35127 12161
rect 35069 12121 35081 12155
rect 35115 12121 35127 12155
rect 35069 12115 35127 12121
rect 35084 12084 35112 12115
rect 31572 12056 35112 12084
rect 1104 11994 36432 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 36432 11994
rect 1104 11920 36432 11942
rect 2406 11840 2412 11892
rect 2464 11840 2470 11892
rect 2961 11883 3019 11889
rect 2961 11849 2973 11883
rect 3007 11880 3019 11883
rect 3142 11880 3148 11892
rect 3007 11852 3148 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 3326 11840 3332 11892
rect 3384 11880 3390 11892
rect 4154 11880 4160 11892
rect 3384 11852 4160 11880
rect 3384 11840 3390 11852
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 4614 11880 4620 11892
rect 4479 11852 4620 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 5902 11840 5908 11892
rect 5960 11840 5966 11892
rect 5994 11840 6000 11892
rect 6052 11840 6058 11892
rect 6457 11883 6515 11889
rect 6457 11849 6469 11883
rect 6503 11880 6515 11883
rect 6546 11880 6552 11892
rect 6503 11852 6552 11880
rect 6503 11849 6515 11852
rect 6457 11843 6515 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 6730 11840 6736 11892
rect 6788 11840 6794 11892
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 7524 11852 7696 11880
rect 7524 11840 7530 11852
rect 6270 11812 6276 11824
rect 3068 11784 6276 11812
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 2623 11747 2681 11753
rect 2623 11744 2635 11747
rect 2556 11716 2635 11744
rect 2556 11704 2562 11716
rect 2623 11713 2635 11716
rect 2669 11713 2681 11747
rect 2623 11707 2681 11713
rect 2774 11704 2780 11756
rect 2832 11704 2838 11756
rect 3068 11753 3096 11784
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 6748 11812 6776 11840
rect 7282 11812 7288 11824
rect 6748 11784 7288 11812
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 4571 11716 4844 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 2884 11676 2912 11707
rect 2884 11648 3096 11676
rect 3068 11620 3096 11648
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 4338 11676 4344 11688
rect 3660 11648 4344 11676
rect 3660 11636 3666 11648
rect 4338 11636 4344 11648
rect 4396 11676 4402 11688
rect 4816 11685 4844 11716
rect 4890 11704 4896 11756
rect 4948 11704 4954 11756
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 4709 11679 4767 11685
rect 4709 11676 4721 11679
rect 4396 11648 4721 11676
rect 4396 11636 4402 11648
rect 4709 11645 4721 11648
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 5000 11676 5028 11707
rect 5258 11704 5264 11756
rect 5316 11704 5322 11756
rect 5442 11704 5448 11756
rect 5500 11704 5506 11756
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11744 5595 11747
rect 5626 11744 5632 11756
rect 5583 11716 5632 11744
rect 5583 11713 5595 11716
rect 5537 11707 5595 11713
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 5997 11747 6055 11753
rect 5997 11744 6009 11747
rect 5868 11716 6009 11744
rect 5868 11704 5874 11716
rect 5997 11713 6009 11716
rect 6043 11713 6055 11747
rect 5997 11707 6055 11713
rect 6178 11704 6184 11756
rect 6236 11704 6242 11756
rect 6638 11753 6644 11756
rect 6636 11744 6644 11753
rect 6599 11716 6644 11744
rect 6636 11707 6644 11716
rect 6638 11704 6644 11707
rect 6696 11704 6702 11756
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 6822 11704 6828 11756
rect 6880 11704 6886 11756
rect 7116 11753 7144 11784
rect 7282 11772 7288 11784
rect 7340 11772 7346 11824
rect 6953 11747 7011 11753
rect 6953 11744 6965 11747
rect 6932 11713 6965 11744
rect 6999 11713 7011 11747
rect 6932 11707 7011 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 5902 11676 5908 11688
rect 5000 11648 5488 11676
rect 4801 11639 4859 11645
rect 3050 11568 3056 11620
rect 3108 11608 3114 11620
rect 3510 11608 3516 11620
rect 3108 11580 3516 11608
rect 3108 11568 3114 11580
rect 3510 11568 3516 11580
rect 3568 11568 3574 11620
rect 4816 11608 4844 11639
rect 5460 11608 5488 11648
rect 5644 11648 5908 11676
rect 5644 11608 5672 11648
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 6932 11676 6960 11707
rect 7190 11704 7196 11756
rect 7248 11704 7254 11756
rect 7374 11704 7380 11756
rect 7432 11744 7438 11756
rect 7668 11753 7696 11852
rect 8662 11840 8668 11892
rect 8720 11840 8726 11892
rect 9125 11883 9183 11889
rect 9125 11849 9137 11883
rect 9171 11880 9183 11883
rect 9398 11880 9404 11892
rect 9171 11852 9404 11880
rect 9171 11849 9183 11852
rect 9125 11843 9183 11849
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9548 11852 9873 11880
rect 9548 11840 9554 11852
rect 9861 11849 9873 11852
rect 9907 11880 9919 11883
rect 9950 11880 9956 11892
rect 9907 11852 9956 11880
rect 9907 11849 9919 11852
rect 9861 11843 9919 11849
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10042 11840 10048 11892
rect 10100 11840 10106 11892
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10686 11880 10692 11892
rect 10376 11852 10692 11880
rect 10376 11840 10382 11852
rect 10686 11840 10692 11852
rect 10744 11880 10750 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10744 11852 10977 11880
rect 10744 11840 10750 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 10965 11843 11023 11849
rect 11072 11852 15608 11880
rect 8110 11812 8116 11824
rect 7760 11784 8116 11812
rect 7760 11753 7788 11784
rect 8110 11772 8116 11784
rect 8168 11812 8174 11824
rect 8680 11812 8708 11840
rect 11072 11812 11100 11852
rect 8168 11784 8708 11812
rect 9692 11784 11100 11812
rect 8168 11772 8174 11784
rect 7469 11747 7527 11753
rect 7469 11744 7481 11747
rect 7432 11716 7481 11744
rect 7432 11704 7438 11716
rect 7469 11713 7481 11716
rect 7515 11713 7527 11747
rect 7469 11707 7527 11713
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 7668 11676 7696 11707
rect 6144 11648 7696 11676
rect 7944 11676 7972 11707
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11744 8539 11747
rect 8588 11744 8616 11784
rect 8527 11716 8616 11744
rect 8665 11747 8723 11753
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 8665 11713 8677 11747
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 8570 11676 8576 11688
rect 7944 11648 8576 11676
rect 6144 11636 6150 11648
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 8680 11676 8708 11707
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 8911 11747 8969 11753
rect 8911 11713 8923 11747
rect 8957 11744 8969 11747
rect 9582 11744 9588 11756
rect 8957 11716 9588 11744
rect 8957 11713 8969 11716
rect 8911 11707 8969 11713
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 9692 11753 9720 11784
rect 10244 11753 10272 11784
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 12032 11784 12434 11812
rect 12032 11772 12038 11784
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 9956 11747 10014 11753
rect 9956 11713 9968 11747
rect 10002 11713 10014 11747
rect 9956 11707 10014 11713
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 9217 11679 9275 11685
rect 9217 11676 9229 11679
rect 8680 11648 9229 11676
rect 9217 11645 9229 11648
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 9968 11676 9996 11707
rect 10594 11704 10600 11756
rect 10652 11744 10658 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 10652 11716 10701 11744
rect 10652 11704 10658 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11296 11716 11713 11744
rect 11296 11704 11302 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11713 12311 11747
rect 12406 11744 12434 11784
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 15470 11812 15476 11824
rect 14240 11784 15476 11812
rect 14240 11772 14246 11784
rect 15470 11772 15476 11784
rect 15528 11772 15534 11824
rect 15580 11812 15608 11852
rect 16666 11840 16672 11892
rect 16724 11840 16730 11892
rect 16758 11840 16764 11892
rect 16816 11840 16822 11892
rect 19702 11880 19708 11892
rect 17604 11852 19708 11880
rect 16776 11812 16804 11840
rect 17405 11815 17463 11821
rect 17405 11812 17417 11815
rect 15580 11784 16804 11812
rect 16960 11784 17417 11812
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12406 11716 13001 11744
rect 12253 11707 12311 11713
rect 12989 11713 13001 11716
rect 13035 11744 13047 11747
rect 13170 11744 13176 11756
rect 13035 11716 13176 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 9364 11648 9996 11676
rect 10413 11679 10471 11685
rect 9364 11636 9370 11648
rect 10413 11645 10425 11679
rect 10459 11676 10471 11679
rect 10502 11676 10508 11688
rect 10459 11648 10508 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 11514 11636 11520 11688
rect 11572 11636 11578 11688
rect 4816 11580 5304 11608
rect 5460 11580 5672 11608
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 4948 11512 5181 11540
rect 4948 11500 4954 11512
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 5276 11540 5304 11580
rect 5718 11568 5724 11620
rect 5776 11608 5782 11620
rect 7193 11611 7251 11617
rect 7193 11608 7205 11611
rect 5776 11580 7205 11608
rect 5776 11568 5782 11580
rect 7193 11577 7205 11580
rect 7239 11577 7251 11611
rect 7193 11571 7251 11577
rect 7374 11568 7380 11620
rect 7432 11608 7438 11620
rect 7469 11611 7527 11617
rect 7469 11608 7481 11611
rect 7432 11580 7481 11608
rect 7432 11568 7438 11580
rect 7469 11577 7481 11580
rect 7515 11577 7527 11611
rect 7469 11571 7527 11577
rect 7745 11611 7803 11617
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 8846 11608 8852 11620
rect 7791 11580 8852 11608
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 8846 11568 8852 11580
rect 8904 11568 8910 11620
rect 9585 11611 9643 11617
rect 9585 11577 9597 11611
rect 9631 11608 9643 11611
rect 12268 11608 12296 11707
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 13446 11744 13452 11756
rect 13311 11716 13452 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13446 11704 13452 11716
rect 13504 11744 13510 11756
rect 14550 11744 14556 11756
rect 13504 11716 14556 11744
rect 13504 11704 13510 11716
rect 14550 11704 14556 11716
rect 14608 11704 14614 11756
rect 15194 11704 15200 11756
rect 15252 11744 15258 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 15252 11716 15393 11744
rect 15252 11704 15258 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 15746 11744 15752 11756
rect 15611 11716 15752 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12492 11648 12541 11676
rect 12492 11636 12498 11648
rect 12529 11645 12541 11648
rect 12575 11676 12587 11679
rect 12802 11676 12808 11688
rect 12575 11648 12808 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 12802 11636 12808 11648
rect 12860 11676 12866 11688
rect 13354 11676 13360 11688
rect 12860 11648 13360 11676
rect 12860 11636 12866 11648
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 15396 11676 15424 11707
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 16850 11747 16856 11756
rect 16776 11744 16856 11747
rect 15856 11719 16856 11744
rect 15856 11716 16804 11719
rect 15856 11676 15884 11716
rect 16850 11704 16856 11719
rect 16908 11704 16914 11756
rect 15396 11648 15884 11676
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 16960 11676 16988 11784
rect 17405 11781 17417 11784
rect 17451 11781 17463 11815
rect 17405 11775 17463 11781
rect 17604 11756 17632 11852
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 19886 11840 19892 11892
rect 19944 11880 19950 11892
rect 20530 11880 20536 11892
rect 19944 11852 20536 11880
rect 19944 11840 19950 11852
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 23014 11840 23020 11892
rect 23072 11880 23078 11892
rect 23109 11883 23167 11889
rect 23109 11880 23121 11883
rect 23072 11852 23121 11880
rect 23072 11840 23078 11852
rect 23109 11849 23121 11852
rect 23155 11880 23167 11883
rect 23474 11880 23480 11892
rect 23155 11852 23480 11880
rect 23155 11849 23167 11852
rect 23109 11843 23167 11849
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 26694 11840 26700 11892
rect 26752 11840 26758 11892
rect 27522 11840 27528 11892
rect 27580 11880 27586 11892
rect 27580 11852 27844 11880
rect 27580 11840 27586 11852
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 20220 11784 20668 11812
rect 20220 11772 20226 11784
rect 17218 11704 17224 11756
rect 17276 11744 17282 11756
rect 17313 11747 17371 11753
rect 17313 11744 17325 11747
rect 17276 11716 17325 11744
rect 17276 11704 17282 11716
rect 17313 11713 17325 11716
rect 17359 11713 17371 11747
rect 17313 11707 17371 11713
rect 17586 11704 17592 11756
rect 17644 11704 17650 11756
rect 17678 11704 17684 11756
rect 17736 11704 17742 11756
rect 17862 11704 17868 11756
rect 17920 11704 17926 11756
rect 17954 11704 17960 11756
rect 18012 11704 18018 11756
rect 19150 11704 19156 11756
rect 19208 11744 19214 11756
rect 19886 11744 19892 11756
rect 19208 11716 19892 11744
rect 19208 11704 19214 11716
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 20254 11704 20260 11756
rect 20312 11744 20318 11756
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 20312 11716 20361 11744
rect 20312 11704 20318 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 20530 11704 20536 11756
rect 20588 11704 20594 11756
rect 20640 11753 20668 11784
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 23198 11812 23204 11824
rect 22336 11784 23204 11812
rect 22336 11772 22342 11784
rect 23198 11772 23204 11784
rect 23256 11772 23262 11824
rect 25038 11772 25044 11824
rect 25096 11812 25102 11824
rect 25096 11784 27752 11812
rect 25096 11772 25102 11784
rect 27724 11756 27752 11784
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11713 20683 11747
rect 20625 11707 20683 11713
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 21542 11744 21548 11756
rect 20763 11716 21548 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 23293 11747 23351 11753
rect 23293 11713 23305 11747
rect 23339 11713 23351 11747
rect 23293 11707 23351 11713
rect 16816 11648 16988 11676
rect 17037 11679 17095 11685
rect 16816 11636 16822 11648
rect 17037 11645 17049 11679
rect 17083 11676 17095 11679
rect 17494 11676 17500 11688
rect 17083 11648 17500 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 23308 11676 23336 11707
rect 24026 11704 24032 11756
rect 24084 11744 24090 11756
rect 26605 11747 26663 11753
rect 26605 11744 26617 11747
rect 24084 11716 26617 11744
rect 24084 11704 24090 11716
rect 26605 11713 26617 11716
rect 26651 11744 26663 11747
rect 26694 11744 26700 11756
rect 26651 11716 26700 11744
rect 26651 11713 26663 11716
rect 26605 11707 26663 11713
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 26789 11747 26847 11753
rect 26789 11713 26801 11747
rect 26835 11744 26847 11747
rect 27154 11744 27160 11756
rect 26835 11716 27160 11744
rect 26835 11713 26847 11716
rect 26789 11707 26847 11713
rect 27154 11704 27160 11716
rect 27212 11704 27218 11756
rect 27246 11704 27252 11756
rect 27304 11704 27310 11756
rect 27433 11747 27491 11753
rect 27433 11713 27445 11747
rect 27479 11744 27491 11747
rect 27614 11744 27620 11756
rect 27479 11716 27620 11744
rect 27479 11713 27491 11716
rect 27433 11707 27491 11713
rect 27614 11704 27620 11716
rect 27672 11704 27678 11756
rect 27706 11704 27712 11756
rect 27764 11704 27770 11756
rect 27816 11744 27844 11852
rect 30558 11840 30564 11892
rect 30616 11880 30622 11892
rect 30745 11883 30803 11889
rect 30745 11880 30757 11883
rect 30616 11852 30757 11880
rect 30616 11840 30622 11852
rect 30745 11849 30757 11852
rect 30791 11849 30803 11883
rect 30745 11843 30803 11849
rect 31018 11840 31024 11892
rect 31076 11840 31082 11892
rect 31481 11883 31539 11889
rect 31481 11849 31493 11883
rect 31527 11880 31539 11883
rect 31754 11880 31760 11892
rect 31527 11852 31760 11880
rect 31527 11849 31539 11852
rect 31481 11843 31539 11849
rect 31754 11840 31760 11852
rect 31812 11840 31818 11892
rect 31849 11883 31907 11889
rect 31849 11849 31861 11883
rect 31895 11880 31907 11883
rect 32766 11880 32772 11892
rect 31895 11852 32772 11880
rect 31895 11849 31907 11852
rect 31849 11843 31907 11849
rect 28261 11815 28319 11821
rect 28261 11781 28273 11815
rect 28307 11812 28319 11815
rect 29362 11812 29368 11824
rect 28307 11784 29368 11812
rect 28307 11781 28319 11784
rect 28261 11775 28319 11781
rect 29362 11772 29368 11784
rect 29420 11772 29426 11824
rect 30469 11815 30527 11821
rect 30469 11781 30481 11815
rect 30515 11812 30527 11815
rect 30650 11812 30656 11824
rect 30515 11784 30656 11812
rect 30515 11781 30527 11784
rect 30469 11775 30527 11781
rect 30650 11772 30656 11784
rect 30708 11772 30714 11824
rect 31036 11812 31064 11840
rect 31864 11812 31892 11843
rect 32766 11840 32772 11852
rect 32824 11840 32830 11892
rect 32858 11840 32864 11892
rect 32916 11880 32922 11892
rect 34330 11880 34336 11892
rect 32916 11852 34336 11880
rect 32916 11840 32922 11852
rect 34330 11840 34336 11852
rect 34388 11840 34394 11892
rect 30944 11784 31064 11812
rect 31312 11784 31892 11812
rect 28994 11744 29000 11756
rect 27816 11716 29000 11744
rect 28994 11704 29000 11716
rect 29052 11704 29058 11756
rect 29181 11747 29239 11753
rect 29181 11713 29193 11747
rect 29227 11713 29239 11747
rect 29181 11707 29239 11713
rect 25314 11676 25320 11688
rect 23308 11648 25320 11676
rect 25314 11636 25320 11648
rect 25372 11636 25378 11688
rect 27341 11679 27399 11685
rect 27341 11645 27353 11679
rect 27387 11676 27399 11679
rect 29196 11676 29224 11707
rect 30098 11704 30104 11756
rect 30156 11704 30162 11756
rect 30282 11753 30288 11756
rect 30259 11747 30288 11753
rect 30259 11713 30271 11747
rect 30259 11707 30288 11713
rect 30282 11704 30288 11707
rect 30340 11704 30346 11756
rect 30374 11704 30380 11756
rect 30432 11704 30438 11756
rect 30561 11747 30619 11753
rect 30561 11713 30573 11747
rect 30607 11744 30619 11747
rect 30944 11744 30972 11784
rect 30607 11716 30972 11744
rect 30607 11713 30619 11716
rect 30561 11707 30619 11713
rect 31018 11704 31024 11756
rect 31076 11744 31082 11756
rect 31312 11753 31340 11784
rect 32950 11772 32956 11824
rect 33008 11772 33014 11824
rect 34514 11772 34520 11824
rect 34572 11812 34578 11824
rect 34572 11784 34638 11812
rect 34572 11772 34578 11784
rect 31297 11747 31355 11753
rect 31297 11744 31309 11747
rect 31076 11716 31309 11744
rect 31076 11704 31082 11716
rect 31297 11713 31309 11716
rect 31343 11713 31355 11747
rect 31297 11707 31355 11713
rect 31386 11704 31392 11756
rect 31444 11744 31450 11756
rect 31665 11747 31723 11753
rect 31665 11744 31677 11747
rect 31444 11716 31677 11744
rect 31444 11704 31450 11716
rect 31665 11713 31677 11716
rect 31711 11744 31723 11747
rect 32309 11747 32367 11753
rect 32309 11744 32321 11747
rect 31711 11716 32321 11744
rect 31711 11713 31723 11716
rect 31665 11707 31723 11713
rect 32309 11713 32321 11716
rect 32355 11713 32367 11747
rect 32309 11707 32367 11713
rect 32674 11704 32680 11756
rect 32732 11704 32738 11756
rect 32398 11676 32404 11688
rect 27387 11648 28212 11676
rect 29196 11648 32404 11676
rect 27387 11645 27399 11648
rect 27341 11639 27399 11645
rect 12713 11611 12771 11617
rect 12713 11608 12725 11611
rect 9631 11580 10640 11608
rect 12268 11580 12725 11608
rect 9631 11577 9643 11580
rect 9585 11571 9643 11577
rect 10612 11552 10640 11580
rect 12713 11577 12725 11580
rect 12759 11577 12771 11611
rect 12713 11571 12771 11577
rect 13630 11568 13636 11620
rect 13688 11608 13694 11620
rect 17862 11608 17868 11620
rect 13688 11580 17868 11608
rect 13688 11568 13694 11580
rect 17862 11568 17868 11580
rect 17920 11568 17926 11620
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18012 11580 21128 11608
rect 18012 11568 18018 11580
rect 5626 11540 5632 11552
rect 5276 11512 5632 11540
rect 5169 11503 5227 11509
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 8021 11543 8079 11549
rect 8021 11509 8033 11543
rect 8067 11540 8079 11543
rect 8938 11540 8944 11552
rect 8067 11512 8944 11540
rect 8067 11509 8079 11512
rect 8021 11503 8079 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9493 11543 9551 11549
rect 9493 11509 9505 11543
rect 9539 11540 9551 11543
rect 10502 11540 10508 11552
rect 9539 11512 10508 11540
rect 9539 11509 9551 11512
rect 9493 11503 9551 11509
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 10594 11500 10600 11552
rect 10652 11500 10658 11552
rect 12894 11500 12900 11552
rect 12952 11500 12958 11552
rect 15194 11500 15200 11552
rect 15252 11500 15258 11552
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 16853 11543 16911 11549
rect 16853 11540 16865 11543
rect 16816 11512 16865 11540
rect 16816 11500 16822 11512
rect 16853 11509 16865 11512
rect 16899 11509 16911 11543
rect 16853 11503 16911 11509
rect 18506 11500 18512 11552
rect 18564 11540 18570 11552
rect 19702 11540 19708 11552
rect 18564 11512 19708 11540
rect 18564 11500 18570 11512
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 20714 11500 20720 11552
rect 20772 11540 20778 11552
rect 20993 11543 21051 11549
rect 20993 11540 21005 11543
rect 20772 11512 21005 11540
rect 20772 11500 20778 11512
rect 20993 11509 21005 11512
rect 21039 11509 21051 11543
rect 21100 11540 21128 11580
rect 21450 11568 21456 11620
rect 21508 11608 21514 11620
rect 26973 11611 27031 11617
rect 26973 11608 26985 11611
rect 21508 11580 26985 11608
rect 21508 11568 21514 11580
rect 26973 11577 26985 11580
rect 27019 11577 27031 11611
rect 26973 11571 27031 11577
rect 27080 11580 27660 11608
rect 22646 11540 22652 11552
rect 21100 11512 22652 11540
rect 20993 11503 21051 11509
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 27080 11540 27108 11580
rect 25556 11512 27108 11540
rect 25556 11500 25562 11512
rect 27522 11500 27528 11552
rect 27580 11500 27586 11552
rect 27632 11540 27660 11580
rect 28074 11568 28080 11620
rect 28132 11568 28138 11620
rect 28184 11608 28212 11648
rect 32398 11636 32404 11648
rect 32456 11636 32462 11688
rect 35434 11636 35440 11688
rect 35492 11676 35498 11688
rect 35805 11679 35863 11685
rect 35805 11676 35817 11679
rect 35492 11648 35817 11676
rect 35492 11636 35498 11648
rect 35805 11645 35817 11648
rect 35851 11645 35863 11679
rect 35805 11639 35863 11645
rect 36078 11636 36084 11688
rect 36136 11636 36142 11688
rect 29454 11608 29460 11620
rect 28184 11580 29460 11608
rect 29454 11568 29460 11580
rect 29512 11568 29518 11620
rect 29546 11568 29552 11620
rect 29604 11608 29610 11620
rect 34698 11608 34704 11620
rect 29604 11580 34704 11608
rect 29604 11568 29610 11580
rect 34698 11568 34704 11580
rect 34756 11568 34762 11620
rect 28905 11543 28963 11549
rect 28905 11540 28917 11543
rect 27632 11512 28917 11540
rect 28905 11509 28917 11512
rect 28951 11540 28963 11543
rect 28994 11540 29000 11552
rect 28951 11512 29000 11540
rect 28951 11509 28963 11512
rect 28905 11503 28963 11509
rect 28994 11500 29000 11512
rect 29052 11500 29058 11552
rect 33042 11500 33048 11552
rect 33100 11500 33106 11552
rect 34333 11543 34391 11549
rect 34333 11509 34345 11543
rect 34379 11540 34391 11543
rect 34790 11540 34796 11552
rect 34379 11512 34796 11540
rect 34379 11509 34391 11512
rect 34333 11503 34391 11509
rect 34790 11500 34796 11512
rect 34848 11500 34854 11552
rect 1104 11450 36432 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 36432 11450
rect 1104 11376 36432 11398
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2866 11336 2872 11348
rect 2363 11308 2872 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11305 3111 11339
rect 6454 11336 6460 11348
rect 3053 11299 3111 11305
rect 3896 11308 6460 11336
rect 2406 11228 2412 11280
rect 2464 11268 2470 11280
rect 3068 11268 3096 11299
rect 2464 11240 3096 11268
rect 2464 11228 2470 11240
rect 3326 11228 3332 11280
rect 3384 11228 3390 11280
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11169 2099 11203
rect 3344 11200 3372 11228
rect 3789 11203 3847 11209
rect 3789 11200 3801 11203
rect 2041 11163 2099 11169
rect 2884 11172 3801 11200
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 2056 11132 2084 11163
rect 2884 11144 2912 11172
rect 3789 11169 3801 11172
rect 3835 11169 3847 11203
rect 3789 11163 3847 11169
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2056 11104 2421 11132
rect 1949 11095 2007 11101
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 1964 11064 1992 11095
rect 2590 11092 2596 11144
rect 2648 11092 2654 11144
rect 2682 11092 2688 11144
rect 2740 11092 2746 11144
rect 2866 11092 2872 11144
rect 2924 11092 2930 11144
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3142 11132 3148 11144
rect 3099 11104 3148 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 1964 11036 2452 11064
rect 2424 10996 2452 11036
rect 2498 11024 2504 11076
rect 2556 11064 2562 11076
rect 2976 11064 3004 11095
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3896 11132 3924 11308
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 10870 11336 10876 11348
rect 10152 11308 10876 11336
rect 4709 11271 4767 11277
rect 4709 11237 4721 11271
rect 4755 11268 4767 11271
rect 5258 11268 5264 11280
rect 4755 11240 5264 11268
rect 4755 11237 4767 11240
rect 4709 11231 4767 11237
rect 5258 11228 5264 11240
rect 5316 11228 5322 11280
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 5721 11271 5779 11277
rect 5721 11268 5733 11271
rect 5592 11240 5733 11268
rect 5592 11228 5598 11240
rect 5721 11237 5733 11240
rect 5767 11268 5779 11271
rect 8478 11268 8484 11280
rect 5767 11240 8484 11268
rect 5767 11237 5779 11240
rect 5721 11231 5779 11237
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 8662 11228 8668 11280
rect 8720 11268 8726 11280
rect 10152 11268 10180 11308
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 11793 11339 11851 11345
rect 11793 11336 11805 11339
rect 11204 11308 11805 11336
rect 11204 11296 11210 11308
rect 11793 11305 11805 11308
rect 11839 11305 11851 11339
rect 11793 11299 11851 11305
rect 12345 11339 12403 11345
rect 12345 11305 12357 11339
rect 12391 11336 12403 11339
rect 12434 11336 12440 11348
rect 12391 11308 12440 11336
rect 12391 11305 12403 11308
rect 12345 11299 12403 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 12526 11296 12532 11348
rect 12584 11296 12590 11348
rect 12894 11296 12900 11348
rect 12952 11296 12958 11348
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 16908 11308 17141 11336
rect 16908 11296 16914 11308
rect 17129 11305 17141 11308
rect 17175 11305 17187 11339
rect 19429 11339 19487 11345
rect 17129 11299 17187 11305
rect 17328 11308 19334 11336
rect 11698 11268 11704 11280
rect 8720 11240 10180 11268
rect 10612 11240 11704 11268
rect 8720 11228 8726 11240
rect 4798 11200 4804 11212
rect 4172 11172 4804 11200
rect 4172 11141 4200 11172
rect 4798 11160 4804 11172
rect 4856 11200 4862 11212
rect 5905 11203 5963 11209
rect 5905 11200 5917 11203
rect 4856 11172 5917 11200
rect 4856 11160 4862 11172
rect 5905 11169 5917 11172
rect 5951 11169 5963 11203
rect 6730 11200 6736 11212
rect 5905 11163 5963 11169
rect 6380 11172 6736 11200
rect 3283 11104 3924 11132
rect 3973 11135 4031 11141
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3973 11101 3985 11135
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 3252 11064 3280 11095
rect 2556 11036 3004 11064
rect 3068 11036 3280 11064
rect 3988 11064 4016 11095
rect 4246 11092 4252 11144
rect 4304 11092 4310 11144
rect 4890 11092 4896 11144
rect 4948 11092 4954 11144
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 5040 11104 5085 11132
rect 5040 11092 5046 11104
rect 5258 11092 5264 11144
rect 5316 11092 5322 11144
rect 5399 11135 5457 11141
rect 5399 11101 5411 11135
rect 5445 11132 5457 11135
rect 5718 11132 5724 11144
rect 5445 11104 5724 11132
rect 5445 11101 5457 11104
rect 5399 11095 5457 11101
rect 5718 11092 5724 11104
rect 5776 11092 5782 11144
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11132 5871 11135
rect 5859 11104 5948 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 4341 11067 4399 11073
rect 4341 11064 4353 11067
rect 3988 11036 4353 11064
rect 2556 11024 2562 11036
rect 3068 11008 3096 11036
rect 4172 11008 4200 11036
rect 4341 11033 4353 11036
rect 4387 11064 4399 11067
rect 5000 11064 5028 11092
rect 5920 11076 5948 11104
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 6380 11141 6408 11172
rect 6730 11160 6736 11172
rect 6788 11200 6794 11212
rect 7374 11200 7380 11212
rect 6788 11172 7380 11200
rect 6788 11160 6794 11172
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8628 11172 8953 11200
rect 8628 11160 8634 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9416 11172 10180 11200
rect 9312 11144 9364 11150
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11101 6423 11135
rect 6365 11095 6423 11101
rect 6454 11092 6460 11144
rect 6512 11092 6518 11144
rect 7006 11092 7012 11144
rect 7064 11132 7070 11144
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 7064 11104 7113 11132
rect 7064 11092 7070 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 7208 11104 7880 11132
rect 4387 11036 5028 11064
rect 5169 11067 5227 11073
rect 4387 11033 4399 11036
rect 4341 11027 4399 11033
rect 5169 11033 5181 11067
rect 5215 11064 5227 11067
rect 5626 11064 5632 11076
rect 5215 11036 5632 11064
rect 5215 11033 5227 11036
rect 5169 11027 5227 11033
rect 5460 11008 5488 11036
rect 5626 11024 5632 11036
rect 5684 11064 5690 11076
rect 5684 11036 5856 11064
rect 5684 11024 5690 11036
rect 3050 10996 3056 11008
rect 2424 10968 3056 10996
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 3421 10999 3479 11005
rect 3421 10965 3433 10999
rect 3467 10996 3479 10999
rect 3694 10996 3700 11008
rect 3467 10968 3700 10996
rect 3467 10965 3479 10968
rect 3421 10959 3479 10965
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 4154 10956 4160 11008
rect 4212 10956 4218 11008
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 4706 10996 4712 11008
rect 4304 10968 4712 10996
rect 4304 10956 4310 10968
rect 4706 10956 4712 10968
rect 4764 10996 4770 11008
rect 4801 10999 4859 11005
rect 4801 10996 4813 10999
rect 4764 10968 4813 10996
rect 4764 10956 4770 10968
rect 4801 10965 4813 10968
rect 4847 10965 4859 10999
rect 4801 10959 4859 10965
rect 5442 10956 5448 11008
rect 5500 10956 5506 11008
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 5828 10996 5856 11036
rect 5902 11024 5908 11076
rect 5960 11024 5966 11076
rect 6273 11067 6331 11073
rect 6273 11033 6285 11067
rect 6319 11064 6331 11067
rect 7024 11064 7052 11092
rect 7208 11064 7236 11104
rect 6319 11036 7052 11064
rect 7116 11036 7236 11064
rect 7653 11067 7711 11073
rect 6319 11033 6331 11036
rect 6273 11027 6331 11033
rect 6822 10996 6828 11008
rect 5828 10968 6828 10996
rect 6822 10956 6828 10968
rect 6880 10996 6886 11008
rect 7116 10996 7144 11036
rect 7653 11033 7665 11067
rect 7699 11064 7711 11067
rect 7742 11064 7748 11076
rect 7699 11036 7748 11064
rect 7699 11033 7711 11036
rect 7653 11027 7711 11033
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 7852 11064 7880 11104
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8481 11135 8539 11141
rect 8481 11132 8493 11135
rect 8352 11104 8493 11132
rect 8352 11092 8358 11104
rect 8481 11101 8493 11104
rect 8527 11132 8539 11135
rect 9122 11132 9128 11144
rect 8527 11104 9128 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9416 11142 9444 11172
rect 9364 11114 9444 11142
rect 9950 11092 9956 11144
rect 10008 11092 10014 11144
rect 10152 11141 10180 11172
rect 10612 11144 10640 11240
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 17218 11268 17224 11280
rect 12406 11240 17224 11268
rect 12406 11200 12434 11240
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 10888 11172 12434 11200
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 9312 11086 9364 11092
rect 8662 11064 8668 11076
rect 7852 11036 8668 11064
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 9968 11064 9996 11092
rect 10336 11064 10364 11095
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 10888 11141 10916 11172
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 13722 11200 13728 11212
rect 12584 11172 13728 11200
rect 12584 11160 12590 11172
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 15286 11200 15292 11212
rect 14844 11172 15292 11200
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 11974 11092 11980 11144
rect 12032 11092 12038 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12710 11132 12716 11144
rect 12207 11104 12716 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11132 12863 11135
rect 13081 11135 13139 11141
rect 12851 11104 13032 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 9968 11036 10364 11064
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 12437 11067 12495 11073
rect 10560 11036 12388 11064
rect 10560 11024 10566 11036
rect 6880 10968 7144 10996
rect 6880 10956 6886 10968
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 9214 10996 9220 11008
rect 8536 10968 9220 10996
rect 8536 10956 8542 10968
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 10226 10956 10232 11008
rect 10284 10956 10290 11008
rect 12360 10996 12388 11036
rect 12437 11033 12449 11067
rect 12483 11064 12495 11067
rect 13004 11064 13032 11104
rect 13081 11101 13093 11135
rect 13127 11132 13139 11135
rect 13446 11132 13452 11144
rect 13127 11104 13452 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14366 11132 14372 11144
rect 14056 11104 14372 11132
rect 14056 11092 14062 11104
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 14550 11092 14556 11144
rect 14608 11092 14614 11144
rect 14642 11092 14648 11144
rect 14700 11092 14706 11144
rect 14844 11141 14872 11172
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 16482 11160 16488 11212
rect 16540 11200 16546 11212
rect 16761 11203 16819 11209
rect 16761 11200 16773 11203
rect 16540 11172 16773 11200
rect 16540 11160 16546 11172
rect 16761 11169 16773 11172
rect 16807 11169 16819 11203
rect 17328 11200 17356 11308
rect 17678 11228 17684 11280
rect 17736 11268 17742 11280
rect 18138 11268 18144 11280
rect 17736 11240 18144 11268
rect 17736 11228 17742 11240
rect 18138 11228 18144 11240
rect 18196 11228 18202 11280
rect 19306 11268 19334 11308
rect 19429 11305 19441 11339
rect 19475 11305 19487 11339
rect 19429 11299 19487 11305
rect 19444 11268 19472 11299
rect 19610 11296 19616 11348
rect 19668 11296 19674 11348
rect 19702 11296 19708 11348
rect 19760 11336 19766 11348
rect 22094 11336 22100 11348
rect 19760 11308 22100 11336
rect 19760 11296 19766 11308
rect 22094 11296 22100 11308
rect 22152 11336 22158 11348
rect 23014 11336 23020 11348
rect 22152 11308 23020 11336
rect 22152 11296 22158 11308
rect 23014 11296 23020 11308
rect 23072 11296 23078 11348
rect 23201 11339 23259 11345
rect 23201 11305 23213 11339
rect 23247 11336 23259 11339
rect 23290 11336 23296 11348
rect 23247 11308 23296 11336
rect 23247 11305 23259 11308
rect 23201 11299 23259 11305
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 23474 11296 23480 11348
rect 23532 11296 23538 11348
rect 24302 11296 24308 11348
rect 24360 11336 24366 11348
rect 26602 11336 26608 11348
rect 24360 11308 26608 11336
rect 24360 11296 24366 11308
rect 26602 11296 26608 11308
rect 26660 11296 26666 11348
rect 26786 11296 26792 11348
rect 26844 11336 26850 11348
rect 27614 11336 27620 11348
rect 26844 11308 27620 11336
rect 26844 11296 26850 11308
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 29730 11336 29736 11348
rect 28000 11308 29736 11336
rect 19978 11268 19984 11280
rect 19306 11240 19380 11268
rect 19444 11240 19984 11268
rect 19352 11200 19380 11240
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 27246 11228 27252 11280
rect 27304 11268 27310 11280
rect 28000 11268 28028 11308
rect 29730 11296 29736 11308
rect 29788 11296 29794 11348
rect 31573 11339 31631 11345
rect 31573 11305 31585 11339
rect 31619 11336 31631 11339
rect 31754 11336 31760 11348
rect 31619 11308 31760 11336
rect 31619 11305 31631 11308
rect 31573 11299 31631 11305
rect 31754 11296 31760 11308
rect 31812 11296 31818 11348
rect 32582 11296 32588 11348
rect 32640 11296 32646 11348
rect 33042 11336 33048 11348
rect 32876 11308 33048 11336
rect 27304 11240 28028 11268
rect 27304 11228 27310 11240
rect 19610 11200 19616 11212
rect 16761 11163 16819 11169
rect 16960 11172 17356 11200
rect 17604 11172 19288 11200
rect 19352 11172 19616 11200
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11101 14887 11135
rect 14829 11095 14887 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11132 14979 11135
rect 16666 11132 16672 11144
rect 14967 11104 16672 11132
rect 14967 11101 14979 11104
rect 14921 11095 14979 11101
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 16960 11141 16988 11172
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11101 17003 11135
rect 16945 11095 17003 11101
rect 17494 11092 17500 11144
rect 17552 11092 17558 11144
rect 15194 11064 15200 11076
rect 12483 11036 12940 11064
rect 13004 11036 15200 11064
rect 12483 11033 12495 11036
rect 12437 11027 12495 11033
rect 12526 10996 12532 11008
rect 12360 10968 12532 10996
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 12912 10996 12940 11036
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 17218 11024 17224 11076
rect 17276 11064 17282 11076
rect 17604 11064 17632 11172
rect 19260 11141 19288 11172
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 19702 11160 19708 11212
rect 19760 11200 19766 11212
rect 20162 11200 20168 11212
rect 19760 11172 20168 11200
rect 19760 11160 19766 11172
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 24762 11200 24768 11212
rect 22848 11172 24768 11200
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11134 18475 11135
rect 19245 11135 19303 11141
rect 18463 11106 18552 11134
rect 18463 11101 18475 11106
rect 18417 11095 18475 11101
rect 17276 11036 17632 11064
rect 18524 11064 18552 11106
rect 19245 11101 19257 11135
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 20530 11132 20536 11144
rect 19475 11104 20536 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 20530 11092 20536 11104
rect 20588 11132 20594 11144
rect 20588 11104 20760 11132
rect 20588 11092 20594 11104
rect 20622 11064 20628 11076
rect 18524 11036 20628 11064
rect 17276 11024 17282 11036
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 20732 11064 20760 11104
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 22738 11092 22744 11144
rect 22796 11092 22802 11144
rect 22848 11064 22876 11172
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 26510 11160 26516 11212
rect 26568 11200 26574 11212
rect 26786 11200 26792 11212
rect 26568 11172 26792 11200
rect 26568 11160 26574 11172
rect 26786 11160 26792 11172
rect 26844 11160 26850 11212
rect 27798 11200 27804 11212
rect 27356 11172 27804 11200
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 20732 11036 22876 11064
rect 22940 11064 22968 11095
rect 23014 11092 23020 11144
rect 23072 11092 23078 11144
rect 23382 11092 23388 11144
rect 23440 11092 23446 11144
rect 27356 11132 27384 11172
rect 27798 11160 27804 11172
rect 27856 11160 27862 11212
rect 27893 11203 27951 11209
rect 27893 11169 27905 11203
rect 27939 11200 27951 11203
rect 28000 11200 28028 11240
rect 28534 11228 28540 11280
rect 28592 11268 28598 11280
rect 29917 11271 29975 11277
rect 29917 11268 29929 11271
rect 28592 11240 29929 11268
rect 28592 11228 28598 11240
rect 29917 11237 29929 11240
rect 29963 11237 29975 11271
rect 29917 11231 29975 11237
rect 31294 11228 31300 11280
rect 31352 11268 31358 11280
rect 31389 11271 31447 11277
rect 31389 11268 31401 11271
rect 31352 11240 31401 11268
rect 31352 11228 31358 11240
rect 31389 11237 31401 11240
rect 31435 11237 31447 11271
rect 31389 11231 31447 11237
rect 31662 11228 31668 11280
rect 31720 11268 31726 11280
rect 31720 11240 32260 11268
rect 31720 11228 31726 11240
rect 27939 11172 28028 11200
rect 28184 11172 29224 11200
rect 27939 11169 27951 11172
rect 27893 11163 27951 11169
rect 28184 11144 28212 11172
rect 23676 11104 27384 11132
rect 27433 11135 27491 11141
rect 23106 11064 23112 11076
rect 22940 11036 23112 11064
rect 23106 11024 23112 11036
rect 23164 11064 23170 11076
rect 23400 11064 23428 11092
rect 23676 11073 23704 11104
rect 27433 11101 27445 11135
rect 27479 11101 27491 11135
rect 27433 11095 27491 11101
rect 27617 11135 27675 11141
rect 27617 11101 27629 11135
rect 27663 11132 27675 11135
rect 27663 11104 27752 11132
rect 27663 11101 27675 11104
rect 27617 11095 27675 11101
rect 23661 11067 23719 11073
rect 23661 11064 23673 11067
rect 23164 11036 23336 11064
rect 23400 11036 23673 11064
rect 23164 11024 23170 11036
rect 13446 10996 13452 11008
rect 12912 10968 13452 10996
rect 13446 10956 13452 10968
rect 13504 10956 13510 11008
rect 14642 10956 14648 11008
rect 14700 10996 14706 11008
rect 17405 10999 17463 11005
rect 17405 10996 17417 10999
rect 14700 10968 17417 10996
rect 14700 10956 14706 10968
rect 17405 10965 17417 10968
rect 17451 10996 17463 10999
rect 18046 10996 18052 11008
rect 17451 10968 18052 10996
rect 17451 10965 17463 10968
rect 17405 10959 17463 10965
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 18230 10956 18236 11008
rect 18288 10956 18294 11008
rect 18506 10956 18512 11008
rect 18564 10996 18570 11008
rect 20254 10996 20260 11008
rect 18564 10968 20260 10996
rect 18564 10956 18570 10968
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 23308 11005 23336 11036
rect 23661 11033 23673 11036
rect 23707 11033 23719 11067
rect 23661 11027 23719 11033
rect 24394 11024 24400 11076
rect 24452 11024 24458 11076
rect 24581 11067 24639 11073
rect 24581 11033 24593 11067
rect 24627 11064 24639 11067
rect 24854 11064 24860 11076
rect 24627 11036 24860 11064
rect 24627 11033 24639 11036
rect 24581 11027 24639 11033
rect 24854 11024 24860 11036
rect 24912 11064 24918 11076
rect 25314 11064 25320 11076
rect 24912 11036 25320 11064
rect 24912 11024 24918 11036
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 27154 11024 27160 11076
rect 27212 11064 27218 11076
rect 27448 11064 27476 11095
rect 27212 11036 27476 11064
rect 27212 11024 27218 11036
rect 23293 10999 23351 11005
rect 23293 10965 23305 10999
rect 23339 10965 23351 10999
rect 23293 10959 23351 10965
rect 23461 10999 23519 11005
rect 23461 10965 23473 10999
rect 23507 10996 23519 10999
rect 23566 10996 23572 11008
rect 23507 10968 23572 10996
rect 23507 10965 23519 10968
rect 23461 10959 23519 10965
rect 23566 10956 23572 10968
rect 23624 10996 23630 11008
rect 24210 10996 24216 11008
rect 23624 10968 24216 10996
rect 23624 10956 23630 10968
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 27724 10996 27752 11104
rect 27982 11092 27988 11144
rect 28040 11092 28046 11144
rect 28166 11092 28172 11144
rect 28224 11092 28230 11144
rect 28350 11092 28356 11144
rect 28408 11092 28414 11144
rect 28810 11092 28816 11144
rect 28868 11132 28874 11144
rect 28905 11135 28963 11141
rect 28905 11132 28917 11135
rect 28868 11104 28917 11132
rect 28868 11092 28874 11104
rect 28905 11101 28917 11104
rect 28951 11101 28963 11135
rect 28905 11095 28963 11101
rect 28994 11092 29000 11144
rect 29052 11092 29058 11144
rect 29086 11092 29092 11144
rect 29144 11092 29150 11144
rect 29196 11141 29224 11172
rect 31938 11160 31944 11212
rect 31996 11160 32002 11212
rect 32232 11200 32260 11240
rect 32398 11228 32404 11280
rect 32456 11268 32462 11280
rect 32677 11271 32735 11277
rect 32677 11268 32689 11271
rect 32456 11240 32689 11268
rect 32456 11228 32462 11240
rect 32677 11237 32689 11240
rect 32723 11268 32735 11271
rect 32766 11268 32772 11280
rect 32723 11240 32772 11268
rect 32723 11237 32735 11240
rect 32677 11231 32735 11237
rect 32766 11228 32772 11240
rect 32824 11228 32830 11280
rect 32876 11200 32904 11308
rect 33042 11296 33048 11308
rect 33100 11296 33106 11348
rect 33134 11296 33140 11348
rect 33192 11336 33198 11348
rect 33229 11339 33287 11345
rect 33229 11336 33241 11339
rect 33192 11308 33241 11336
rect 33192 11296 33198 11308
rect 33229 11305 33241 11308
rect 33275 11305 33287 11339
rect 33229 11299 33287 11305
rect 34514 11296 34520 11348
rect 34572 11296 34578 11348
rect 34698 11296 34704 11348
rect 34756 11336 34762 11348
rect 34882 11336 34888 11348
rect 34756 11308 34888 11336
rect 34756 11296 34762 11308
rect 34882 11296 34888 11308
rect 34940 11296 34946 11348
rect 34532 11268 34560 11296
rect 34974 11268 34980 11280
rect 34532 11240 34980 11268
rect 34974 11228 34980 11240
rect 35032 11228 35038 11280
rect 32232 11172 32904 11200
rect 29181 11135 29239 11141
rect 29181 11101 29193 11135
rect 29227 11101 29239 11135
rect 29181 11095 29239 11101
rect 28261 11067 28319 11073
rect 28261 11033 28273 11067
rect 28307 11064 28319 11067
rect 28534 11064 28540 11076
rect 28307 11036 28540 11064
rect 28307 11033 28319 11036
rect 28261 11027 28319 11033
rect 28534 11024 28540 11036
rect 28592 11024 28598 11076
rect 28629 11067 28687 11073
rect 28629 11033 28641 11067
rect 28675 11064 28687 11067
rect 28675 11036 29040 11064
rect 28675 11033 28687 11036
rect 28629 11027 28687 11033
rect 29012 11008 29040 11036
rect 28442 10996 28448 11008
rect 27724 10968 28448 10996
rect 28442 10956 28448 10968
rect 28500 10956 28506 11008
rect 28718 10956 28724 11008
rect 28776 10956 28782 11008
rect 28994 10956 29000 11008
rect 29052 10956 29058 11008
rect 29104 10996 29132 11092
rect 29196 11064 29224 11095
rect 29546 11092 29552 11144
rect 29604 11092 29610 11144
rect 30101 11135 30159 11141
rect 30101 11101 30113 11135
rect 30147 11132 30159 11135
rect 31386 11132 31392 11144
rect 30147 11104 31392 11132
rect 30147 11101 30159 11104
rect 30101 11095 30159 11101
rect 31386 11092 31392 11104
rect 31444 11092 31450 11144
rect 31726 11132 31846 11148
rect 31588 11120 31892 11132
rect 31588 11104 31754 11120
rect 31818 11104 31892 11120
rect 31588 11076 31616 11104
rect 31570 11073 31576 11076
rect 31557 11067 31576 11073
rect 31557 11064 31569 11067
rect 29196 11036 31569 11064
rect 31557 11033 31569 11036
rect 31557 11027 31576 11033
rect 31570 11024 31576 11027
rect 31628 11024 31634 11076
rect 31662 11024 31668 11076
rect 31720 11064 31726 11076
rect 31757 11067 31815 11073
rect 31757 11064 31769 11067
rect 31720 11036 31769 11064
rect 31720 11024 31726 11036
rect 31757 11033 31769 11036
rect 31803 11033 31815 11067
rect 31864 11064 31892 11104
rect 32030 11092 32036 11144
rect 32088 11141 32094 11144
rect 32232 11141 32260 11172
rect 34514 11160 34520 11212
rect 34572 11200 34578 11212
rect 35069 11203 35127 11209
rect 35069 11200 35081 11203
rect 34572 11172 35081 11200
rect 34572 11160 34578 11172
rect 35069 11169 35081 11172
rect 35115 11169 35127 11203
rect 35069 11163 35127 11169
rect 32088 11135 32137 11141
rect 32088 11101 32091 11135
rect 32125 11101 32137 11135
rect 32088 11095 32137 11101
rect 32217 11135 32275 11141
rect 32217 11101 32229 11135
rect 32263 11101 32275 11135
rect 32217 11095 32275 11101
rect 32088 11092 32094 11095
rect 32306 11092 32312 11144
rect 32364 11092 32370 11144
rect 32401 11135 32459 11141
rect 32401 11101 32413 11135
rect 32447 11132 32459 11135
rect 32858 11132 32864 11144
rect 32447 11104 32864 11132
rect 32447 11101 32459 11104
rect 32401 11095 32459 11101
rect 32858 11092 32864 11104
rect 32916 11092 32922 11144
rect 34790 11092 34796 11144
rect 34848 11092 34854 11144
rect 35342 11092 35348 11144
rect 35400 11092 35406 11144
rect 32953 11067 33011 11073
rect 32953 11064 32965 11067
rect 31864 11036 32965 11064
rect 31757 11027 31815 11033
rect 32953 11033 32965 11036
rect 32999 11033 33011 11067
rect 32953 11027 33011 11033
rect 33042 11024 33048 11076
rect 33100 11024 33106 11076
rect 29546 10996 29552 11008
rect 29104 10968 29552 10996
rect 29546 10956 29552 10968
rect 29604 10956 29610 11008
rect 29730 10956 29736 11008
rect 29788 10956 29794 11008
rect 31846 10956 31852 11008
rect 31904 10996 31910 11008
rect 32861 10999 32919 11005
rect 32861 10996 32873 10999
rect 31904 10968 32873 10996
rect 31904 10956 31910 10968
rect 32861 10965 32873 10968
rect 32907 10965 32919 10999
rect 32861 10959 32919 10965
rect 1104 10906 36432 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 36432 10906
rect 1104 10832 36432 10854
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3418 10792 3424 10804
rect 3200 10764 3424 10792
rect 3200 10752 3206 10764
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 5442 10792 5448 10804
rect 5184 10764 5448 10792
rect 2958 10724 2964 10736
rect 2898 10696 2964 10724
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 3694 10684 3700 10736
rect 3752 10684 3758 10736
rect 5184 10724 5212 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5534 10752 5540 10804
rect 5592 10752 5598 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 7064 10764 7941 10792
rect 7064 10752 7070 10764
rect 7929 10761 7941 10764
rect 7975 10761 7987 10795
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 7929 10755 7987 10761
rect 8312 10764 9996 10792
rect 5552 10724 5580 10752
rect 4632 10696 5212 10724
rect 5276 10696 5580 10724
rect 1394 10616 1400 10668
rect 1452 10616 1458 10668
rect 3234 10616 3240 10668
rect 3292 10616 3298 10668
rect 3391 10659 3449 10665
rect 3391 10625 3403 10659
rect 3437 10656 3449 10659
rect 3602 10656 3608 10668
rect 3437 10628 3608 10656
rect 3437 10625 3449 10628
rect 3391 10619 3449 10625
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3936 10628 3985 10656
rect 3936 10616 3942 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 3786 10588 3792 10600
rect 1719 10560 3792 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 4632 10588 4660 10696
rect 4798 10616 4804 10668
rect 4856 10616 4862 10668
rect 5276 10665 5304 10696
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 8312 10724 8340 10764
rect 8570 10724 8576 10736
rect 5868 10696 8340 10724
rect 8404 10696 8576 10724
rect 5868 10684 5874 10696
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5445 10659 5503 10665
rect 5445 10625 5457 10659
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 3896 10560 4660 10588
rect 1670 10412 1676 10464
rect 1728 10452 1734 10464
rect 2314 10452 2320 10464
rect 1728 10424 2320 10452
rect 1728 10412 1734 10424
rect 2314 10412 2320 10424
rect 2372 10452 2378 10464
rect 3326 10452 3332 10464
rect 2372 10424 3332 10452
rect 2372 10412 2378 10424
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3421 10455 3479 10461
rect 3421 10421 3433 10455
rect 3467 10452 3479 10455
rect 3602 10452 3608 10464
rect 3467 10424 3608 10452
rect 3467 10421 3479 10424
rect 3421 10415 3479 10421
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 3896 10461 3924 10560
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 5460 10588 5488 10619
rect 4764 10560 5488 10588
rect 4764 10548 4770 10560
rect 5077 10523 5135 10529
rect 5077 10520 5089 10523
rect 3988 10492 5089 10520
rect 3988 10464 4016 10492
rect 5077 10489 5089 10492
rect 5123 10489 5135 10523
rect 5077 10483 5135 10489
rect 5258 10480 5264 10532
rect 5316 10520 5322 10532
rect 5552 10520 5580 10619
rect 8128 10588 8156 10619
rect 8294 10616 8300 10668
rect 8352 10616 8358 10668
rect 8404 10665 8432 10696
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 8754 10684 8760 10736
rect 8812 10724 8818 10736
rect 9968 10733 9996 10764
rect 10060 10764 10517 10792
rect 9953 10727 10011 10733
rect 8812 10696 9628 10724
rect 8812 10684 8818 10696
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 8527 10628 8800 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 8496 10588 8524 10619
rect 8128 10560 8524 10588
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10588 8631 10591
rect 8662 10588 8668 10600
rect 8619 10560 8668 10588
rect 8619 10557 8631 10560
rect 8573 10551 8631 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8772 10588 8800 10628
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 9180 10628 9229 10656
rect 9180 10616 9186 10628
rect 9217 10625 9229 10628
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 9398 10616 9404 10668
rect 9456 10616 9462 10668
rect 9490 10616 9496 10668
rect 9548 10616 9554 10668
rect 9600 10665 9628 10696
rect 9953 10693 9965 10727
rect 9999 10693 10011 10727
rect 9953 10687 10011 10693
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 10060 10656 10088 10764
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 10505 10755 10563 10761
rect 12710 10752 12716 10804
rect 12768 10792 12774 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 12768 10764 15025 10792
rect 12768 10752 12774 10764
rect 15013 10761 15025 10764
rect 15059 10761 15071 10795
rect 15013 10755 15071 10761
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21266 10792 21272 10804
rect 21140 10764 21272 10792
rect 21140 10752 21146 10764
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 21637 10795 21695 10801
rect 21637 10761 21649 10795
rect 21683 10792 21695 10795
rect 21818 10792 21824 10804
rect 21683 10764 21824 10792
rect 21683 10761 21695 10764
rect 21637 10755 21695 10761
rect 21818 10752 21824 10764
rect 21876 10752 21882 10804
rect 23842 10752 23848 10804
rect 23900 10792 23906 10804
rect 24029 10795 24087 10801
rect 24029 10792 24041 10795
rect 23900 10764 24041 10792
rect 23900 10752 23906 10764
rect 24029 10761 24041 10764
rect 24075 10761 24087 10795
rect 24029 10755 24087 10761
rect 24210 10752 24216 10804
rect 24268 10792 24274 10804
rect 25130 10792 25136 10804
rect 24268 10764 25136 10792
rect 24268 10752 24274 10764
rect 25130 10752 25136 10764
rect 25188 10792 25194 10804
rect 25225 10795 25283 10801
rect 25225 10792 25237 10795
rect 25188 10764 25237 10792
rect 25188 10752 25194 10764
rect 25225 10761 25237 10764
rect 25271 10761 25283 10795
rect 25225 10755 25283 10761
rect 25774 10752 25780 10804
rect 25832 10792 25838 10804
rect 27706 10792 27712 10804
rect 25832 10764 27712 10792
rect 25832 10752 25838 10764
rect 27706 10752 27712 10764
rect 27764 10752 27770 10804
rect 27798 10752 27804 10804
rect 27856 10792 27862 10804
rect 27893 10795 27951 10801
rect 27893 10792 27905 10795
rect 27856 10764 27905 10792
rect 27856 10752 27862 10764
rect 27893 10761 27905 10764
rect 27939 10792 27951 10795
rect 28350 10792 28356 10804
rect 27939 10764 28356 10792
rect 27939 10761 27951 10764
rect 27893 10755 27951 10761
rect 28350 10752 28356 10764
rect 28408 10752 28414 10804
rect 28810 10752 28816 10804
rect 28868 10792 28874 10804
rect 29365 10795 29423 10801
rect 29365 10792 29377 10795
rect 28868 10764 29377 10792
rect 28868 10752 28874 10764
rect 29365 10761 29377 10764
rect 29411 10761 29423 10795
rect 29365 10755 29423 10761
rect 29457 10795 29515 10801
rect 29457 10761 29469 10795
rect 29503 10792 29515 10795
rect 29503 10764 29592 10792
rect 29503 10761 29515 10764
rect 29457 10755 29515 10761
rect 10137 10727 10195 10733
rect 10137 10693 10149 10727
rect 10183 10724 10195 10727
rect 10410 10724 10416 10736
rect 10183 10696 10416 10724
rect 10183 10693 10195 10696
rect 10137 10687 10195 10693
rect 10410 10684 10416 10696
rect 10468 10684 10474 10736
rect 11974 10684 11980 10736
rect 12032 10724 12038 10736
rect 18506 10724 18512 10736
rect 12032 10696 18512 10724
rect 12032 10684 12038 10696
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 18693 10727 18751 10733
rect 18693 10693 18705 10727
rect 18739 10724 18751 10727
rect 18782 10724 18788 10736
rect 18739 10696 18788 10724
rect 18739 10693 18751 10696
rect 18693 10687 18751 10693
rect 18782 10684 18788 10696
rect 18840 10684 18846 10736
rect 20622 10684 20628 10736
rect 20680 10724 20686 10736
rect 20680 10696 20944 10724
rect 20680 10684 20686 10696
rect 9631 10628 10088 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 10318 10616 10324 10668
rect 10376 10616 10382 10668
rect 10686 10616 10692 10668
rect 10744 10616 10750 10668
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 10226 10588 10232 10600
rect 8772 10560 10232 10588
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 15212 10588 15240 10619
rect 15286 10616 15292 10668
rect 15344 10616 15350 10668
rect 15470 10616 15476 10668
rect 15528 10616 15534 10668
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10625 17647 10659
rect 17589 10619 17647 10625
rect 15562 10588 15568 10600
rect 15212 10560 15568 10588
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 6638 10520 6644 10532
rect 5316 10492 6644 10520
rect 5316 10480 5322 10492
rect 6638 10480 6644 10492
rect 6696 10520 6702 10532
rect 8110 10520 8116 10532
rect 6696 10492 8116 10520
rect 6696 10480 6702 10492
rect 8110 10480 8116 10492
rect 8168 10520 8174 10532
rect 12066 10520 12072 10532
rect 8168 10492 12072 10520
rect 8168 10480 8174 10492
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 3881 10455 3939 10461
rect 3881 10421 3893 10455
rect 3927 10421 3939 10455
rect 3881 10415 3939 10421
rect 3970 10412 3976 10464
rect 4028 10412 4034 10464
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4341 10455 4399 10461
rect 4341 10452 4353 10455
rect 4120 10424 4353 10452
rect 4120 10412 4126 10424
rect 4341 10421 4353 10424
rect 4387 10421 4399 10455
rect 4341 10415 4399 10421
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4890 10452 4896 10464
rect 4479 10424 4896 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 9125 10455 9183 10461
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 9490 10452 9496 10464
rect 9171 10424 9496 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9858 10412 9864 10464
rect 9916 10412 9922 10464
rect 15010 10412 15016 10464
rect 15068 10452 15074 10464
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 15068 10424 15209 10452
rect 15068 10412 15074 10424
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 15197 10415 15255 10421
rect 17402 10412 17408 10464
rect 17460 10412 17466 10464
rect 17604 10452 17632 10619
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17828 10628 17877 10656
rect 17828 10616 17834 10628
rect 17865 10625 17877 10628
rect 17911 10656 17923 10659
rect 17954 10656 17960 10668
rect 17911 10628 17960 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 18046 10616 18052 10668
rect 18104 10616 18110 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 18966 10656 18972 10668
rect 18371 10628 18972 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 19150 10616 19156 10668
rect 19208 10616 19214 10668
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19613 10659 19671 10665
rect 19613 10656 19625 10659
rect 19392 10628 19625 10656
rect 19392 10616 19398 10628
rect 19613 10625 19625 10628
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 20714 10616 20720 10668
rect 20772 10616 20778 10668
rect 20916 10665 20944 10696
rect 20990 10684 20996 10736
rect 21048 10724 21054 10736
rect 21048 10696 21220 10724
rect 21048 10684 21054 10696
rect 20901 10659 20959 10665
rect 20901 10625 20913 10659
rect 20947 10625 20959 10659
rect 20901 10619 20959 10625
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 18601 10591 18659 10597
rect 17736 10560 18552 10588
rect 17736 10548 17742 10560
rect 17773 10523 17831 10529
rect 17773 10489 17785 10523
rect 17819 10520 17831 10523
rect 18141 10523 18199 10529
rect 18141 10520 18153 10523
rect 17819 10492 18153 10520
rect 17819 10489 17831 10492
rect 17773 10483 17831 10489
rect 18141 10489 18153 10492
rect 18187 10489 18199 10523
rect 18524 10520 18552 10560
rect 18601 10557 18613 10591
rect 18647 10588 18659 10591
rect 18690 10588 18696 10600
rect 18647 10560 18696 10588
rect 18647 10557 18659 10560
rect 18601 10551 18659 10557
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 19061 10591 19119 10597
rect 19061 10557 19073 10591
rect 19107 10588 19119 10591
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19107 10560 19441 10588
rect 19107 10557 19119 10560
rect 19061 10551 19119 10557
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 19518 10548 19524 10600
rect 19576 10588 19582 10600
rect 19886 10588 19892 10600
rect 19576 10560 19892 10588
rect 19576 10548 19582 10560
rect 19886 10548 19892 10560
rect 19944 10548 19950 10600
rect 19337 10523 19395 10529
rect 18524 10492 19288 10520
rect 18141 10483 18199 10489
rect 17862 10452 17868 10464
rect 17604 10424 17868 10452
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 18322 10412 18328 10464
rect 18380 10452 18386 10464
rect 18506 10452 18512 10464
rect 18380 10424 18512 10452
rect 18380 10412 18386 10424
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 19058 10412 19064 10464
rect 19116 10412 19122 10464
rect 19260 10452 19288 10492
rect 19337 10489 19349 10523
rect 19383 10520 19395 10523
rect 20625 10523 20683 10529
rect 20625 10520 20637 10523
rect 19383 10492 20637 10520
rect 19383 10489 19395 10492
rect 19337 10483 19395 10489
rect 20625 10489 20637 10492
rect 20671 10489 20683 10523
rect 20916 10520 20944 10619
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 21192 10665 21220 10696
rect 22922 10684 22928 10736
rect 22980 10684 22986 10736
rect 24397 10727 24455 10733
rect 24397 10693 24409 10727
rect 24443 10693 24455 10727
rect 24397 10687 24455 10693
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10656 21235 10659
rect 21266 10656 21272 10668
rect 21223 10628 21272 10656
rect 21223 10625 21235 10628
rect 21177 10619 21235 10625
rect 21266 10616 21272 10628
rect 21324 10616 21330 10668
rect 21450 10616 21456 10668
rect 21508 10616 21514 10668
rect 23106 10616 23112 10668
rect 23164 10616 23170 10668
rect 24412 10656 24440 10687
rect 24762 10684 24768 10736
rect 24820 10724 24826 10736
rect 28261 10727 28319 10733
rect 28261 10724 28273 10727
rect 24820 10696 28273 10724
rect 24820 10684 24826 10696
rect 28261 10693 28273 10696
rect 28307 10693 28319 10727
rect 28261 10687 28319 10693
rect 28902 10684 28908 10736
rect 28960 10724 28966 10736
rect 29089 10727 29147 10733
rect 29089 10724 29101 10727
rect 28960 10696 29101 10724
rect 28960 10684 28966 10696
rect 29089 10693 29101 10696
rect 29135 10693 29147 10727
rect 29564 10724 29592 10764
rect 29638 10752 29644 10804
rect 29696 10752 29702 10804
rect 30193 10795 30251 10801
rect 30193 10792 30205 10795
rect 29840 10764 30205 10792
rect 29840 10736 29868 10764
rect 30193 10761 30205 10764
rect 30239 10761 30251 10795
rect 30193 10755 30251 10761
rect 31662 10752 31668 10804
rect 31720 10792 31726 10804
rect 31720 10764 31800 10792
rect 31720 10752 31726 10764
rect 29822 10724 29828 10736
rect 29564 10696 29828 10724
rect 29089 10687 29147 10693
rect 29822 10684 29828 10696
rect 29880 10684 29886 10736
rect 29917 10727 29975 10733
rect 29917 10693 29929 10727
rect 29963 10724 29975 10727
rect 30742 10724 30748 10736
rect 29963 10696 30748 10724
rect 29963 10693 29975 10696
rect 29917 10687 29975 10693
rect 30742 10684 30748 10696
rect 30800 10724 30806 10736
rect 31110 10724 31116 10736
rect 30800 10696 31116 10724
rect 30800 10684 30806 10696
rect 31110 10684 31116 10696
rect 31168 10684 31174 10736
rect 31772 10724 31800 10764
rect 32398 10752 32404 10804
rect 32456 10752 32462 10804
rect 31313 10696 31800 10724
rect 24578 10656 24584 10668
rect 24412 10628 24584 10656
rect 24578 10616 24584 10628
rect 24636 10656 24642 10668
rect 27985 10659 28043 10665
rect 27985 10656 27997 10659
rect 24636 10628 27997 10656
rect 24636 10616 24642 10628
rect 27985 10625 27997 10628
rect 28031 10656 28043 10659
rect 28074 10656 28080 10668
rect 28031 10628 28080 10656
rect 28031 10625 28043 10628
rect 27985 10619 28043 10625
rect 28074 10616 28080 10628
rect 28132 10616 28138 10668
rect 28718 10616 28724 10668
rect 28776 10616 28782 10668
rect 28994 10616 29000 10668
rect 29052 10616 29058 10668
rect 29273 10659 29331 10665
rect 29273 10625 29285 10659
rect 29319 10656 29331 10659
rect 29472 10656 29592 10660
rect 29730 10656 29736 10668
rect 29319 10632 29736 10656
rect 29319 10628 29500 10632
rect 29564 10628 29736 10632
rect 29319 10625 29331 10628
rect 29273 10619 29331 10625
rect 29730 10616 29736 10628
rect 29788 10616 29794 10668
rect 30374 10616 30380 10668
rect 30432 10656 30438 10668
rect 31313 10656 31341 10696
rect 30432 10628 31341 10656
rect 30432 10616 30438 10628
rect 31662 10616 31668 10668
rect 31720 10616 31726 10668
rect 20990 10548 20996 10600
rect 21048 10588 21054 10600
rect 21361 10591 21419 10597
rect 21361 10588 21373 10591
rect 21048 10560 21373 10588
rect 21048 10548 21054 10560
rect 21361 10557 21373 10560
rect 21407 10588 21419 10591
rect 22738 10588 22744 10600
rect 21407 10560 22744 10588
rect 21407 10557 21419 10560
rect 21361 10551 21419 10557
rect 22738 10548 22744 10560
rect 22796 10548 22802 10600
rect 23293 10591 23351 10597
rect 23293 10557 23305 10591
rect 23339 10588 23351 10591
rect 23842 10588 23848 10600
rect 23339 10560 23848 10588
rect 23339 10557 23351 10560
rect 23293 10551 23351 10557
rect 23842 10548 23848 10560
rect 23900 10548 23906 10600
rect 25685 10591 25743 10597
rect 25685 10557 25697 10591
rect 25731 10588 25743 10591
rect 27614 10588 27620 10600
rect 25731 10560 27620 10588
rect 25731 10557 25743 10560
rect 25685 10551 25743 10557
rect 27614 10548 27620 10560
rect 27672 10588 27678 10600
rect 28534 10588 28540 10600
rect 27672 10560 28540 10588
rect 27672 10548 27678 10560
rect 28534 10548 28540 10560
rect 28592 10588 28598 10600
rect 28810 10588 28816 10600
rect 28592 10560 28816 10588
rect 28592 10548 28598 10560
rect 28810 10548 28816 10560
rect 28868 10548 28874 10600
rect 29546 10548 29552 10600
rect 29604 10588 29610 10600
rect 30558 10588 30564 10600
rect 29604 10560 30564 10588
rect 29604 10548 29610 10560
rect 30558 10548 30564 10560
rect 30616 10588 30622 10600
rect 31570 10588 31576 10600
rect 30616 10560 31576 10588
rect 30616 10548 30622 10560
rect 31570 10548 31576 10560
rect 31628 10548 31634 10600
rect 31772 10588 31800 10696
rect 31864 10696 32719 10724
rect 31864 10665 31892 10696
rect 31849 10659 31907 10665
rect 31849 10625 31861 10659
rect 31895 10625 31907 10659
rect 31849 10619 31907 10625
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10656 32367 10659
rect 32398 10656 32404 10668
rect 32355 10628 32404 10656
rect 32355 10625 32367 10628
rect 32309 10619 32367 10625
rect 32324 10588 32352 10619
rect 32398 10616 32404 10628
rect 32456 10616 32462 10668
rect 32691 10665 32719 10696
rect 32766 10684 32772 10736
rect 32824 10724 32830 10736
rect 32824 10696 33088 10724
rect 32824 10684 32830 10696
rect 32493 10659 32551 10665
rect 32493 10625 32505 10659
rect 32539 10625 32551 10659
rect 32493 10619 32551 10625
rect 32677 10659 32735 10665
rect 32677 10625 32689 10659
rect 32723 10646 32735 10659
rect 32723 10625 32812 10646
rect 32677 10619 32812 10625
rect 31772 10560 32352 10588
rect 20916 10492 22094 10520
rect 20625 10483 20683 10489
rect 19797 10455 19855 10461
rect 19797 10452 19809 10455
rect 19260 10424 19809 10452
rect 19797 10421 19809 10424
rect 19843 10452 19855 10455
rect 19886 10452 19892 10464
rect 19843 10424 19892 10452
rect 19843 10421 19855 10424
rect 19797 10415 19855 10421
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 20254 10412 20260 10464
rect 20312 10452 20318 10464
rect 20349 10455 20407 10461
rect 20349 10452 20361 10455
rect 20312 10424 20361 10452
rect 20312 10412 20318 10424
rect 20349 10421 20361 10424
rect 20395 10421 20407 10455
rect 20349 10415 20407 10421
rect 20806 10412 20812 10464
rect 20864 10412 20870 10464
rect 20990 10412 20996 10464
rect 21048 10452 21054 10464
rect 21177 10455 21235 10461
rect 21177 10452 21189 10455
rect 21048 10424 21189 10452
rect 21048 10412 21054 10424
rect 21177 10421 21189 10424
rect 21223 10421 21235 10455
rect 22066 10452 22094 10492
rect 22554 10480 22560 10532
rect 22612 10520 22618 10532
rect 24762 10520 24768 10532
rect 22612 10492 24768 10520
rect 22612 10480 22618 10492
rect 24762 10480 24768 10492
rect 24820 10480 24826 10532
rect 25409 10523 25467 10529
rect 25409 10489 25421 10523
rect 25455 10520 25467 10523
rect 27522 10520 27528 10532
rect 25455 10492 27528 10520
rect 25455 10489 25467 10492
rect 25409 10483 25467 10489
rect 27522 10480 27528 10492
rect 27580 10480 27586 10532
rect 28905 10523 28963 10529
rect 28905 10489 28917 10523
rect 28951 10520 28963 10523
rect 29086 10520 29092 10532
rect 28951 10492 29092 10520
rect 28951 10489 28963 10492
rect 28905 10483 28963 10489
rect 29086 10480 29092 10492
rect 29144 10480 29150 10532
rect 31754 10480 31760 10532
rect 31812 10520 31818 10532
rect 31849 10523 31907 10529
rect 31849 10520 31861 10523
rect 31812 10492 31861 10520
rect 31812 10480 31818 10492
rect 31849 10489 31861 10492
rect 31895 10489 31907 10523
rect 31849 10483 31907 10489
rect 23842 10452 23848 10464
rect 22066 10424 23848 10452
rect 21177 10415 21235 10421
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 24213 10455 24271 10461
rect 24213 10421 24225 10455
rect 24259 10452 24271 10455
rect 24394 10452 24400 10464
rect 24259 10424 24400 10452
rect 24259 10421 24271 10424
rect 24213 10415 24271 10421
rect 24394 10412 24400 10424
rect 24452 10412 24458 10464
rect 26234 10412 26240 10464
rect 26292 10452 26298 10464
rect 26602 10452 26608 10464
rect 26292 10424 26608 10452
rect 26292 10412 26298 10424
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 28074 10412 28080 10464
rect 28132 10452 28138 10464
rect 28442 10452 28448 10464
rect 28132 10424 28448 10452
rect 28132 10412 28138 10424
rect 28442 10412 28448 10424
rect 28500 10412 28506 10464
rect 29178 10412 29184 10464
rect 29236 10452 29242 10464
rect 29546 10452 29552 10464
rect 29236 10424 29552 10452
rect 29236 10412 29242 10424
rect 29546 10412 29552 10424
rect 29604 10452 29610 10464
rect 30009 10455 30067 10461
rect 30009 10452 30021 10455
rect 29604 10424 30021 10452
rect 29604 10412 29610 10424
rect 30009 10421 30021 10424
rect 30055 10452 30067 10455
rect 30282 10452 30288 10464
rect 30055 10424 30288 10452
rect 30055 10421 30067 10424
rect 30009 10415 30067 10421
rect 30282 10412 30288 10424
rect 30340 10412 30346 10464
rect 32508 10452 32536 10619
rect 32691 10618 32812 10619
rect 32784 10520 32812 10618
rect 32858 10616 32864 10668
rect 32916 10616 32922 10668
rect 33060 10665 33088 10696
rect 34422 10684 34428 10736
rect 34480 10724 34486 10736
rect 34517 10727 34575 10733
rect 34517 10724 34529 10727
rect 34480 10696 34529 10724
rect 34480 10684 34486 10696
rect 34517 10693 34529 10696
rect 34563 10693 34575 10727
rect 34517 10687 34575 10693
rect 34974 10684 34980 10736
rect 35032 10684 35038 10736
rect 33045 10659 33103 10665
rect 33045 10625 33057 10659
rect 33091 10625 33103 10659
rect 33045 10619 33103 10625
rect 33502 10548 33508 10600
rect 33560 10588 33566 10600
rect 34241 10591 34299 10597
rect 34241 10588 34253 10591
rect 33560 10560 34253 10588
rect 33560 10548 33566 10560
rect 34241 10557 34253 10560
rect 34287 10557 34299 10591
rect 34241 10551 34299 10557
rect 34146 10520 34152 10532
rect 32784 10492 34152 10520
rect 34146 10480 34152 10492
rect 34204 10480 34210 10532
rect 33229 10455 33287 10461
rect 33229 10452 33241 10455
rect 32508 10424 33241 10452
rect 33229 10421 33241 10424
rect 33275 10452 33287 10455
rect 33410 10452 33416 10464
rect 33275 10424 33416 10452
rect 33275 10421 33287 10424
rect 33229 10415 33287 10421
rect 33410 10412 33416 10424
rect 33468 10412 33474 10464
rect 34330 10412 34336 10464
rect 34388 10452 34394 10464
rect 34974 10452 34980 10464
rect 34388 10424 34980 10452
rect 34388 10412 34394 10424
rect 34974 10412 34980 10424
rect 35032 10412 35038 10464
rect 35526 10412 35532 10464
rect 35584 10452 35590 10464
rect 35989 10455 36047 10461
rect 35989 10452 36001 10455
rect 35584 10424 36001 10452
rect 35584 10412 35590 10424
rect 35989 10421 36001 10424
rect 36035 10421 36047 10455
rect 35989 10415 36047 10421
rect 1104 10362 36432 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 36432 10362
rect 1104 10288 36432 10310
rect 1765 10251 1823 10257
rect 1765 10217 1777 10251
rect 1811 10248 1823 10251
rect 2590 10248 2596 10260
rect 1811 10220 2596 10248
rect 1811 10217 1823 10220
rect 1765 10211 1823 10217
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 3786 10208 3792 10260
rect 3844 10208 3850 10260
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 3936 10220 4721 10248
rect 3936 10208 3942 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 5960 10220 6960 10248
rect 5960 10208 5966 10220
rect 6932 10192 6960 10220
rect 8496 10220 11713 10248
rect 2866 10180 2872 10192
rect 1964 10152 2872 10180
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 1964 10053 1992 10152
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 3234 10140 3240 10192
rect 3292 10180 3298 10192
rect 4890 10180 4896 10192
rect 3292 10152 4896 10180
rect 3292 10140 3298 10152
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2317 10115 2375 10121
rect 2317 10112 2329 10115
rect 2087 10084 2329 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 2317 10081 2329 10084
rect 2363 10081 2375 10115
rect 2317 10075 2375 10081
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 1949 10007 2007 10013
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10013 2191 10047
rect 2133 10007 2191 10013
rect 1872 9976 1900 10007
rect 2148 9976 2176 10007
rect 2406 10004 2412 10056
rect 2464 10004 2470 10056
rect 3344 10053 3372 10152
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 5994 10180 6000 10192
rect 5828 10152 6000 10180
rect 3602 10072 3608 10124
rect 3660 10112 3666 10124
rect 3660 10084 4108 10112
rect 3660 10072 3666 10084
rect 3328 10047 3386 10053
rect 3328 10013 3340 10047
rect 3374 10013 3386 10047
rect 3328 10007 3386 10013
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 3878 10044 3884 10056
rect 3476 10016 3884 10044
rect 3476 10004 3482 10016
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 3970 10004 3976 10056
rect 4028 10004 4034 10056
rect 4080 10053 4108 10084
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5408 10084 5580 10112
rect 5408 10072 5414 10084
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 4154 10004 4160 10056
rect 4212 10004 4218 10056
rect 4246 10004 4252 10056
rect 4304 10053 4310 10056
rect 4304 10047 4333 10053
rect 4321 10013 4333 10047
rect 4304 10007 4333 10013
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4304 10004 4310 10007
rect 2498 9976 2504 9988
rect 1872 9948 1992 9976
rect 2148 9948 2504 9976
rect 1964 9908 1992 9948
rect 2498 9936 2504 9948
rect 2556 9976 2562 9988
rect 3053 9979 3111 9985
rect 3053 9976 3065 9979
rect 2556 9948 3065 9976
rect 2556 9936 2562 9948
rect 3053 9945 3065 9948
rect 3099 9945 3111 9979
rect 3053 9939 3111 9945
rect 3142 9936 3148 9988
rect 3200 9976 3206 9988
rect 3200 9948 4200 9976
rect 3200 9936 3206 9948
rect 2406 9908 2412 9920
rect 1964 9880 2412 9908
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 2777 9911 2835 9917
rect 2777 9877 2789 9911
rect 2823 9908 2835 9911
rect 3970 9908 3976 9920
rect 2823 9880 3976 9908
rect 2823 9877 2835 9880
rect 2777 9871 2835 9877
rect 3970 9868 3976 9880
rect 4028 9868 4034 9920
rect 4172 9908 4200 9948
rect 4448 9908 4476 10007
rect 4706 10004 4712 10056
rect 4764 10004 4770 10056
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5552 10053 5580 10084
rect 5828 10053 5856 10152
rect 5994 10140 6000 10152
rect 6052 10180 6058 10192
rect 6457 10183 6515 10189
rect 6457 10180 6469 10183
rect 6052 10152 6469 10180
rect 6052 10140 6058 10152
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 4948 10016 5089 10044
rect 4948 10004 4954 10016
rect 5077 10013 5089 10016
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 5538 10047 5596 10053
rect 5538 10013 5550 10047
rect 5584 10013 5596 10047
rect 5538 10007 5596 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 5460 9976 5488 10007
rect 5902 10004 5908 10056
rect 5960 10053 5966 10056
rect 5960 10044 5968 10053
rect 6104 10044 6132 10152
rect 6457 10149 6469 10152
rect 6503 10149 6515 10183
rect 6457 10143 6515 10149
rect 6914 10140 6920 10192
rect 6972 10180 6978 10192
rect 8294 10180 8300 10192
rect 6972 10152 8300 10180
rect 6972 10140 6978 10152
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 8496 10180 8524 10220
rect 11701 10217 11713 10220
rect 11747 10217 11759 10251
rect 11701 10211 11759 10217
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12345 10251 12403 10257
rect 12345 10248 12357 10251
rect 12124 10220 12357 10248
rect 12124 10208 12130 10220
rect 12345 10217 12357 10220
rect 12391 10217 12403 10251
rect 12345 10211 12403 10217
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10217 12587 10251
rect 12529 10211 12587 10217
rect 14737 10251 14795 10257
rect 14737 10217 14749 10251
rect 14783 10248 14795 10251
rect 15470 10248 15476 10260
rect 14783 10220 15476 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 8404 10152 8524 10180
rect 10781 10183 10839 10189
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6362 10112 6368 10124
rect 6227 10084 6368 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 6362 10072 6368 10084
rect 6420 10112 6426 10124
rect 8404 10112 8432 10152
rect 10781 10149 10793 10183
rect 10827 10180 10839 10183
rect 11882 10180 11888 10192
rect 10827 10152 11888 10180
rect 10827 10149 10839 10152
rect 10781 10143 10839 10149
rect 6420 10084 6868 10112
rect 6420 10072 6426 10084
rect 6840 10053 6868 10084
rect 7484 10084 8432 10112
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 5960 10016 6005 10044
rect 6104 10016 6745 10044
rect 5960 10007 5968 10016
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 6826 10047 6884 10053
rect 6826 10013 6838 10047
rect 6872 10013 6884 10047
rect 7484 10044 7512 10084
rect 6826 10007 6884 10013
rect 7116 10016 7512 10044
rect 7561 10047 7619 10053
rect 5960 10004 5966 10007
rect 5626 9976 5632 9988
rect 5460 9948 5632 9976
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 5718 9936 5724 9988
rect 5776 9976 5782 9988
rect 6270 9976 6276 9988
rect 5776 9948 6276 9976
rect 5776 9936 5782 9948
rect 6270 9936 6276 9948
rect 6328 9976 6334 9988
rect 7116 9976 7144 10016
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 7650 10044 7656 10056
rect 7607 10016 7656 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 7650 10004 7656 10016
rect 7708 10044 7714 10056
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 7708 10016 7757 10044
rect 7708 10004 7714 10016
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 7834 10004 7840 10056
rect 7892 10044 7898 10056
rect 7929 10047 7987 10053
rect 7929 10044 7941 10047
rect 7892 10016 7941 10044
rect 7892 10004 7898 10016
rect 7929 10013 7941 10016
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 8404 10053 8432 10084
rect 8754 10072 8760 10124
rect 8812 10112 8818 10124
rect 9030 10112 9036 10124
rect 8812 10084 9036 10112
rect 8812 10072 8818 10084
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 11256 10121 11284 10152
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 12544 10124 12572 10211
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 17405 10251 17463 10257
rect 17405 10248 17417 10251
rect 15620 10220 17417 10248
rect 15620 10208 15626 10220
rect 17405 10217 17417 10220
rect 17451 10217 17463 10251
rect 17405 10211 17463 10217
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 20070 10248 20076 10260
rect 19668 10220 20076 10248
rect 19668 10208 19674 10220
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20806 10208 20812 10260
rect 20864 10208 20870 10260
rect 20990 10208 20996 10260
rect 21048 10208 21054 10260
rect 22646 10208 22652 10260
rect 22704 10248 22710 10260
rect 23017 10251 23075 10257
rect 23017 10248 23029 10251
rect 22704 10220 23029 10248
rect 22704 10208 22710 10220
rect 23017 10217 23029 10220
rect 23063 10217 23075 10251
rect 23017 10211 23075 10217
rect 23198 10208 23204 10260
rect 23256 10248 23262 10260
rect 24394 10248 24400 10260
rect 23256 10220 24400 10248
rect 23256 10208 23262 10220
rect 24394 10208 24400 10220
rect 24452 10208 24458 10260
rect 24486 10208 24492 10260
rect 24544 10208 24550 10260
rect 25038 10208 25044 10260
rect 25096 10208 25102 10260
rect 25498 10208 25504 10260
rect 25556 10248 25562 10260
rect 25774 10248 25780 10260
rect 25556 10220 25780 10248
rect 25556 10208 25562 10220
rect 25774 10208 25780 10220
rect 25832 10208 25838 10260
rect 26881 10251 26939 10257
rect 26881 10217 26893 10251
rect 26927 10217 26939 10251
rect 26881 10211 26939 10217
rect 17034 10180 17040 10192
rect 15258 10152 17040 10180
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 11664 10084 12081 10112
rect 11664 10072 11670 10084
rect 12069 10081 12081 10084
rect 12115 10112 12127 10115
rect 12526 10112 12532 10124
rect 12115 10084 12532 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 15258 10112 15286 10152
rect 17034 10140 17040 10152
rect 17092 10140 17098 10192
rect 17773 10183 17831 10189
rect 17773 10149 17785 10183
rect 17819 10180 17831 10183
rect 18598 10180 18604 10192
rect 17819 10152 18604 10180
rect 17819 10149 17831 10152
rect 17773 10143 17831 10149
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 19978 10140 19984 10192
rect 20036 10180 20042 10192
rect 21008 10180 21036 10208
rect 26697 10183 26755 10189
rect 26697 10180 26709 10183
rect 20036 10152 21036 10180
rect 22388 10152 26709 10180
rect 20036 10140 20042 10152
rect 22388 10112 22416 10152
rect 26697 10149 26709 10152
rect 26743 10149 26755 10183
rect 26697 10143 26755 10149
rect 13964 10084 15286 10112
rect 15488 10084 22416 10112
rect 13964 10072 13970 10084
rect 8206 10047 8264 10053
rect 8206 10013 8218 10047
rect 8252 10013 8264 10047
rect 8206 10007 8264 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8617 10047 8675 10053
rect 8617 10013 8629 10047
rect 8663 10044 8675 10047
rect 8938 10044 8944 10056
rect 8663 10016 8944 10044
rect 8663 10013 8675 10016
rect 8617 10007 8675 10013
rect 6328 9948 7144 9976
rect 6328 9936 6334 9948
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 8220 9976 8248 10007
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 10686 10044 10692 10056
rect 10442 10016 10692 10044
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 10870 10004 10876 10056
rect 10928 10004 10934 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10044 11115 10047
rect 11514 10044 11520 10056
rect 11103 10016 11520 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 12250 10044 12256 10056
rect 11931 10016 12256 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 13446 10004 13452 10056
rect 13504 10044 13510 10056
rect 14921 10047 14979 10053
rect 14921 10044 14933 10047
rect 13504 10016 14933 10044
rect 13504 10004 13510 10016
rect 14921 10013 14933 10016
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 8294 9976 8300 9988
rect 7248 9948 7880 9976
rect 8220 9948 8300 9976
rect 7248 9936 7254 9948
rect 4172 9880 4476 9908
rect 4525 9911 4583 9917
rect 4525 9877 4537 9911
rect 4571 9908 4583 9911
rect 4706 9908 4712 9920
rect 4571 9880 4712 9908
rect 4571 9877 4583 9880
rect 4525 9871 4583 9877
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 5902 9868 5908 9920
rect 5960 9908 5966 9920
rect 6089 9911 6147 9917
rect 6089 9908 6101 9911
rect 5960 9880 6101 9908
rect 5960 9868 5966 9880
rect 6089 9877 6101 9880
rect 6135 9877 6147 9911
rect 6089 9871 6147 9877
rect 6546 9868 6552 9920
rect 6604 9908 6610 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6604 9880 6653 9908
rect 6604 9868 6610 9880
rect 6641 9877 6653 9880
rect 6687 9877 6699 9911
rect 6641 9871 6699 9877
rect 7098 9868 7104 9920
rect 7156 9868 7162 9920
rect 7466 9868 7472 9920
rect 7524 9868 7530 9920
rect 7852 9917 7880 9948
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 8478 9936 8484 9988
rect 8536 9936 8542 9988
rect 9306 9936 9312 9988
rect 9364 9936 9370 9988
rect 12710 9936 12716 9988
rect 12768 9936 12774 9988
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 14936 9976 14964 10007
rect 15010 10004 15016 10056
rect 15068 10004 15074 10056
rect 15212 10053 15240 10084
rect 15197 10047 15255 10053
rect 15197 10013 15209 10047
rect 15243 10013 15255 10047
rect 15197 10007 15255 10013
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10044 15347 10047
rect 15378 10044 15384 10056
rect 15335 10016 15384 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 15488 9976 15516 10084
rect 22462 10072 22468 10124
rect 22520 10112 22526 10124
rect 25593 10115 25651 10121
rect 25593 10112 25605 10115
rect 22520 10084 25605 10112
rect 22520 10072 22526 10084
rect 25593 10081 25605 10084
rect 25639 10112 25651 10115
rect 26050 10112 26056 10124
rect 25639 10084 26056 10112
rect 25639 10081 25651 10084
rect 25593 10075 25651 10081
rect 26050 10072 26056 10084
rect 26108 10072 26114 10124
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 12860 9948 14688 9976
rect 14936 9948 15516 9976
rect 17604 9976 17632 10007
rect 17770 10004 17776 10056
rect 17828 10044 17834 10056
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17828 10016 17877 10044
rect 17828 10004 17834 10016
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 18141 10047 18199 10053
rect 18141 10013 18153 10047
rect 18187 10044 18199 10047
rect 18230 10044 18236 10056
rect 18187 10016 18236 10044
rect 18187 10013 18199 10016
rect 18141 10007 18199 10013
rect 18156 9976 18184 10007
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 21085 10047 21143 10053
rect 21085 10013 21097 10047
rect 21131 10013 21143 10047
rect 21085 10007 21143 10013
rect 17604 9948 18184 9976
rect 21100 9976 21128 10007
rect 21174 10004 21180 10056
rect 21232 10004 21238 10056
rect 21542 10004 21548 10056
rect 21600 10044 21606 10056
rect 24673 10047 24731 10053
rect 24673 10044 24685 10047
rect 21600 10016 24685 10044
rect 21600 10004 21606 10016
rect 21450 9976 21456 9988
rect 21100 9948 21456 9976
rect 12860 9936 12866 9948
rect 7837 9911 7895 9917
rect 7837 9877 7849 9911
rect 7883 9908 7895 9911
rect 8110 9908 8116 9920
rect 7883 9880 8116 9908
rect 7883 9877 7895 9880
rect 7837 9871 7895 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 8757 9911 8815 9917
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 8938 9908 8944 9920
rect 8803 9880 8944 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 12513 9911 12571 9917
rect 12513 9877 12525 9911
rect 12559 9908 12571 9911
rect 14550 9908 14556 9920
rect 12559 9880 14556 9908
rect 12559 9877 12571 9880
rect 12513 9871 12571 9877
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 14660 9908 14688 9948
rect 17880 9920 17908 9948
rect 21450 9936 21456 9948
rect 21508 9936 21514 9988
rect 23385 9979 23443 9985
rect 23385 9945 23397 9979
rect 23431 9976 23443 9979
rect 23842 9976 23848 9988
rect 23431 9948 23848 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 23842 9936 23848 9948
rect 23900 9936 23906 9988
rect 17402 9908 17408 9920
rect 14660 9880 17408 9908
rect 17402 9868 17408 9880
rect 17460 9868 17466 9920
rect 17862 9868 17868 9920
rect 17920 9868 17926 9920
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18325 9911 18383 9917
rect 18325 9908 18337 9911
rect 18104 9880 18337 9908
rect 18104 9868 18110 9880
rect 18325 9877 18337 9880
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 23201 9911 23259 9917
rect 23201 9908 23213 9911
rect 22980 9880 23213 9908
rect 22980 9868 22986 9880
rect 23201 9877 23213 9880
rect 23247 9877 23259 9911
rect 24320 9908 24348 10016
rect 24673 10013 24685 10016
rect 24719 10013 24731 10047
rect 24673 10007 24731 10013
rect 24854 10004 24860 10056
rect 24912 10004 24918 10056
rect 25314 10004 25320 10056
rect 25372 10004 25378 10056
rect 25406 10004 25412 10056
rect 25464 10004 25470 10056
rect 25777 10047 25835 10053
rect 25777 10013 25789 10047
rect 25823 10044 25835 10047
rect 25869 10047 25927 10053
rect 25869 10044 25881 10047
rect 25823 10016 25881 10044
rect 25823 10013 25835 10016
rect 25777 10007 25835 10013
rect 25869 10013 25881 10016
rect 25915 10044 25927 10047
rect 25958 10044 25964 10056
rect 25915 10016 25964 10044
rect 25915 10013 25927 10016
rect 25869 10007 25927 10013
rect 24394 9936 24400 9988
rect 24452 9976 24458 9988
rect 25332 9976 25360 10004
rect 24452 9948 25360 9976
rect 24452 9936 24458 9948
rect 25792 9908 25820 10007
rect 25958 10004 25964 10016
rect 26016 10004 26022 10056
rect 26234 10004 26240 10056
rect 26292 10004 26298 10056
rect 26896 10044 26924 10211
rect 26970 10208 26976 10260
rect 27028 10248 27034 10260
rect 27028 10220 29960 10248
rect 27028 10208 27034 10220
rect 27522 10140 27528 10192
rect 27580 10180 27586 10192
rect 27580 10152 27936 10180
rect 27580 10140 27586 10152
rect 27157 10115 27215 10121
rect 27157 10081 27169 10115
rect 27203 10112 27215 10115
rect 27246 10112 27252 10124
rect 27203 10084 27252 10112
rect 27203 10081 27215 10084
rect 27157 10075 27215 10081
rect 26344 10016 26924 10044
rect 26050 9936 26056 9988
rect 26108 9976 26114 9988
rect 26344 9976 26372 10016
rect 26970 10004 26976 10056
rect 27028 10004 27034 10056
rect 27062 10004 27068 10056
rect 27120 10004 27126 10056
rect 26108 9948 26372 9976
rect 26108 9936 26114 9948
rect 26510 9936 26516 9988
rect 26568 9976 26574 9988
rect 27172 9976 27200 10075
rect 27246 10072 27252 10084
rect 27304 10072 27310 10124
rect 27433 10115 27491 10121
rect 27433 10081 27445 10115
rect 27479 10112 27491 10115
rect 27614 10112 27620 10124
rect 27479 10084 27620 10112
rect 27479 10081 27491 10084
rect 27433 10075 27491 10081
rect 27614 10072 27620 10084
rect 27672 10072 27678 10124
rect 27908 10112 27936 10152
rect 27982 10140 27988 10192
rect 28040 10180 28046 10192
rect 28813 10183 28871 10189
rect 28813 10180 28825 10183
rect 28040 10152 28825 10180
rect 28040 10140 28046 10152
rect 28813 10149 28825 10152
rect 28859 10149 28871 10183
rect 29822 10180 29828 10192
rect 28813 10143 28871 10149
rect 28920 10152 29828 10180
rect 28920 10112 28948 10152
rect 29822 10140 29828 10152
rect 29880 10140 29886 10192
rect 29932 10180 29960 10220
rect 31202 10208 31208 10260
rect 31260 10208 31266 10260
rect 31662 10208 31668 10260
rect 31720 10248 31726 10260
rect 32858 10248 32864 10260
rect 31720 10220 32864 10248
rect 31720 10208 31726 10220
rect 32858 10208 32864 10220
rect 32916 10208 32922 10260
rect 34422 10208 34428 10260
rect 34480 10208 34486 10260
rect 31294 10180 31300 10192
rect 29932 10152 31300 10180
rect 31294 10140 31300 10152
rect 31352 10140 31358 10192
rect 31570 10140 31576 10192
rect 31628 10180 31634 10192
rect 32585 10183 32643 10189
rect 32585 10180 32597 10183
rect 31628 10152 32597 10180
rect 31628 10140 31634 10152
rect 32585 10149 32597 10152
rect 32631 10149 32643 10183
rect 32585 10143 32643 10149
rect 33505 10183 33563 10189
rect 33505 10149 33517 10183
rect 33551 10180 33563 10183
rect 33870 10180 33876 10192
rect 33551 10152 33876 10180
rect 33551 10149 33563 10152
rect 33505 10143 33563 10149
rect 33870 10140 33876 10152
rect 33928 10140 33934 10192
rect 29178 10112 29184 10124
rect 27908 10084 28948 10112
rect 27522 10004 27528 10056
rect 27580 10004 27586 10056
rect 27706 10004 27712 10056
rect 27764 10044 27770 10056
rect 27985 10047 28043 10053
rect 27985 10044 27997 10047
rect 27764 10016 27997 10044
rect 27764 10004 27770 10016
rect 27985 10013 27997 10016
rect 28031 10013 28043 10047
rect 27985 10007 28043 10013
rect 28074 10004 28080 10056
rect 28132 10004 28138 10056
rect 28350 10004 28356 10056
rect 28408 10004 28414 10056
rect 28442 10004 28448 10056
rect 28500 10004 28506 10056
rect 28629 10047 28687 10053
rect 28629 10013 28641 10047
rect 28675 10044 28687 10047
rect 28718 10044 28724 10056
rect 28675 10016 28724 10044
rect 28675 10013 28687 10016
rect 28629 10007 28687 10013
rect 28718 10004 28724 10016
rect 28776 10004 28782 10056
rect 28920 10053 28948 10084
rect 29012 10084 29184 10112
rect 29012 10053 29040 10084
rect 29178 10072 29184 10084
rect 29236 10072 29242 10124
rect 29270 10072 29276 10124
rect 29328 10112 29334 10124
rect 29733 10115 29791 10121
rect 29733 10112 29745 10115
rect 29328 10084 29745 10112
rect 29328 10072 29334 10084
rect 29733 10081 29745 10084
rect 29779 10081 29791 10115
rect 29733 10075 29791 10081
rect 28905 10047 28963 10053
rect 28905 10013 28917 10047
rect 28951 10013 28963 10047
rect 28905 10007 28963 10013
rect 28997 10047 29055 10053
rect 28997 10013 29009 10047
rect 29043 10013 29055 10047
rect 28997 10007 29055 10013
rect 29086 10004 29092 10056
rect 29144 10044 29150 10056
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 29144 10016 29561 10044
rect 29144 10004 29150 10016
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29840 10044 29868 10140
rect 30190 10072 30196 10124
rect 30248 10112 30254 10124
rect 30248 10084 30604 10112
rect 30248 10072 30254 10084
rect 30576 10053 30604 10084
rect 31386 10072 31392 10124
rect 31444 10072 31450 10124
rect 31938 10112 31944 10124
rect 31496 10084 31944 10112
rect 30285 10047 30343 10053
rect 30285 10044 30297 10047
rect 29840 10016 30297 10044
rect 29549 10007 29607 10013
rect 30285 10013 30297 10016
rect 30331 10013 30343 10047
rect 30285 10007 30343 10013
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10013 30619 10047
rect 30561 10007 30619 10013
rect 31018 10004 31024 10056
rect 31076 10004 31082 10056
rect 31205 10047 31263 10053
rect 31205 10013 31217 10047
rect 31251 10013 31263 10047
rect 31496 10044 31524 10084
rect 31938 10072 31944 10084
rect 31996 10072 32002 10124
rect 32398 10072 32404 10124
rect 32456 10112 32462 10124
rect 34977 10115 35035 10121
rect 34977 10112 34989 10115
rect 32456 10084 34989 10112
rect 32456 10072 32462 10084
rect 31205 10007 31263 10013
rect 31312 10016 31524 10044
rect 31665 10047 31723 10053
rect 26568 9948 27200 9976
rect 27617 9979 27675 9985
rect 26568 9936 26574 9948
rect 27617 9945 27629 9979
rect 27663 9976 27675 9979
rect 27663 9948 28764 9976
rect 27663 9945 27675 9948
rect 27617 9939 27675 9945
rect 24320 9880 25820 9908
rect 23201 9871 23259 9877
rect 27798 9868 27804 9920
rect 27856 9868 27862 9920
rect 28537 9911 28595 9917
rect 28537 9877 28549 9911
rect 28583 9908 28595 9911
rect 28626 9908 28632 9920
rect 28583 9880 28632 9908
rect 28583 9877 28595 9880
rect 28537 9871 28595 9877
rect 28626 9868 28632 9880
rect 28684 9868 28690 9920
rect 28736 9908 28764 9948
rect 28810 9936 28816 9988
rect 28868 9976 28874 9988
rect 30101 9979 30159 9985
rect 30101 9976 30113 9979
rect 28868 9948 30113 9976
rect 28868 9936 28874 9948
rect 30101 9945 30113 9948
rect 30147 9945 30159 9979
rect 30101 9939 30159 9945
rect 30466 9936 30472 9988
rect 30524 9976 30530 9988
rect 31220 9976 31248 10007
rect 30524 9948 31248 9976
rect 30524 9936 30530 9948
rect 28902 9908 28908 9920
rect 28736 9880 28908 9908
rect 28902 9868 28908 9880
rect 28960 9908 28966 9920
rect 29181 9911 29239 9917
rect 29181 9908 29193 9911
rect 28960 9880 29193 9908
rect 28960 9868 28966 9880
rect 29181 9877 29193 9880
rect 29227 9877 29239 9911
rect 29181 9871 29239 9877
rect 29730 9868 29736 9920
rect 29788 9908 29794 9920
rect 30193 9911 30251 9917
rect 30193 9908 30205 9911
rect 29788 9880 30205 9908
rect 29788 9868 29794 9880
rect 30193 9877 30205 9880
rect 30239 9877 30251 9911
rect 30193 9871 30251 9877
rect 30282 9868 30288 9920
rect 30340 9908 30346 9920
rect 30653 9911 30711 9917
rect 30653 9908 30665 9911
rect 30340 9880 30665 9908
rect 30340 9868 30346 9880
rect 30653 9877 30665 9880
rect 30699 9908 30711 9911
rect 31312 9908 31340 10016
rect 31665 10013 31677 10047
rect 31711 10044 31723 10047
rect 31754 10044 31760 10056
rect 31711 10016 31760 10044
rect 31711 10013 31723 10016
rect 31665 10007 31723 10013
rect 31754 10004 31760 10016
rect 31812 10044 31818 10056
rect 32122 10044 32128 10056
rect 31812 10016 32128 10044
rect 31812 10004 31818 10016
rect 32122 10004 32128 10016
rect 32180 10004 32186 10056
rect 32766 10004 32772 10056
rect 32824 10044 32830 10056
rect 33704 10053 33732 10084
rect 34977 10081 34989 10084
rect 35023 10081 35035 10115
rect 34977 10075 35035 10081
rect 35434 10072 35440 10124
rect 35492 10072 35498 10124
rect 33689 10047 33747 10053
rect 32824 10016 33456 10044
rect 32824 10004 32830 10016
rect 32401 9979 32459 9985
rect 32401 9945 32413 9979
rect 32447 9976 32459 9979
rect 32490 9976 32496 9988
rect 32447 9948 32496 9976
rect 32447 9945 32459 9948
rect 32401 9939 32459 9945
rect 32490 9936 32496 9948
rect 32548 9976 32554 9988
rect 33318 9976 33324 9988
rect 32548 9948 33324 9976
rect 32548 9936 32554 9948
rect 33318 9936 33324 9948
rect 33376 9936 33382 9988
rect 33428 9976 33456 10016
rect 33689 10013 33701 10047
rect 33735 10013 33747 10047
rect 33689 10007 33747 10013
rect 33781 10047 33839 10053
rect 33781 10013 33793 10047
rect 33827 10044 33839 10047
rect 33870 10044 33876 10056
rect 33827 10016 33876 10044
rect 33827 10013 33839 10016
rect 33781 10007 33839 10013
rect 33870 10004 33876 10016
rect 33928 10004 33934 10056
rect 34698 10004 34704 10056
rect 34756 10004 34762 10056
rect 34057 9979 34115 9985
rect 34057 9976 34069 9979
rect 33428 9948 34069 9976
rect 34057 9945 34069 9948
rect 34103 9945 34115 9979
rect 34057 9939 34115 9945
rect 34241 9979 34299 9985
rect 34241 9945 34253 9979
rect 34287 9976 34299 9979
rect 34790 9976 34796 9988
rect 34287 9948 34796 9976
rect 34287 9945 34299 9948
rect 34241 9939 34299 9945
rect 34790 9936 34796 9948
rect 34848 9936 34854 9988
rect 35158 9936 35164 9988
rect 35216 9976 35222 9988
rect 35452 9976 35480 10072
rect 35621 9979 35679 9985
rect 35621 9976 35633 9979
rect 35216 9948 35633 9976
rect 35216 9936 35222 9948
rect 35621 9945 35633 9948
rect 35667 9945 35679 9979
rect 35621 9939 35679 9945
rect 35986 9936 35992 9988
rect 36044 9936 36050 9988
rect 30699 9880 31340 9908
rect 30699 9877 30711 9880
rect 30653 9871 30711 9877
rect 31386 9868 31392 9920
rect 31444 9908 31450 9920
rect 33134 9908 33140 9920
rect 31444 9880 33140 9908
rect 31444 9868 31450 9880
rect 33134 9868 33140 9880
rect 33192 9868 33198 9920
rect 34146 9868 34152 9920
rect 34204 9908 34210 9920
rect 34330 9908 34336 9920
rect 34204 9880 34336 9908
rect 34204 9868 34210 9880
rect 34330 9868 34336 9880
rect 34388 9868 34394 9920
rect 1104 9818 36432 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 36432 9818
rect 1104 9744 36432 9766
rect 3145 9707 3203 9713
rect 3145 9673 3157 9707
rect 3191 9704 3203 9707
rect 3418 9704 3424 9716
rect 3191 9676 3424 9704
rect 3191 9673 3203 9676
rect 3145 9667 3203 9673
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 5445 9707 5503 9713
rect 3896 9676 4752 9704
rect 2314 9596 2320 9648
rect 2372 9596 2378 9648
rect 2682 9596 2688 9648
rect 2740 9596 2746 9648
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2464 9540 2513 9568
rect 2464 9528 2470 9540
rect 2501 9537 2513 9540
rect 2547 9568 2559 9571
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2547 9540 2973 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2961 9537 2973 9540
rect 3007 9568 3019 9571
rect 3896 9568 3924 9676
rect 4614 9636 4620 9648
rect 3988 9608 4620 9636
rect 3988 9577 4016 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 4724 9636 4752 9676
rect 5445 9673 5457 9707
rect 5491 9704 5503 9707
rect 5626 9704 5632 9716
rect 5491 9676 5632 9704
rect 5491 9673 5503 9676
rect 5445 9667 5503 9673
rect 5626 9664 5632 9676
rect 5684 9664 5690 9716
rect 6932 9676 7604 9704
rect 6932 9636 6960 9676
rect 4724 9608 6960 9636
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7466 9636 7472 9648
rect 7055 9608 7472 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 7576 9636 7604 9676
rect 8478 9664 8484 9716
rect 8536 9704 8542 9716
rect 8754 9704 8760 9716
rect 8536 9676 8760 9704
rect 8536 9664 8542 9676
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 8941 9707 8999 9713
rect 8941 9673 8953 9707
rect 8987 9704 8999 9707
rect 9306 9704 9312 9716
rect 8987 9676 9312 9704
rect 8987 9673 8999 9676
rect 8941 9667 8999 9673
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 10870 9704 10876 9716
rect 9692 9676 10876 9704
rect 7742 9636 7748 9648
rect 7576 9608 7748 9636
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 9692 9636 9720 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13265 9707 13323 9713
rect 13265 9704 13277 9707
rect 12768 9676 13277 9704
rect 12768 9664 12774 9676
rect 11974 9636 11980 9648
rect 8404 9608 8800 9636
rect 3007 9540 3924 9568
rect 3973 9571 4031 9577
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4157 9571 4215 9577
rect 4157 9568 4169 9571
rect 4120 9540 4169 9568
rect 4120 9528 4126 9540
rect 4157 9537 4169 9540
rect 4203 9568 4215 9571
rect 4203 9540 4384 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 3050 9500 3056 9512
rect 2823 9472 3056 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 3050 9460 3056 9472
rect 3108 9460 3114 9512
rect 4356 9500 4384 9540
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5258 9568 5264 9580
rect 5215 9540 5264 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5442 9568 5448 9580
rect 5403 9540 5448 9568
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5552 9540 6009 9568
rect 5077 9503 5135 9509
rect 5077 9500 5089 9503
rect 4356 9472 5089 9500
rect 5077 9469 5089 9472
rect 5123 9500 5135 9503
rect 5552 9500 5580 9540
rect 5997 9537 6009 9540
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 5123 9472 5580 9500
rect 5905 9503 5963 9509
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5905 9469 5917 9503
rect 5951 9500 5963 9503
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 5951 9472 6101 9500
rect 5951 9469 5963 9472
rect 5905 9463 5963 9469
rect 6089 9469 6101 9472
rect 6135 9469 6147 9503
rect 6196 9500 6224 9531
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 6914 9577 6920 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6912 9568 6920 9577
rect 6875 9540 6920 9568
rect 6549 9531 6607 9537
rect 6912 9531 6920 9540
rect 6564 9500 6592 9531
rect 6914 9528 6920 9531
rect 6972 9528 6978 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 7024 9540 7113 9568
rect 7024 9512 7052 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 7284 9571 7342 9577
rect 7284 9537 7296 9571
rect 7330 9537 7342 9571
rect 7284 9531 7342 9537
rect 6196 9472 6592 9500
rect 6089 9463 6147 9469
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 4890 9432 4896 9444
rect 4028 9404 4896 9432
rect 4028 9392 4034 9404
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 6564 9432 6592 9472
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 7300 9500 7328 9531
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7650 9528 7656 9580
rect 7708 9528 7714 9580
rect 7834 9528 7840 9580
rect 7892 9528 7898 9580
rect 8202 9528 8208 9580
rect 8260 9528 8266 9580
rect 8404 9577 8432 9608
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8665 9571 8723 9577
rect 8665 9568 8677 9571
rect 8389 9531 8447 9537
rect 8496 9540 8677 9568
rect 7466 9500 7472 9512
rect 7300 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 8018 9460 8024 9512
rect 8076 9460 8082 9512
rect 8202 9432 8208 9444
rect 6564 9404 8208 9432
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 4065 9367 4123 9373
rect 4065 9333 4077 9367
rect 4111 9364 4123 9367
rect 4798 9364 4804 9376
rect 4111 9336 4804 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 5166 9324 5172 9376
rect 5224 9364 5230 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 5224 9336 5273 9364
rect 5224 9324 5230 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 5261 9327 5319 9333
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 5902 9364 5908 9376
rect 5859 9336 5908 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6549 9367 6607 9373
rect 6549 9333 6561 9367
rect 6595 9364 6607 9367
rect 6638 9364 6644 9376
rect 6595 9336 6644 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 6730 9324 6736 9376
rect 6788 9324 6794 9376
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8496 9364 8524 9540
rect 8665 9537 8677 9540
rect 8711 9537 8723 9571
rect 8665 9531 8723 9537
rect 8772 9500 8800 9608
rect 9416 9608 9720 9636
rect 10704 9608 11980 9636
rect 8846 9528 8852 9580
rect 8904 9528 8910 9580
rect 9030 9528 9036 9580
rect 9088 9568 9094 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 9088 9540 9137 9568
rect 9088 9528 9094 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9214 9528 9220 9580
rect 9272 9528 9278 9580
rect 9416 9577 9444 9608
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 9858 9568 9864 9580
rect 9539 9540 9864 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10410 9528 10416 9580
rect 10468 9528 10474 9580
rect 10704 9577 10732 9608
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 12820 9645 12848 9676
rect 13265 9673 13277 9676
rect 13311 9704 13323 9707
rect 13354 9704 13360 9716
rect 13311 9676 13360 9704
rect 13311 9673 13323 9676
rect 13265 9667 13323 9673
rect 13354 9664 13360 9676
rect 13412 9704 13418 9716
rect 14642 9704 14648 9716
rect 13412 9676 14648 9704
rect 13412 9664 13418 9676
rect 14642 9664 14648 9676
rect 14700 9704 14706 9716
rect 15010 9704 15016 9716
rect 14700 9676 15016 9704
rect 14700 9664 14706 9676
rect 15010 9664 15016 9676
rect 15068 9664 15074 9716
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 20898 9704 20904 9716
rect 19116 9676 20904 9704
rect 19116 9664 19122 9676
rect 12605 9639 12663 9645
rect 12605 9605 12617 9639
rect 12651 9636 12663 9639
rect 12805 9639 12863 9645
rect 12651 9608 12756 9636
rect 12651 9605 12663 9608
rect 12605 9599 12663 9605
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9568 10931 9571
rect 10962 9568 10968 9580
rect 10919 9540 10968 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 9582 9500 9588 9512
rect 8772 9472 9588 9500
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9500 10379 9503
rect 10594 9500 10600 9512
rect 10367 9472 10600 9500
rect 10367 9469 10379 9472
rect 10321 9463 10379 9469
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10796 9500 10824 9531
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11698 9568 11704 9580
rect 11195 9540 11704 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11072 9500 11100 9531
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 12728 9568 12756 9608
rect 12805 9605 12817 9639
rect 12851 9605 12863 9639
rect 12805 9599 12863 9605
rect 12894 9596 12900 9648
rect 12952 9596 12958 9648
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 13004 9608 13308 9636
rect 13004 9568 13032 9608
rect 12728 9540 13032 9568
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13127 9540 13216 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 10796 9472 11008 9500
rect 11072 9472 11529 9500
rect 8757 9435 8815 9441
rect 8757 9401 8769 9435
rect 8803 9432 8815 9435
rect 9398 9432 9404 9444
rect 8803 9404 9404 9432
rect 8803 9401 8815 9404
rect 8757 9395 8815 9401
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 10870 9432 10876 9444
rect 10428 9404 10876 9432
rect 7800 9336 8524 9364
rect 7800 9324 7806 9336
rect 8570 9324 8576 9376
rect 8628 9324 8634 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 10045 9367 10103 9373
rect 10045 9364 10057 9367
rect 9180 9336 10057 9364
rect 9180 9324 9186 9336
rect 10045 9333 10057 9336
rect 10091 9333 10103 9367
rect 10045 9327 10103 9333
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 10428 9373 10456 9404
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10980 9432 11008 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 11606 9432 11612 9444
rect 10980 9404 11612 9432
rect 11606 9392 11612 9404
rect 11664 9392 11670 9444
rect 11701 9435 11759 9441
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 12526 9432 12532 9444
rect 11747 9404 12532 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 10376 9336 10425 9364
rect 10376 9324 10382 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10413 9327 10471 9333
rect 10502 9324 10508 9376
rect 10560 9324 10566 9376
rect 12434 9324 12440 9376
rect 12492 9324 12498 9376
rect 12621 9367 12679 9373
rect 12621 9333 12633 9367
rect 12667 9364 12679 9367
rect 12710 9364 12716 9376
rect 12667 9336 12716 9364
rect 12667 9333 12679 9336
rect 12621 9327 12679 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 13188 9364 13216 9540
rect 13280 9500 13308 9608
rect 15120 9608 16681 9636
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9568 13415 9571
rect 13446 9568 13452 9580
rect 13403 9540 13452 9568
rect 13403 9537 13415 9540
rect 13357 9531 13415 9537
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9568 13875 9571
rect 13906 9568 13912 9580
rect 13863 9540 13912 9568
rect 13863 9537 13875 9540
rect 13817 9531 13875 9537
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 14734 9528 14740 9580
rect 14792 9528 14798 9580
rect 14826 9528 14832 9580
rect 14884 9568 14890 9580
rect 15120 9568 15148 9608
rect 16669 9605 16681 9608
rect 16715 9605 16727 9639
rect 16669 9599 16727 9605
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17862 9636 17868 9648
rect 17083 9608 17868 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 19352 9645 19380 9676
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 22462 9704 22468 9716
rect 22112 9676 22468 9704
rect 19337 9639 19395 9645
rect 19337 9605 19349 9639
rect 19383 9605 19395 9639
rect 19337 9599 19395 9605
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 19521 9639 19579 9645
rect 19521 9636 19533 9639
rect 19484 9608 19533 9636
rect 19484 9596 19490 9608
rect 19521 9605 19533 9608
rect 19567 9605 19579 9639
rect 19521 9599 19579 9605
rect 14884 9540 15148 9568
rect 14884 9528 14890 9540
rect 15194 9528 15200 9580
rect 15252 9528 15258 9580
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9568 17187 9571
rect 17678 9568 17684 9580
rect 17175 9540 17684 9568
rect 17175 9537 17187 9540
rect 17129 9531 17187 9537
rect 13280 9472 13952 9500
rect 13538 9392 13544 9444
rect 13596 9432 13602 9444
rect 13633 9435 13691 9441
rect 13633 9432 13645 9435
rect 13596 9404 13645 9432
rect 13596 9392 13602 9404
rect 13633 9401 13645 9404
rect 13679 9401 13691 9435
rect 13924 9432 13952 9472
rect 13998 9460 14004 9512
rect 14056 9460 14062 9512
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9500 15071 9503
rect 15562 9500 15568 9512
rect 15059 9472 15568 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 16868 9500 16896 9531
rect 17678 9528 17684 9540
rect 17736 9528 17742 9580
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 19153 9571 19211 9577
rect 19153 9568 19165 9571
rect 18196 9540 19165 9568
rect 18196 9528 18202 9540
rect 19153 9537 19165 9540
rect 19199 9537 19211 9571
rect 19153 9531 19211 9537
rect 20806 9528 20812 9580
rect 20864 9528 20870 9580
rect 20898 9528 20904 9580
rect 20956 9528 20962 9580
rect 20990 9528 20996 9580
rect 21048 9528 21054 9580
rect 22112 9577 22140 9676
rect 22462 9664 22468 9676
rect 22520 9664 22526 9716
rect 22554 9664 22560 9716
rect 22612 9664 22618 9716
rect 23842 9704 23848 9716
rect 22664 9676 23848 9704
rect 22664 9636 22692 9676
rect 23842 9664 23848 9676
rect 23900 9664 23906 9716
rect 26326 9664 26332 9716
rect 26384 9704 26390 9716
rect 27062 9704 27068 9716
rect 26384 9676 27068 9704
rect 26384 9664 26390 9676
rect 27062 9664 27068 9676
rect 27120 9664 27126 9716
rect 28442 9704 28448 9716
rect 27172 9676 28448 9704
rect 22388 9608 22692 9636
rect 22725 9639 22783 9645
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 22077 9571 22140 9577
rect 22077 9537 22089 9571
rect 22123 9540 22140 9571
rect 22123 9537 22135 9540
rect 22077 9531 22135 9537
rect 18046 9500 18052 9512
rect 16868 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 19886 9460 19892 9512
rect 19944 9500 19950 9512
rect 21192 9500 21220 9531
rect 22186 9528 22192 9580
rect 22244 9528 22250 9580
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9558 22339 9571
rect 22388 9558 22416 9608
rect 22725 9605 22737 9639
rect 22771 9636 22783 9639
rect 22925 9639 22983 9645
rect 22771 9608 22876 9636
rect 22771 9605 22783 9608
rect 22725 9599 22783 9605
rect 22327 9537 22416 9558
rect 22281 9531 22416 9537
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9568 22600 9571
rect 22848 9568 22876 9608
rect 22925 9605 22937 9639
rect 22971 9636 22983 9639
rect 23014 9636 23020 9648
rect 22971 9608 23020 9636
rect 22971 9605 22983 9608
rect 22925 9599 22983 9605
rect 23014 9596 23020 9608
rect 23072 9596 23078 9648
rect 25222 9596 25228 9648
rect 25280 9636 25286 9648
rect 26344 9636 26372 9664
rect 25280 9608 25728 9636
rect 25280 9596 25286 9608
rect 23382 9568 23388 9580
rect 22511 9543 22784 9568
rect 22511 9537 22523 9543
rect 22572 9540 22784 9543
rect 22848 9540 23388 9568
rect 22465 9531 22523 9537
rect 22296 9530 22416 9531
rect 19944 9472 22324 9500
rect 19944 9460 19950 9472
rect 22296 9444 22324 9472
rect 20625 9435 20683 9441
rect 20625 9432 20637 9435
rect 13924 9404 20637 9432
rect 13633 9395 13691 9401
rect 20625 9401 20637 9404
rect 20671 9401 20683 9435
rect 20625 9395 20683 9401
rect 20898 9392 20904 9444
rect 20956 9432 20962 9444
rect 20956 9404 21956 9432
rect 20956 9392 20962 9404
rect 14093 9367 14151 9373
rect 14093 9364 14105 9367
rect 13188 9336 14105 9364
rect 14093 9333 14105 9336
rect 14139 9364 14151 9367
rect 14182 9364 14188 9376
rect 14139 9336 14188 9364
rect 14139 9333 14151 9336
rect 14093 9327 14151 9333
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 14458 9324 14464 9376
rect 14516 9324 14522 9376
rect 14921 9367 14979 9373
rect 14921 9333 14933 9367
rect 14967 9364 14979 9367
rect 15194 9364 15200 9376
rect 14967 9336 15200 9364
rect 14967 9333 14979 9336
rect 14921 9327 14979 9333
rect 15194 9324 15200 9336
rect 15252 9364 15258 9376
rect 15838 9364 15844 9376
rect 15252 9336 15844 9364
rect 15252 9324 15258 9336
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 18046 9324 18052 9376
rect 18104 9364 18110 9376
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 18104 9336 21833 9364
rect 18104 9324 18110 9336
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 21928 9364 21956 9404
rect 22278 9392 22284 9444
rect 22336 9392 22342 9444
rect 22756 9373 22784 9540
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 23658 9528 23664 9580
rect 23716 9568 23722 9580
rect 25593 9571 25651 9577
rect 25593 9568 25605 9571
rect 23716 9540 25605 9568
rect 23716 9528 23722 9540
rect 25593 9537 25605 9540
rect 25639 9537 25651 9571
rect 25700 9568 25728 9608
rect 26252 9608 26372 9636
rect 26050 9568 26056 9580
rect 25700 9540 26056 9568
rect 25593 9531 25651 9537
rect 26050 9528 26056 9540
rect 26108 9528 26114 9580
rect 25777 9503 25835 9509
rect 25777 9469 25789 9503
rect 25823 9500 25835 9503
rect 26252 9500 26280 9608
rect 26418 9596 26424 9648
rect 26476 9596 26482 9648
rect 26712 9608 27108 9636
rect 26712 9577 26740 9608
rect 26329 9571 26387 9577
rect 26329 9537 26341 9571
rect 26375 9568 26387 9571
rect 26513 9571 26571 9577
rect 26375 9540 26464 9568
rect 26375 9537 26387 9540
rect 26329 9531 26387 9537
rect 25823 9472 26280 9500
rect 25823 9469 25835 9472
rect 25777 9463 25835 9469
rect 25685 9435 25743 9441
rect 25685 9401 25697 9435
rect 25731 9432 25743 9435
rect 26145 9435 26203 9441
rect 26145 9432 26157 9435
rect 25731 9404 26157 9432
rect 25731 9401 25743 9404
rect 25685 9395 25743 9401
rect 26145 9401 26157 9404
rect 26191 9401 26203 9435
rect 26145 9395 26203 9401
rect 22741 9367 22799 9373
rect 22741 9364 22753 9367
rect 21928 9336 22753 9364
rect 21821 9327 21879 9333
rect 22741 9333 22753 9336
rect 22787 9364 22799 9367
rect 23198 9364 23204 9376
rect 22787 9336 23204 9364
rect 22787 9333 22799 9336
rect 22741 9327 22799 9333
rect 23198 9324 23204 9336
rect 23256 9324 23262 9376
rect 23290 9324 23296 9376
rect 23348 9364 23354 9376
rect 25317 9367 25375 9373
rect 25317 9364 25329 9367
rect 23348 9336 25329 9364
rect 23348 9324 23354 9336
rect 25317 9333 25329 9336
rect 25363 9333 25375 9367
rect 25317 9327 25375 9333
rect 25866 9324 25872 9376
rect 25924 9324 25930 9376
rect 26436 9364 26464 9540
rect 26513 9537 26525 9571
rect 26559 9537 26571 9571
rect 26513 9531 26571 9537
rect 26697 9571 26755 9577
rect 26697 9537 26709 9571
rect 26743 9537 26755 9571
rect 26697 9531 26755 9537
rect 26528 9500 26556 9531
rect 26970 9528 26976 9580
rect 27028 9528 27034 9580
rect 26786 9500 26792 9512
rect 26528 9472 26792 9500
rect 26786 9460 26792 9472
rect 26844 9460 26850 9512
rect 27080 9500 27108 9608
rect 27172 9580 27200 9676
rect 28442 9664 28448 9676
rect 28500 9664 28506 9716
rect 28534 9664 28540 9716
rect 28592 9704 28598 9716
rect 31018 9704 31024 9716
rect 28592 9676 31024 9704
rect 28592 9664 28598 9676
rect 31018 9664 31024 9676
rect 31076 9664 31082 9716
rect 32214 9664 32220 9716
rect 32272 9664 32278 9716
rect 34698 9664 34704 9716
rect 34756 9704 34762 9716
rect 35253 9707 35311 9713
rect 35253 9704 35265 9707
rect 34756 9676 35265 9704
rect 34756 9664 34762 9676
rect 35253 9673 35265 9676
rect 35299 9673 35311 9707
rect 35253 9667 35311 9673
rect 28350 9596 28356 9648
rect 28408 9636 28414 9648
rect 31846 9636 31852 9648
rect 28408 9608 31852 9636
rect 28408 9596 28414 9608
rect 31846 9596 31852 9608
rect 31904 9636 31910 9648
rect 33321 9639 33379 9645
rect 31904 9608 32352 9636
rect 31904 9596 31910 9608
rect 27154 9528 27160 9580
rect 27212 9528 27218 9580
rect 27246 9528 27252 9580
rect 27304 9528 27310 9580
rect 29822 9528 29828 9580
rect 29880 9568 29886 9580
rect 30282 9568 30288 9580
rect 29880 9540 30288 9568
rect 29880 9528 29886 9540
rect 30282 9528 30288 9540
rect 30340 9528 30346 9580
rect 30466 9528 30472 9580
rect 30524 9528 30530 9580
rect 30653 9571 30711 9577
rect 30653 9537 30665 9571
rect 30699 9568 30711 9571
rect 31018 9568 31024 9580
rect 30699 9540 31024 9568
rect 30699 9537 30711 9540
rect 30653 9531 30711 9537
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 31386 9528 31392 9580
rect 31444 9528 31450 9580
rect 31570 9528 31576 9580
rect 31628 9528 31634 9580
rect 32324 9577 32352 9608
rect 33321 9605 33333 9639
rect 33367 9636 33379 9639
rect 33686 9636 33692 9648
rect 33367 9608 33692 9636
rect 33367 9605 33379 9608
rect 33321 9599 33379 9605
rect 33686 9596 33692 9608
rect 33744 9596 33750 9648
rect 33778 9596 33784 9648
rect 33836 9596 33842 9648
rect 34422 9596 34428 9648
rect 34480 9596 34486 9648
rect 35158 9596 35164 9648
rect 35216 9636 35222 9648
rect 35713 9639 35771 9645
rect 35713 9636 35725 9639
rect 35216 9608 35725 9636
rect 35216 9596 35222 9608
rect 35713 9605 35725 9608
rect 35759 9605 35771 9639
rect 35713 9599 35771 9605
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 27522 9500 27528 9512
rect 27080 9472 27528 9500
rect 27522 9460 27528 9472
rect 27580 9500 27586 9512
rect 28166 9500 28172 9512
rect 27580 9472 28172 9500
rect 27580 9460 27586 9472
rect 28166 9460 28172 9472
rect 28224 9460 28230 9512
rect 29546 9460 29552 9512
rect 29604 9500 29610 9512
rect 29641 9503 29699 9509
rect 29641 9500 29653 9503
rect 29604 9472 29653 9500
rect 29604 9460 29610 9472
rect 29641 9469 29653 9472
rect 29687 9469 29699 9503
rect 31754 9500 31760 9512
rect 29641 9463 29699 9469
rect 31036 9472 31760 9500
rect 26973 9435 27031 9441
rect 26973 9401 26985 9435
rect 27019 9432 27031 9435
rect 27062 9432 27068 9444
rect 27019 9404 27068 9432
rect 27019 9401 27031 9404
rect 26973 9395 27031 9401
rect 27062 9392 27068 9404
rect 27120 9392 27126 9444
rect 27614 9392 27620 9444
rect 27672 9432 27678 9444
rect 30009 9435 30067 9441
rect 30009 9432 30021 9435
rect 27672 9404 30021 9432
rect 27672 9392 27678 9404
rect 30009 9401 30021 9404
rect 30055 9401 30067 9435
rect 30009 9395 30067 9401
rect 30377 9435 30435 9441
rect 30377 9401 30389 9435
rect 30423 9432 30435 9435
rect 30926 9432 30932 9444
rect 30423 9404 30932 9432
rect 30423 9401 30435 9404
rect 30377 9395 30435 9401
rect 30926 9392 30932 9404
rect 30984 9392 30990 9444
rect 27338 9364 27344 9376
rect 26436 9336 27344 9364
rect 27338 9324 27344 9336
rect 27396 9364 27402 9376
rect 31036 9364 31064 9472
rect 31754 9460 31760 9472
rect 31812 9460 31818 9512
rect 32324 9500 32352 9531
rect 32398 9528 32404 9580
rect 32456 9528 32462 9580
rect 33042 9528 33048 9580
rect 33100 9568 33106 9580
rect 33229 9571 33287 9577
rect 33229 9568 33241 9571
rect 33100 9540 33241 9568
rect 33100 9528 33106 9540
rect 33229 9537 33241 9540
rect 33275 9537 33287 9571
rect 33229 9531 33287 9537
rect 33413 9571 33471 9577
rect 33413 9537 33425 9571
rect 33459 9537 33471 9571
rect 33413 9531 33471 9537
rect 33428 9500 33456 9531
rect 33502 9528 33508 9580
rect 33560 9528 33566 9580
rect 35066 9528 35072 9580
rect 35124 9568 35130 9580
rect 35124 9540 35480 9568
rect 35124 9528 35130 9540
rect 35342 9500 35348 9512
rect 32324 9472 35348 9500
rect 35342 9460 35348 9472
rect 35400 9460 35406 9512
rect 35452 9500 35480 9540
rect 35526 9528 35532 9580
rect 35584 9528 35590 9580
rect 35618 9500 35624 9512
rect 35452 9472 35624 9500
rect 35618 9460 35624 9472
rect 35676 9460 35682 9512
rect 35250 9392 35256 9444
rect 35308 9432 35314 9444
rect 35434 9432 35440 9444
rect 35308 9404 35440 9432
rect 35308 9392 35314 9404
rect 35434 9392 35440 9404
rect 35492 9392 35498 9444
rect 35710 9392 35716 9444
rect 35768 9432 35774 9444
rect 35897 9435 35955 9441
rect 35897 9432 35909 9435
rect 35768 9404 35909 9432
rect 35768 9392 35774 9404
rect 35897 9401 35909 9404
rect 35943 9401 35955 9435
rect 35897 9395 35955 9401
rect 27396 9336 31064 9364
rect 27396 9324 27402 9336
rect 31386 9324 31392 9376
rect 31444 9364 31450 9376
rect 32582 9364 32588 9376
rect 31444 9336 32588 9364
rect 31444 9324 31450 9336
rect 32582 9324 32588 9336
rect 32640 9324 32646 9376
rect 32766 9324 32772 9376
rect 32824 9364 32830 9376
rect 35345 9367 35403 9373
rect 35345 9364 35357 9367
rect 32824 9336 35357 9364
rect 32824 9324 32830 9336
rect 35345 9333 35357 9336
rect 35391 9333 35403 9367
rect 35345 9327 35403 9333
rect 1104 9274 36432 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 36432 9274
rect 1104 9200 36432 9222
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 4338 9160 4344 9172
rect 3651 9132 4344 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 6420 9132 7021 9160
rect 6420 9120 6426 9132
rect 7009 9129 7021 9132
rect 7055 9129 7067 9163
rect 7009 9123 7067 9129
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8352 9132 8677 9160
rect 8352 9120 8358 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 8665 9123 8723 9129
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 10284 9132 10916 9160
rect 10284 9120 10290 9132
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 2556 9064 7604 9092
rect 2556 9052 2562 9064
rect 4706 9024 4712 9036
rect 3344 8996 4712 9024
rect 3344 8965 3372 8996
rect 3804 8965 3832 8996
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 4890 8984 4896 9036
rect 4948 9024 4954 9036
rect 4985 9027 5043 9033
rect 4985 9024 4997 9027
rect 4948 8996 4997 9024
rect 4948 8984 4954 8996
rect 4985 8993 4997 8996
rect 5031 9024 5043 9027
rect 6086 9024 6092 9036
rect 5031 8996 6092 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6270 8984 6276 9036
rect 6328 8984 6334 9036
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 6604 8996 7236 9024
rect 6604 8984 6610 8996
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3513 8891 3571 8897
rect 3513 8857 3525 8891
rect 3559 8857 3571 8891
rect 3620 8888 3648 8919
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 4120 8928 4537 8956
rect 4120 8916 4126 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 5166 8916 5172 8968
rect 5224 8916 5230 8968
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8956 5503 8959
rect 5626 8956 5632 8968
rect 5491 8928 5632 8956
rect 5491 8925 5503 8928
rect 5445 8919 5503 8925
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8956 5779 8959
rect 6181 8959 6239 8965
rect 6181 8956 6193 8959
rect 5767 8928 6193 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 6181 8925 6193 8928
rect 6227 8925 6239 8959
rect 6288 8956 6316 8984
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 6288 8928 6377 8956
rect 6181 8919 6239 8925
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 4080 8888 4108 8916
rect 4341 8891 4399 8897
rect 4341 8888 4353 8891
rect 3620 8860 4108 8888
rect 4172 8860 4353 8888
rect 3513 8851 3571 8857
rect 3528 8820 3556 8851
rect 3881 8823 3939 8829
rect 3881 8820 3893 8823
rect 3528 8792 3893 8820
rect 3881 8789 3893 8792
rect 3927 8820 3939 8823
rect 4172 8820 4200 8860
rect 4341 8857 4353 8860
rect 4387 8888 4399 8891
rect 4614 8888 4620 8900
rect 4387 8860 4620 8888
rect 4387 8857 4399 8860
rect 4341 8851 4399 8857
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 5350 8888 5356 8900
rect 4908 8860 5356 8888
rect 3927 8792 4200 8820
rect 4249 8823 4307 8829
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4522 8820 4528 8832
rect 4295 8792 4528 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4908 8829 4936 8860
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 5994 8888 6000 8900
rect 5592 8860 6000 8888
rect 5592 8848 5598 8860
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 6472 8888 6500 8919
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 7098 8956 7104 8968
rect 6932 8928 7104 8956
rect 6932 8888 6960 8928
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 7208 8965 7236 8996
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 7466 8956 7472 8968
rect 7239 8928 7472 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7576 8956 7604 9064
rect 8754 9052 8760 9104
rect 8812 9092 8818 9104
rect 8812 9064 9352 9092
rect 8812 9052 8818 9064
rect 8570 8984 8576 9036
rect 8628 9024 8634 9036
rect 8628 8996 9168 9024
rect 8628 8984 8634 8996
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7576 8928 7849 8956
rect 7837 8925 7849 8928
rect 7883 8956 7895 8959
rect 8478 8956 8484 8968
rect 7883 8928 8484 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8720 8928 8769 8956
rect 8720 8916 8726 8928
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 8757 8919 8815 8925
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9140 8965 9168 8996
rect 9324 8965 9352 9064
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 9024 9919 9027
rect 10502 9024 10508 9036
rect 9907 8996 10508 9024
rect 9907 8993 9919 8996
rect 9861 8987 9919 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10888 9024 10916 9132
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11333 9163 11391 9169
rect 11333 9160 11345 9163
rect 11020 9132 11345 9160
rect 11020 9120 11026 9132
rect 11333 9129 11345 9132
rect 11379 9129 11391 9163
rect 11333 9123 11391 9129
rect 11698 9120 11704 9172
rect 11756 9120 11762 9172
rect 16390 9120 16396 9172
rect 16448 9120 16454 9172
rect 16853 9163 16911 9169
rect 16853 9129 16865 9163
rect 16899 9160 16911 9163
rect 18325 9163 18383 9169
rect 18325 9160 18337 9163
rect 16899 9132 18337 9160
rect 16899 9129 16911 9132
rect 16853 9123 16911 9129
rect 18325 9129 18337 9132
rect 18371 9129 18383 9163
rect 18325 9123 18383 9129
rect 22554 9120 22560 9172
rect 22612 9160 22618 9172
rect 22922 9160 22928 9172
rect 22612 9132 22928 9160
rect 22612 9120 22618 9132
rect 22922 9120 22928 9132
rect 22980 9160 22986 9172
rect 23382 9160 23388 9172
rect 22980 9132 23388 9160
rect 22980 9120 22986 9132
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 25866 9120 25872 9172
rect 25924 9160 25930 9172
rect 28445 9163 28503 9169
rect 28445 9160 28457 9163
rect 25924 9132 28457 9160
rect 25924 9120 25930 9132
rect 28445 9129 28457 9132
rect 28491 9129 28503 9163
rect 29362 9160 29368 9172
rect 28445 9123 28503 9129
rect 28966 9132 29368 9160
rect 12526 9052 12532 9104
rect 12584 9092 12590 9104
rect 12584 9064 12940 9092
rect 12584 9052 12590 9064
rect 10888 8996 11560 9024
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 11532 8965 11560 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12492 8996 12817 9024
rect 12492 8984 12498 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 9585 8959 9643 8965
rect 9585 8956 9597 8959
rect 9548 8928 9597 8956
rect 9548 8916 9554 8928
rect 9585 8925 9597 8928
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11606 8916 11612 8968
rect 11664 8956 11670 8968
rect 11701 8959 11759 8965
rect 11701 8956 11713 8959
rect 11664 8928 11713 8956
rect 11664 8916 11670 8928
rect 11701 8925 11713 8928
rect 11747 8925 11759 8959
rect 11701 8919 11759 8925
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8956 12771 8959
rect 12912 8956 12940 9064
rect 14182 9052 14188 9104
rect 14240 9092 14246 9104
rect 16574 9092 16580 9104
rect 14240 9064 16580 9092
rect 14240 9052 14246 9064
rect 16574 9052 16580 9064
rect 16632 9052 16638 9104
rect 17586 9052 17592 9104
rect 17644 9052 17650 9104
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 19058 9092 19064 9104
rect 17828 9064 19064 9092
rect 17828 9052 17834 9064
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 20990 9052 20996 9104
rect 21048 9092 21054 9104
rect 23569 9095 23627 9101
rect 21048 9064 23520 9092
rect 21048 9052 21054 9064
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 9024 16727 9027
rect 17126 9024 17132 9036
rect 16715 8996 17132 9024
rect 16715 8993 16727 8996
rect 16669 8987 16727 8993
rect 17126 8984 17132 8996
rect 17184 9024 17190 9036
rect 19334 9024 19340 9036
rect 17184 8996 18092 9024
rect 17184 8984 17190 8996
rect 18064 8968 18092 8996
rect 18616 8996 19340 9024
rect 12759 8928 12940 8956
rect 16945 8959 17003 8965
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 16945 8925 16957 8959
rect 16991 8925 17003 8959
rect 16945 8919 17003 8925
rect 6472 8860 6960 8888
rect 7285 8891 7343 8897
rect 7285 8857 7297 8891
rect 7331 8857 7343 8891
rect 7285 8851 7343 8857
rect 4709 8823 4767 8829
rect 4709 8789 4721 8823
rect 4755 8820 4767 8823
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4755 8792 4905 8820
rect 4755 8789 4767 8792
rect 4709 8783 4767 8789
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 4893 8783 4951 8789
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5077 8823 5135 8829
rect 5077 8820 5089 8823
rect 5040 8792 5089 8820
rect 5040 8780 5046 8792
rect 5077 8789 5089 8792
rect 5123 8789 5135 8823
rect 5077 8783 5135 8789
rect 5258 8780 5264 8832
rect 5316 8780 5322 8832
rect 5629 8823 5687 8829
rect 5629 8789 5641 8823
rect 5675 8820 5687 8823
rect 6362 8820 6368 8832
rect 5675 8792 6368 8820
rect 5675 8789 5687 8792
rect 5629 8783 5687 8789
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 7300 8820 7328 8851
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 9217 8891 9275 8897
rect 9217 8888 9229 8891
rect 8168 8860 9229 8888
rect 8168 8848 8174 8860
rect 9217 8857 9229 8860
rect 9263 8857 9275 8891
rect 11146 8888 11152 8900
rect 11086 8860 11152 8888
rect 9217 8851 9275 8857
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 6604 8792 7328 8820
rect 7653 8823 7711 8829
rect 6604 8780 6610 8792
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 8754 8820 8760 8832
rect 7699 8792 8760 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 9493 8823 9551 8829
rect 9493 8820 9505 8823
rect 9364 8792 9505 8820
rect 9364 8780 9370 8792
rect 9493 8789 9505 8792
rect 9539 8789 9551 8823
rect 9493 8783 9551 8789
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 10226 8820 10232 8832
rect 10100 8792 10232 8820
rect 10100 8780 10106 8792
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 12032 8792 12265 8820
rect 12032 8780 12038 8792
rect 12253 8789 12265 8792
rect 12299 8789 12311 8823
rect 12253 8783 12311 8789
rect 12618 8780 12624 8832
rect 12676 8780 12682 8832
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 16960 8820 16988 8919
rect 17034 8916 17040 8968
rect 17092 8916 17098 8968
rect 17770 8916 17776 8968
rect 17828 8916 17834 8968
rect 17862 8916 17868 8968
rect 17920 8916 17926 8968
rect 18046 8916 18052 8968
rect 18104 8916 18110 8968
rect 18138 8916 18144 8968
rect 18196 8916 18202 8968
rect 18616 8965 18644 8996
rect 19334 8984 19340 8996
rect 19392 9024 19398 9036
rect 19702 9024 19708 9036
rect 19392 8996 19708 9024
rect 19392 8984 19398 8996
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 20070 8984 20076 9036
rect 20128 8984 20134 9036
rect 20254 8984 20260 9036
rect 20312 8984 20318 9036
rect 23106 9024 23112 9036
rect 20364 8996 23112 9024
rect 18581 8959 18644 8965
rect 18581 8925 18593 8959
rect 18627 8928 18644 8959
rect 18693 8959 18751 8965
rect 18627 8925 18639 8928
rect 18581 8919 18639 8925
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 17405 8891 17463 8897
rect 17405 8857 17417 8891
rect 17451 8888 17463 8891
rect 18230 8888 18236 8900
rect 17451 8860 18236 8888
rect 17451 8857 17463 8860
rect 17405 8851 17463 8857
rect 18230 8848 18236 8860
rect 18288 8848 18294 8900
rect 18708 8888 18736 8919
rect 18782 8916 18788 8968
rect 18840 8916 18846 8968
rect 18966 8916 18972 8968
rect 19024 8916 19030 8968
rect 20364 8956 20392 8996
rect 23106 8984 23112 8996
rect 23164 8984 23170 9036
rect 23492 9024 23520 9064
rect 23569 9061 23581 9095
rect 23615 9092 23627 9095
rect 25038 9092 25044 9104
rect 23615 9064 25044 9092
rect 23615 9061 23627 9064
rect 23569 9055 23627 9061
rect 25038 9052 25044 9064
rect 25096 9052 25102 9104
rect 27341 9095 27399 9101
rect 27341 9061 27353 9095
rect 27387 9092 27399 9095
rect 28350 9092 28356 9104
rect 27387 9064 28356 9092
rect 27387 9061 27399 9064
rect 27341 9055 27399 9061
rect 28350 9052 28356 9064
rect 28408 9052 28414 9104
rect 27798 9024 27804 9036
rect 23492 8996 27804 9024
rect 27798 8984 27804 8996
rect 27856 8984 27862 9036
rect 28966 9024 28994 9132
rect 29362 9120 29368 9132
rect 29420 9120 29426 9172
rect 30742 9120 30748 9172
rect 30800 9120 30806 9172
rect 31389 9163 31447 9169
rect 31389 9129 31401 9163
rect 31435 9160 31447 9163
rect 31478 9160 31484 9172
rect 31435 9132 31484 9160
rect 31435 9129 31447 9132
rect 31389 9123 31447 9129
rect 31478 9120 31484 9132
rect 31536 9120 31542 9172
rect 32674 9120 32680 9172
rect 32732 9160 32738 9172
rect 32861 9163 32919 9169
rect 32861 9160 32873 9163
rect 32732 9132 32873 9160
rect 32732 9120 32738 9132
rect 32861 9129 32873 9132
rect 32907 9129 32919 9163
rect 36354 9160 36360 9172
rect 32861 9123 32919 9129
rect 32968 9132 36360 9160
rect 29086 9052 29092 9104
rect 29144 9092 29150 9104
rect 30466 9092 30472 9104
rect 29144 9064 30472 9092
rect 29144 9052 29150 9064
rect 30466 9052 30472 9064
rect 30524 9052 30530 9104
rect 30929 9095 30987 9101
rect 30929 9061 30941 9095
rect 30975 9061 30987 9095
rect 30929 9055 30987 9061
rect 28460 8996 28994 9024
rect 30944 9024 30972 9055
rect 31938 9052 31944 9104
rect 31996 9092 32002 9104
rect 32968 9092 32996 9132
rect 36354 9120 36360 9132
rect 36412 9120 36418 9172
rect 31996 9064 32996 9092
rect 34057 9095 34115 9101
rect 31996 9052 32002 9064
rect 34057 9061 34069 9095
rect 34103 9061 34115 9095
rect 34057 9055 34115 9061
rect 31757 9027 31815 9033
rect 31757 9024 31769 9027
rect 30944 8996 31769 9024
rect 20180 8928 20392 8956
rect 20441 8959 20499 8965
rect 18524 8860 18736 8888
rect 18524 8832 18552 8860
rect 19242 8848 19248 8900
rect 19300 8888 19306 8900
rect 20180 8888 20208 8928
rect 20441 8925 20453 8959
rect 20487 8925 20499 8959
rect 20441 8919 20499 8925
rect 19300 8860 20208 8888
rect 19300 8848 19306 8860
rect 20346 8848 20352 8900
rect 20404 8888 20410 8900
rect 20456 8888 20484 8919
rect 20530 8916 20536 8968
rect 20588 8956 20594 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20588 8928 20637 8956
rect 20588 8916 20594 8928
rect 20625 8925 20637 8928
rect 20671 8956 20683 8959
rect 23290 8956 23296 8968
rect 20671 8928 23296 8956
rect 20671 8925 20683 8928
rect 20625 8919 20683 8925
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 23382 8916 23388 8968
rect 23440 8916 23446 8968
rect 23477 8959 23535 8965
rect 23477 8925 23489 8959
rect 23523 8925 23535 8959
rect 23477 8919 23535 8925
rect 23201 8891 23259 8897
rect 23201 8888 23213 8891
rect 20404 8860 23213 8888
rect 20404 8848 20410 8860
rect 23201 8857 23213 8860
rect 23247 8857 23259 8891
rect 23201 8851 23259 8857
rect 23492 8888 23520 8919
rect 23658 8916 23664 8968
rect 23716 8916 23722 8968
rect 23768 8928 26832 8956
rect 23566 8888 23572 8900
rect 23492 8860 23572 8888
rect 18322 8820 18328 8832
rect 12860 8792 18328 8820
rect 12860 8780 12866 8792
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 18506 8780 18512 8832
rect 18564 8780 18570 8832
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 23106 8820 23112 8832
rect 19116 8792 23112 8820
rect 19116 8780 19122 8792
rect 23106 8780 23112 8792
rect 23164 8780 23170 8832
rect 23290 8780 23296 8832
rect 23348 8820 23354 8832
rect 23492 8820 23520 8860
rect 23566 8848 23572 8860
rect 23624 8888 23630 8900
rect 23768 8888 23796 8928
rect 23624 8860 23796 8888
rect 23624 8848 23630 8860
rect 26694 8848 26700 8900
rect 26752 8848 26758 8900
rect 26804 8888 26832 8928
rect 27062 8916 27068 8968
rect 27120 8956 27126 8968
rect 27157 8959 27215 8965
rect 27157 8956 27169 8959
rect 27120 8928 27169 8956
rect 27120 8916 27126 8928
rect 27157 8925 27169 8928
rect 27203 8925 27215 8959
rect 27157 8919 27215 8925
rect 27338 8916 27344 8968
rect 27396 8956 27402 8968
rect 28460 8965 28488 8996
rect 27433 8959 27491 8965
rect 27433 8956 27445 8959
rect 27396 8928 27445 8956
rect 27396 8916 27402 8928
rect 27433 8925 27445 8928
rect 27479 8925 27491 8959
rect 27433 8919 27491 8925
rect 28445 8959 28503 8965
rect 28445 8925 28457 8959
rect 28491 8925 28503 8959
rect 28721 8959 28779 8965
rect 28721 8956 28733 8959
rect 28445 8919 28503 8925
rect 28552 8928 28733 8956
rect 27614 8888 27620 8900
rect 26804 8860 27620 8888
rect 27614 8848 27620 8860
rect 27672 8848 27678 8900
rect 23348 8792 23520 8820
rect 23348 8780 23354 8792
rect 25314 8780 25320 8832
rect 25372 8820 25378 8832
rect 28552 8820 28580 8928
rect 28721 8925 28733 8928
rect 28767 8956 28779 8959
rect 29086 8956 29092 8968
rect 28767 8928 29092 8956
rect 28767 8925 28779 8928
rect 28721 8919 28779 8925
rect 29086 8916 29092 8928
rect 29144 8916 29150 8968
rect 29181 8959 29239 8965
rect 29181 8925 29193 8959
rect 29227 8925 29239 8959
rect 29181 8919 29239 8925
rect 28629 8891 28687 8897
rect 28629 8857 28641 8891
rect 28675 8888 28687 8891
rect 29196 8888 29224 8919
rect 29362 8916 29368 8968
rect 29420 8956 29426 8968
rect 30101 8959 30159 8965
rect 29420 8928 29960 8956
rect 29420 8916 29426 8928
rect 29822 8888 29828 8900
rect 28675 8860 29828 8888
rect 28675 8857 28687 8860
rect 28629 8851 28687 8857
rect 29822 8848 29828 8860
rect 29880 8848 29886 8900
rect 29932 8832 29960 8928
rect 30101 8925 30113 8959
rect 30147 8956 30159 8959
rect 30944 8956 30972 8996
rect 31757 8993 31769 8996
rect 31803 9024 31815 9027
rect 33781 9027 33839 9033
rect 33781 9024 33793 9027
rect 31803 8996 33793 9024
rect 31803 8993 31815 8996
rect 31757 8987 31815 8993
rect 31864 8965 31892 8996
rect 30147 8928 30972 8956
rect 31573 8959 31631 8965
rect 30147 8925 30159 8928
rect 30101 8919 30159 8925
rect 31573 8925 31585 8959
rect 31619 8925 31631 8959
rect 31573 8919 31631 8925
rect 31849 8959 31907 8965
rect 31849 8925 31861 8959
rect 31895 8925 31907 8959
rect 31849 8919 31907 8925
rect 30285 8891 30343 8897
rect 30285 8857 30297 8891
rect 30331 8888 30343 8891
rect 31205 8891 31263 8897
rect 31205 8888 31217 8891
rect 30331 8860 31217 8888
rect 30331 8857 30343 8860
rect 30285 8851 30343 8857
rect 31205 8857 31217 8860
rect 31251 8888 31263 8891
rect 31588 8888 31616 8919
rect 31938 8916 31944 8968
rect 31996 8956 32002 8968
rect 32309 8959 32367 8965
rect 32309 8956 32321 8959
rect 31996 8928 32321 8956
rect 31996 8916 32002 8928
rect 32309 8925 32321 8928
rect 32355 8956 32367 8959
rect 32398 8956 32404 8968
rect 32355 8928 32404 8956
rect 32355 8925 32367 8928
rect 32309 8919 32367 8925
rect 32398 8916 32404 8928
rect 32456 8916 32462 8968
rect 33060 8965 33088 8996
rect 33781 8993 33793 8996
rect 33827 9024 33839 9027
rect 33962 9024 33968 9036
rect 33827 8996 33968 9024
rect 33827 8993 33839 8996
rect 33781 8987 33839 8993
rect 33962 8984 33968 8996
rect 34020 8984 34026 9036
rect 32493 8959 32551 8965
rect 32493 8925 32505 8959
rect 32539 8956 32551 8959
rect 32861 8959 32919 8965
rect 32861 8956 32873 8959
rect 32539 8928 32873 8956
rect 32539 8925 32551 8928
rect 32493 8919 32551 8925
rect 32861 8925 32873 8928
rect 32907 8925 32919 8959
rect 32861 8919 32919 8925
rect 33045 8959 33103 8965
rect 33045 8925 33057 8959
rect 33091 8925 33103 8959
rect 34072 8956 34100 9055
rect 34238 9052 34244 9104
rect 34296 9052 34302 9104
rect 34422 9052 34428 9104
rect 34480 9092 34486 9104
rect 35710 9092 35716 9104
rect 34480 9064 35716 9092
rect 34480 9052 34486 9064
rect 35710 9052 35716 9064
rect 35768 9052 35774 9104
rect 34606 8984 34612 9036
rect 34664 9024 34670 9036
rect 35066 9024 35072 9036
rect 34664 8996 35072 9024
rect 34664 8984 34670 8996
rect 35066 8984 35072 8996
rect 35124 8984 35130 9036
rect 33045 8919 33103 8925
rect 33980 8928 34100 8956
rect 34885 8959 34943 8965
rect 32030 8888 32036 8900
rect 31251 8860 32036 8888
rect 31251 8857 31263 8860
rect 31205 8851 31263 8857
rect 32030 8848 32036 8860
rect 32088 8888 32094 8900
rect 32508 8888 32536 8919
rect 32088 8860 32536 8888
rect 32876 8888 32904 8919
rect 33980 8888 34008 8928
rect 34885 8925 34897 8959
rect 34931 8925 34943 8959
rect 34885 8919 34943 8925
rect 34146 8888 34152 8900
rect 32876 8860 34152 8888
rect 32088 8848 32094 8860
rect 34146 8848 34152 8860
rect 34204 8848 34210 8900
rect 34238 8848 34244 8900
rect 34296 8888 34302 8900
rect 34900 8888 34928 8919
rect 35158 8916 35164 8968
rect 35216 8956 35222 8968
rect 35253 8959 35311 8965
rect 35253 8956 35265 8959
rect 35216 8928 35265 8956
rect 35216 8916 35222 8928
rect 35253 8925 35265 8928
rect 35299 8956 35311 8959
rect 35434 8956 35440 8968
rect 35299 8928 35440 8956
rect 35299 8925 35311 8928
rect 35253 8919 35311 8925
rect 35434 8916 35440 8928
rect 35492 8916 35498 8968
rect 35618 8888 35624 8900
rect 34296 8860 35624 8888
rect 34296 8848 34302 8860
rect 35618 8848 35624 8860
rect 35676 8848 35682 8900
rect 25372 8792 28580 8820
rect 25372 8780 25378 8792
rect 29086 8780 29092 8832
rect 29144 8820 29150 8832
rect 29454 8820 29460 8832
rect 29144 8792 29460 8820
rect 29144 8780 29150 8792
rect 29454 8780 29460 8792
rect 29512 8780 29518 8832
rect 29914 8780 29920 8832
rect 29972 8820 29978 8832
rect 30009 8823 30067 8829
rect 30009 8820 30021 8823
rect 29972 8792 30021 8820
rect 29972 8780 29978 8792
rect 30009 8789 30021 8792
rect 30055 8789 30067 8823
rect 30009 8783 30067 8789
rect 30098 8780 30104 8832
rect 30156 8820 30162 8832
rect 33226 8820 33232 8832
rect 30156 8792 33232 8820
rect 30156 8780 30162 8792
rect 33226 8780 33232 8792
rect 33284 8780 33290 8832
rect 34330 8780 34336 8832
rect 34388 8820 34394 8832
rect 34882 8820 34888 8832
rect 34388 8792 34888 8820
rect 34388 8780 34394 8792
rect 34882 8780 34888 8792
rect 34940 8820 34946 8832
rect 35069 8823 35127 8829
rect 35069 8820 35081 8823
rect 34940 8792 35081 8820
rect 34940 8780 34946 8792
rect 35069 8789 35081 8792
rect 35115 8789 35127 8823
rect 35069 8783 35127 8789
rect 35437 8823 35495 8829
rect 35437 8789 35449 8823
rect 35483 8820 35495 8823
rect 35526 8820 35532 8832
rect 35483 8792 35532 8820
rect 35483 8789 35495 8792
rect 35437 8783 35495 8789
rect 35526 8780 35532 8792
rect 35584 8780 35590 8832
rect 1104 8730 36432 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 36432 8730
rect 1104 8656 36432 8678
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 4264 8548 4292 8579
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 4614 8616 4620 8628
rect 4396 8588 4620 8616
rect 4396 8576 4402 8588
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 6013 8619 6071 8625
rect 6013 8616 6025 8619
rect 5408 8588 6025 8616
rect 5408 8576 5414 8588
rect 6013 8585 6025 8588
rect 6059 8585 6071 8619
rect 6013 8579 6071 8585
rect 6362 8576 6368 8628
rect 6420 8576 6426 8628
rect 8018 8616 8024 8628
rect 7024 8588 8024 8616
rect 4890 8548 4896 8560
rect 4264 8520 4896 8548
rect 4890 8508 4896 8520
rect 4948 8508 4954 8560
rect 4985 8551 5043 8557
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 5276 8548 5304 8576
rect 5031 8520 5304 8548
rect 5813 8551 5871 8557
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 5813 8517 5825 8551
rect 5859 8548 5871 8551
rect 6270 8548 6276 8560
rect 5859 8520 6276 8548
rect 5859 8517 5871 8520
rect 5813 8511 5871 8517
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 2498 8480 2504 8492
rect 1452 8452 2504 8480
rect 1452 8440 1458 8452
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 4430 8480 4436 8492
rect 3910 8452 4436 8480
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 4522 8440 4528 8492
rect 4580 8480 4586 8492
rect 4801 8483 4859 8489
rect 4580 8452 4752 8480
rect 4580 8440 4586 8452
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8412 2835 8415
rect 4724 8412 4752 8452
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 5074 8480 5080 8492
rect 4847 8452 5080 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5166 8440 5172 8492
rect 5224 8440 5230 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5442 8480 5448 8492
rect 5399 8452 5448 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 4890 8412 4896 8424
rect 2823 8384 4660 8412
rect 4724 8384 4896 8412
rect 2823 8381 2835 8384
rect 2777 8375 2835 8381
rect 4632 8353 4660 8384
rect 4890 8372 4896 8384
rect 4948 8412 4954 8424
rect 5276 8412 5304 8443
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5828 8480 5856 8511
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 5583 8452 5856 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 6546 8440 6552 8492
rect 6604 8480 6610 8492
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 6604 8452 6653 8480
rect 6604 8440 6610 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6788 8452 6929 8480
rect 6788 8440 6794 8452
rect 6917 8449 6929 8452
rect 6963 8480 6975 8483
rect 7024 8480 7052 8588
rect 8018 8576 8024 8588
rect 8076 8616 8082 8628
rect 8662 8616 8668 8628
rect 8076 8588 8668 8616
rect 8076 8576 8082 8588
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 9214 8576 9220 8628
rect 9272 8576 9278 8628
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 10042 8616 10048 8628
rect 9723 8588 10048 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 10042 8576 10048 8588
rect 10100 8616 10106 8628
rect 10410 8616 10416 8628
rect 10100 8588 10416 8616
rect 10100 8576 10106 8588
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 12158 8616 12164 8628
rect 11716 8588 12164 8616
rect 7742 8508 7748 8560
rect 7800 8508 7806 8560
rect 8478 8508 8484 8560
rect 8536 8508 8542 8560
rect 9232 8548 9260 8576
rect 10962 8548 10968 8560
rect 9232 8520 9628 8548
rect 6963 8452 7052 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7098 8440 7104 8492
rect 7156 8440 7162 8492
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8480 7435 8483
rect 7466 8480 7472 8492
rect 7423 8452 7472 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 4948 8384 5304 8412
rect 4948 8372 4954 8384
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6144 8384 6377 8412
rect 6144 8372 6150 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 7576 8412 7604 8443
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 9306 8480 9312 8492
rect 9263 8452 9312 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 7576 8384 7696 8412
rect 6365 8375 6423 8381
rect 4617 8347 4675 8353
rect 4617 8313 4629 8347
rect 4663 8313 4675 8347
rect 4617 8307 4675 8313
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 6181 8347 6239 8353
rect 5500 8316 6040 8344
rect 5500 8304 5506 8316
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 5074 8276 5080 8288
rect 3936 8248 5080 8276
rect 3936 8236 3942 8248
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5721 8279 5779 8285
rect 5721 8245 5733 8279
rect 5767 8276 5779 8279
rect 5902 8276 5908 8288
rect 5767 8248 5908 8276
rect 5767 8245 5779 8248
rect 5721 8239 5779 8245
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 6012 8285 6040 8316
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 6227 8316 6561 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 7006 8344 7012 8356
rect 6871 8316 7012 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 7668 8344 7696 8384
rect 8938 8372 8944 8424
rect 8996 8372 9002 8424
rect 9030 8372 9036 8424
rect 9088 8372 9094 8424
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 9508 8412 9536 8443
rect 9171 8384 9536 8412
rect 9600 8412 9628 8520
rect 9692 8520 10968 8548
rect 9692 8492 9720 8520
rect 9674 8440 9680 8492
rect 9732 8440 9738 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 9600 8384 9781 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 9140 8344 9168 8375
rect 7668 8316 9168 8344
rect 9508 8344 9536 8384
rect 9769 8381 9781 8384
rect 9815 8381 9827 8415
rect 10244 8412 10272 8443
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10428 8489 10456 8520
rect 10962 8508 10968 8520
rect 11020 8508 11026 8560
rect 11348 8548 11376 8576
rect 11164 8520 11376 8548
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 10594 8440 10600 8492
rect 10652 8440 10658 8492
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 10870 8480 10876 8492
rect 10827 8452 10876 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 10870 8440 10876 8452
rect 10928 8480 10934 8492
rect 11164 8489 11192 8520
rect 11716 8492 11744 8588
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 12713 8619 12771 8625
rect 12713 8616 12725 8619
rect 12676 8588 12725 8616
rect 12676 8576 12682 8588
rect 12713 8585 12725 8588
rect 12759 8585 12771 8619
rect 12713 8579 12771 8585
rect 16025 8619 16083 8625
rect 16025 8585 16037 8619
rect 16071 8616 16083 8619
rect 16114 8616 16120 8628
rect 16071 8588 16120 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 18782 8616 18788 8628
rect 18248 8588 18788 8616
rect 12529 8551 12587 8557
rect 11808 8520 12204 8548
rect 11149 8483 11207 8489
rect 10928 8452 11100 8480
rect 10928 8440 10934 8452
rect 10244 8384 10824 8412
rect 9769 8375 9827 8381
rect 10226 8344 10232 8356
rect 9508 8316 10232 8344
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 10796 8288 10824 8384
rect 11072 8344 11100 8452
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 11606 8480 11612 8492
rect 11379 8452 11612 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 11808 8489 11836 8520
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11974 8440 11980 8492
rect 12032 8440 12038 8492
rect 12176 8489 12204 8520
rect 12529 8517 12541 8551
rect 12575 8548 12587 8551
rect 13170 8548 13176 8560
rect 12575 8520 13176 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 16485 8551 16543 8557
rect 16485 8517 16497 8551
rect 16531 8548 16543 8551
rect 18138 8548 18144 8560
rect 16531 8520 18144 8548
rect 16531 8517 16543 8520
rect 16485 8511 16543 8517
rect 18138 8508 18144 8520
rect 18196 8508 18202 8560
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8480 12219 8483
rect 14458 8480 14464 8492
rect 12207 8452 14464 8480
rect 12207 8449 12219 8452
rect 12161 8443 12219 8449
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8412 11299 8415
rect 12084 8412 12112 8443
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8480 16267 8483
rect 16853 8483 16911 8489
rect 16255 8452 16436 8480
rect 16255 8449 16267 8452
rect 16209 8443 16267 8449
rect 11287 8384 12112 8412
rect 16301 8415 16359 8421
rect 11287 8381 11299 8384
rect 11241 8375 11299 8381
rect 16301 8381 16313 8415
rect 16347 8381 16359 8415
rect 16408 8412 16436 8452
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 16666 8412 16672 8424
rect 16408 8384 16672 8412
rect 16301 8375 16359 8381
rect 12802 8344 12808 8356
rect 11072 8316 12808 8344
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 13170 8304 13176 8356
rect 13228 8344 13234 8356
rect 16316 8344 16344 8375
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 16868 8412 16896 8443
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8480 17279 8483
rect 17310 8480 17316 8492
rect 17267 8452 17316 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 17402 8440 17408 8492
rect 17460 8480 17466 8492
rect 17586 8480 17592 8492
rect 17460 8452 17592 8480
rect 17460 8440 17466 8452
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18248 8489 18276 8588
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 19794 8576 19800 8628
rect 19852 8616 19858 8628
rect 20257 8619 20315 8625
rect 20257 8616 20269 8619
rect 19852 8588 20269 8616
rect 19852 8576 19858 8588
rect 20257 8585 20269 8588
rect 20303 8585 20315 8619
rect 20257 8579 20315 8585
rect 21542 8576 21548 8628
rect 21600 8616 21606 8628
rect 23201 8619 23259 8625
rect 23201 8616 23213 8619
rect 21600 8588 23213 8616
rect 21600 8576 21606 8588
rect 23201 8585 23213 8588
rect 23247 8585 23259 8619
rect 23201 8579 23259 8585
rect 23474 8576 23480 8628
rect 23532 8616 23538 8628
rect 23750 8616 23756 8628
rect 23532 8588 23756 8616
rect 23532 8576 23538 8588
rect 23750 8576 23756 8588
rect 23808 8576 23814 8628
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 25317 8619 25375 8625
rect 25317 8616 25329 8619
rect 24820 8588 25329 8616
rect 24820 8576 24826 8588
rect 25317 8585 25329 8588
rect 25363 8585 25375 8619
rect 25317 8579 25375 8585
rect 25406 8576 25412 8628
rect 25464 8616 25470 8628
rect 26602 8616 26608 8628
rect 25464 8588 26608 8616
rect 25464 8576 25470 8588
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 33042 8616 33048 8628
rect 30944 8588 33048 8616
rect 30944 8560 30972 8588
rect 33042 8576 33048 8588
rect 33100 8576 33106 8628
rect 33502 8576 33508 8628
rect 33560 8616 33566 8628
rect 36078 8616 36084 8628
rect 33560 8588 36084 8616
rect 33560 8576 33566 8588
rect 36078 8576 36084 8588
rect 36136 8576 36142 8628
rect 18322 8508 18328 8560
rect 18380 8508 18386 8560
rect 18506 8508 18512 8560
rect 18564 8548 18570 8560
rect 29086 8548 29092 8560
rect 18564 8520 29092 8548
rect 18564 8508 18570 8520
rect 18616 8489 18644 8520
rect 29086 8508 29092 8520
rect 29144 8508 29150 8560
rect 30009 8551 30067 8557
rect 30009 8548 30021 8551
rect 29196 8520 30021 8548
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 18012 8452 18245 8480
rect 18012 8440 18018 8452
rect 18233 8449 18245 8452
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 19058 8440 19064 8492
rect 19116 8480 19122 8492
rect 20254 8480 20260 8492
rect 19116 8452 20260 8480
rect 19116 8440 19122 8452
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 20530 8440 20536 8492
rect 20588 8440 20594 8492
rect 20622 8440 20628 8492
rect 20680 8440 20686 8492
rect 23290 8480 23296 8492
rect 22066 8452 23296 8480
rect 17034 8412 17040 8424
rect 16868 8384 17040 8412
rect 17034 8372 17040 8384
rect 17092 8372 17098 8424
rect 18785 8415 18843 8421
rect 18785 8381 18797 8415
rect 18831 8381 18843 8415
rect 18785 8375 18843 8381
rect 16758 8344 16764 8356
rect 13228 8316 14412 8344
rect 16316 8316 16764 8344
rect 13228 8304 13234 8316
rect 5997 8279 6055 8285
rect 5997 8245 6009 8279
rect 6043 8245 6055 8279
rect 5997 8239 6055 8245
rect 7190 8236 7196 8288
rect 7248 8236 7254 8288
rect 8757 8279 8815 8285
rect 8757 8245 8769 8279
rect 8803 8276 8815 8279
rect 8846 8276 8852 8288
rect 8803 8248 8852 8276
rect 8803 8245 8815 8248
rect 8757 8239 8815 8245
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 10778 8236 10784 8288
rect 10836 8236 10842 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 11517 8279 11575 8285
rect 11517 8276 11529 8279
rect 11480 8248 11529 8276
rect 11480 8236 11486 8248
rect 11517 8245 11529 8248
rect 11563 8245 11575 8279
rect 11517 8239 11575 8245
rect 11606 8236 11612 8288
rect 11664 8276 11670 8288
rect 11882 8276 11888 8288
rect 11664 8248 11888 8276
rect 11664 8236 11670 8248
rect 11882 8236 11888 8248
rect 11940 8276 11946 8288
rect 12529 8279 12587 8285
rect 12529 8276 12541 8279
rect 11940 8248 12541 8276
rect 11940 8236 11946 8248
rect 12529 8245 12541 8248
rect 12575 8276 12587 8279
rect 14274 8276 14280 8288
rect 12575 8248 14280 8276
rect 12575 8245 12587 8248
rect 12529 8239 12587 8245
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 14384 8276 14412 8316
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 15930 8276 15936 8288
rect 14384 8248 15936 8276
rect 15930 8236 15936 8248
rect 15988 8236 15994 8288
rect 16485 8279 16543 8285
rect 16485 8245 16497 8279
rect 16531 8276 16543 8279
rect 16669 8279 16727 8285
rect 16669 8276 16681 8279
rect 16531 8248 16681 8276
rect 16531 8245 16543 8248
rect 16485 8239 16543 8245
rect 16669 8245 16681 8248
rect 16715 8245 16727 8279
rect 18800 8276 18828 8375
rect 18966 8372 18972 8424
rect 19024 8412 19030 8424
rect 20714 8412 20720 8424
rect 19024 8384 20720 8412
rect 19024 8372 19030 8384
rect 20714 8372 20720 8384
rect 20772 8412 20778 8424
rect 21542 8412 21548 8424
rect 20772 8384 21548 8412
rect 20772 8372 20778 8384
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 22066 8412 22094 8452
rect 23290 8440 23296 8452
rect 23348 8440 23354 8492
rect 23385 8483 23443 8489
rect 23385 8449 23397 8483
rect 23431 8449 23443 8483
rect 23661 8483 23719 8489
rect 23661 8480 23673 8483
rect 23385 8443 23443 8449
rect 23492 8452 23673 8480
rect 21744 8384 22094 8412
rect 19306 8316 21588 8344
rect 19306 8276 19334 8316
rect 18800 8248 19334 8276
rect 16669 8239 16727 8245
rect 20346 8236 20352 8288
rect 20404 8276 20410 8288
rect 20441 8279 20499 8285
rect 20441 8276 20453 8279
rect 20404 8248 20453 8276
rect 20404 8236 20410 8248
rect 20441 8245 20453 8248
rect 20487 8245 20499 8279
rect 21560 8276 21588 8316
rect 21744 8276 21772 8384
rect 23198 8372 23204 8424
rect 23256 8412 23262 8424
rect 23400 8412 23428 8443
rect 23256 8384 23428 8412
rect 23256 8372 23262 8384
rect 23106 8304 23112 8356
rect 23164 8344 23170 8356
rect 23492 8344 23520 8452
rect 23661 8449 23673 8452
rect 23707 8480 23719 8483
rect 25406 8480 25412 8492
rect 23707 8452 25412 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 25406 8440 25412 8452
rect 25464 8440 25470 8492
rect 25501 8483 25559 8489
rect 25501 8449 25513 8483
rect 25547 8449 25559 8483
rect 25501 8443 25559 8449
rect 23566 8372 23572 8424
rect 23624 8412 23630 8424
rect 23750 8412 23756 8424
rect 23624 8384 23756 8412
rect 23624 8372 23630 8384
rect 23750 8372 23756 8384
rect 23808 8372 23814 8424
rect 23842 8372 23848 8424
rect 23900 8412 23906 8424
rect 25516 8412 25544 8443
rect 26142 8440 26148 8492
rect 26200 8440 26206 8492
rect 26694 8440 26700 8492
rect 26752 8480 26758 8492
rect 29196 8480 29224 8520
rect 30009 8517 30021 8520
rect 30055 8548 30067 8551
rect 30098 8548 30104 8560
rect 30055 8520 30104 8548
rect 30055 8517 30067 8520
rect 30009 8511 30067 8517
rect 30098 8508 30104 8520
rect 30156 8508 30162 8560
rect 30837 8551 30895 8557
rect 30837 8517 30849 8551
rect 30883 8548 30895 8551
rect 30926 8548 30932 8560
rect 30883 8520 30932 8548
rect 30883 8517 30895 8520
rect 30837 8511 30895 8517
rect 30926 8508 30932 8520
rect 30984 8508 30990 8560
rect 31021 8551 31079 8557
rect 31021 8517 31033 8551
rect 31067 8548 31079 8551
rect 31067 8520 32904 8548
rect 31067 8517 31079 8520
rect 31021 8511 31079 8517
rect 32876 8492 32904 8520
rect 26752 8452 29224 8480
rect 26752 8440 26758 8452
rect 29270 8440 29276 8492
rect 29328 8440 29334 8492
rect 29822 8440 29828 8492
rect 29880 8440 29886 8492
rect 30374 8440 30380 8492
rect 30432 8440 30438 8492
rect 30653 8483 30711 8489
rect 30653 8449 30665 8483
rect 30699 8480 30711 8483
rect 31113 8483 31171 8489
rect 30699 8452 31064 8480
rect 30699 8449 30711 8452
rect 30653 8443 30711 8449
rect 25682 8412 25688 8424
rect 23900 8384 25688 8412
rect 23900 8372 23906 8384
rect 25682 8372 25688 8384
rect 25740 8372 25746 8424
rect 25777 8415 25835 8421
rect 25777 8381 25789 8415
rect 25823 8412 25835 8415
rect 26050 8412 26056 8424
rect 25823 8384 26056 8412
rect 25823 8381 25835 8384
rect 25777 8375 25835 8381
rect 26050 8372 26056 8384
rect 26108 8372 26114 8424
rect 30282 8372 30288 8424
rect 30340 8412 30346 8424
rect 30469 8415 30527 8421
rect 30469 8412 30481 8415
rect 30340 8384 30481 8412
rect 30340 8372 30346 8384
rect 30469 8381 30481 8384
rect 30515 8381 30527 8415
rect 31036 8412 31064 8452
rect 31113 8449 31125 8483
rect 31159 8480 31171 8483
rect 31846 8480 31852 8492
rect 31159 8452 31852 8480
rect 31159 8449 31171 8452
rect 31113 8443 31171 8449
rect 31846 8440 31852 8452
rect 31904 8440 31910 8492
rect 32858 8440 32864 8492
rect 32916 8440 32922 8492
rect 33060 8489 33088 8576
rect 33045 8483 33103 8489
rect 33045 8449 33057 8483
rect 33091 8449 33103 8483
rect 33045 8443 33103 8449
rect 33505 8483 33563 8489
rect 33505 8449 33517 8483
rect 33551 8480 33563 8483
rect 33962 8480 33968 8492
rect 33551 8452 33968 8480
rect 33551 8449 33563 8452
rect 33505 8443 33563 8449
rect 32766 8412 32772 8424
rect 31036 8384 32772 8412
rect 30469 8375 30527 8381
rect 32766 8372 32772 8384
rect 32824 8372 32830 8424
rect 32950 8412 32956 8424
rect 32876 8384 32956 8412
rect 32876 8353 32904 8384
rect 32950 8372 32956 8384
rect 33008 8372 33014 8424
rect 33060 8412 33088 8443
rect 33962 8440 33968 8452
rect 34020 8440 34026 8492
rect 34146 8440 34152 8492
rect 34204 8440 34210 8492
rect 34422 8440 34428 8492
rect 34480 8480 34486 8492
rect 36096 8489 36124 8576
rect 36081 8483 36139 8489
rect 34480 8452 34730 8480
rect 34480 8440 34486 8452
rect 36081 8449 36093 8483
rect 36127 8449 36139 8483
rect 36081 8443 36139 8449
rect 33413 8415 33471 8421
rect 33413 8412 33425 8415
rect 33060 8384 33425 8412
rect 33413 8381 33425 8384
rect 33459 8381 33471 8415
rect 33413 8375 33471 8381
rect 34333 8415 34391 8421
rect 34333 8381 34345 8415
rect 34379 8412 34391 8415
rect 34514 8412 34520 8424
rect 34379 8384 34520 8412
rect 34379 8381 34391 8384
rect 34333 8375 34391 8381
rect 34514 8372 34520 8384
rect 34572 8372 34578 8424
rect 35066 8372 35072 8424
rect 35124 8412 35130 8424
rect 35805 8415 35863 8421
rect 35805 8412 35817 8415
rect 35124 8384 35817 8412
rect 35124 8372 35130 8384
rect 35805 8381 35817 8384
rect 35851 8381 35863 8415
rect 35805 8375 35863 8381
rect 30837 8347 30895 8353
rect 30837 8344 30849 8347
rect 23164 8316 23520 8344
rect 23676 8316 26096 8344
rect 23164 8304 23170 8316
rect 21560 8248 21772 8276
rect 20441 8239 20499 8245
rect 23290 8236 23296 8288
rect 23348 8276 23354 8288
rect 23676 8285 23704 8316
rect 23661 8279 23719 8285
rect 23661 8276 23673 8279
rect 23348 8248 23673 8276
rect 23348 8236 23354 8248
rect 23661 8245 23673 8248
rect 23707 8245 23719 8279
rect 23661 8239 23719 8245
rect 25682 8236 25688 8288
rect 25740 8236 25746 8288
rect 25774 8236 25780 8288
rect 25832 8276 25838 8288
rect 25961 8279 26019 8285
rect 25961 8276 25973 8279
rect 25832 8248 25973 8276
rect 25832 8236 25838 8248
rect 25961 8245 25973 8248
rect 26007 8245 26019 8279
rect 26068 8276 26096 8316
rect 28966 8316 30849 8344
rect 28966 8276 28994 8316
rect 30837 8313 30849 8316
rect 30883 8313 30895 8347
rect 30837 8307 30895 8313
rect 32861 8347 32919 8353
rect 32861 8313 32873 8347
rect 32907 8313 32919 8347
rect 32861 8307 32919 8313
rect 26068 8248 28994 8276
rect 25961 8239 26019 8245
rect 30098 8236 30104 8288
rect 30156 8276 30162 8288
rect 30193 8279 30251 8285
rect 30193 8276 30205 8279
rect 30156 8248 30205 8276
rect 30156 8236 30162 8248
rect 30193 8245 30205 8248
rect 30239 8245 30251 8279
rect 30193 8239 30251 8245
rect 34606 8236 34612 8288
rect 34664 8276 34670 8288
rect 35158 8276 35164 8288
rect 34664 8248 35164 8276
rect 34664 8236 34670 8248
rect 35158 8236 35164 8248
rect 35216 8236 35222 8288
rect 1104 8186 36432 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 36432 8186
rect 1104 8112 36432 8134
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3568 8044 4752 8072
rect 3568 8032 3574 8044
rect 4614 7964 4620 8016
rect 4672 7964 4678 8016
rect 4632 7936 4660 7964
rect 4356 7908 4660 7936
rect 4356 7877 4384 7908
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4724 7868 4752 8044
rect 5442 8032 5448 8084
rect 5500 8072 5506 8084
rect 6365 8075 6423 8081
rect 6365 8072 6377 8075
rect 5500 8044 6377 8072
rect 5500 8032 5506 8044
rect 6365 8041 6377 8044
rect 6411 8041 6423 8075
rect 6365 8035 6423 8041
rect 7561 8075 7619 8081
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 7650 8072 7656 8084
rect 7607 8044 7656 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 9030 8032 9036 8084
rect 9088 8032 9094 8084
rect 10042 8032 10048 8084
rect 10100 8032 10106 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 13262 8072 13268 8084
rect 10836 8044 13268 8072
rect 10836 8032 10842 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 14424 8044 15301 8072
rect 14424 8032 14430 8044
rect 15289 8041 15301 8044
rect 15335 8041 15347 8075
rect 15289 8035 15347 8041
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15841 8075 15899 8081
rect 15841 8072 15853 8075
rect 15436 8044 15853 8072
rect 15436 8032 15442 8044
rect 15841 8041 15853 8044
rect 15887 8072 15899 8075
rect 22094 8072 22100 8084
rect 15887 8044 22100 8072
rect 15887 8041 15899 8044
rect 15841 8035 15899 8041
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 23106 8032 23112 8084
rect 23164 8032 23170 8084
rect 23290 8032 23296 8084
rect 23348 8032 23354 8084
rect 23566 8032 23572 8084
rect 23624 8072 23630 8084
rect 24394 8072 24400 8084
rect 23624 8044 24400 8072
rect 23624 8032 23630 8044
rect 24394 8032 24400 8044
rect 24452 8072 24458 8084
rect 24452 8044 24716 8072
rect 24452 8032 24458 8044
rect 5629 8007 5687 8013
rect 5629 7973 5641 8007
rect 5675 8004 5687 8007
rect 6546 8004 6552 8016
rect 5675 7976 6552 8004
rect 5675 7973 5687 7976
rect 5629 7967 5687 7973
rect 6546 7964 6552 7976
rect 6604 8004 6610 8016
rect 9048 8004 9076 8032
rect 10413 8007 10471 8013
rect 10413 8004 10425 8007
rect 6604 7976 6955 8004
rect 9048 7976 10425 8004
rect 6604 7964 6610 7976
rect 5902 7896 5908 7948
rect 5960 7936 5966 7948
rect 6638 7936 6644 7948
rect 5960 7908 6644 7936
rect 5960 7896 5966 7908
rect 6638 7896 6644 7908
rect 6696 7936 6702 7948
rect 6696 7908 6868 7936
rect 6696 7896 6702 7908
rect 4663 7840 4752 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4540 7800 4568 7831
rect 4798 7828 4804 7880
rect 4856 7828 4862 7880
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 5460 7840 5733 7868
rect 4890 7800 4896 7812
rect 4540 7772 4896 7800
rect 4890 7760 4896 7772
rect 4948 7800 4954 7812
rect 5460 7800 5488 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5721 7831 5779 7837
rect 5828 7840 6009 7868
rect 4948 7772 5488 7800
rect 5629 7803 5687 7809
rect 4948 7760 4954 7772
rect 5629 7769 5641 7803
rect 5675 7800 5687 7803
rect 5828 7800 5856 7840
rect 5997 7837 6009 7840
rect 6043 7868 6055 7871
rect 6270 7868 6276 7880
rect 6043 7840 6276 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6730 7868 6736 7880
rect 6595 7840 6736 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 6840 7877 6868 7908
rect 6927 7877 6955 7976
rect 10413 7973 10425 7976
rect 10459 7973 10471 8007
rect 10413 7967 10471 7973
rect 13541 8007 13599 8013
rect 13541 7973 13553 8007
rect 13587 8004 13599 8007
rect 13814 8004 13820 8016
rect 13587 7976 13820 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 24302 8004 24308 8016
rect 14844 7976 24308 8004
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7936 7435 7939
rect 8662 7936 8668 7948
rect 7423 7908 8668 7936
rect 7423 7905 7435 7908
rect 7377 7899 7435 7905
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8812 7908 9045 7936
rect 8812 7896 8818 7908
rect 9033 7905 9045 7908
rect 9079 7936 9091 7939
rect 9398 7936 9404 7948
rect 9079 7908 9404 7936
rect 9079 7905 9091 7908
rect 9033 7899 9091 7905
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9490 7896 9496 7948
rect 9548 7936 9554 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 9548 7908 11161 7936
rect 9548 7896 9554 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 11422 7896 11428 7948
rect 11480 7896 11486 7948
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 14734 7936 14740 7948
rect 12768 7908 14740 7936
rect 12768 7896 12774 7908
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7868 7711 7871
rect 7742 7868 7748 7880
rect 7699 7840 7748 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 7742 7828 7748 7840
rect 7800 7868 7806 7880
rect 10134 7868 10140 7880
rect 7800 7840 10140 7868
rect 7800 7828 7806 7840
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 10284 7840 10333 7868
rect 10284 7828 10290 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10502 7828 10508 7880
rect 10560 7828 10566 7880
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 13648 7877 13676 7908
rect 14734 7896 14740 7908
rect 14792 7896 14798 7948
rect 13633 7871 13691 7877
rect 13633 7837 13645 7871
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 14182 7868 14188 7880
rect 14139 7840 14188 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 14844 7868 14872 7976
rect 24302 7964 24308 7976
rect 24360 7964 24366 8016
rect 17034 7936 17040 7948
rect 15028 7908 17040 7936
rect 14599 7840 14872 7868
rect 14916 7871 14974 7877
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 14916 7837 14928 7871
rect 14962 7868 14974 7871
rect 15028 7868 15056 7908
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 17310 7896 17316 7948
rect 17368 7936 17374 7948
rect 20254 7936 20260 7948
rect 17368 7908 20260 7936
rect 17368 7896 17374 7908
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 21910 7936 21916 7948
rect 20824 7908 21916 7936
rect 14962 7840 15056 7868
rect 14962 7837 14974 7840
rect 14916 7831 14974 7837
rect 5675 7772 5856 7800
rect 5905 7803 5963 7809
rect 5675 7769 5687 7772
rect 5629 7763 5687 7769
rect 5905 7769 5917 7803
rect 5951 7769 5963 7803
rect 5905 7763 5963 7769
rect 4154 7692 4160 7744
rect 4212 7692 4218 7744
rect 4706 7692 4712 7744
rect 4764 7692 4770 7744
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 5074 7732 5080 7744
rect 4856 7704 5080 7732
rect 4856 7692 4862 7704
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5445 7735 5503 7741
rect 5445 7701 5457 7735
rect 5491 7732 5503 7735
rect 5534 7732 5540 7744
rect 5491 7704 5540 7732
rect 5491 7701 5503 7704
rect 5445 7695 5503 7701
rect 5534 7692 5540 7704
rect 5592 7732 5598 7744
rect 5920 7732 5948 7763
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7926 7800 7932 7812
rect 7064 7772 7932 7800
rect 7064 7760 7070 7772
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 8662 7760 8668 7812
rect 8720 7800 8726 7812
rect 9217 7803 9275 7809
rect 9217 7800 9229 7803
rect 8720 7772 9229 7800
rect 8720 7760 8726 7772
rect 9217 7769 9229 7772
rect 9263 7769 9275 7803
rect 9217 7763 9275 7769
rect 9861 7803 9919 7809
rect 9861 7769 9873 7803
rect 9907 7800 9919 7803
rect 10778 7800 10784 7812
rect 9907 7772 10784 7800
rect 9907 7769 9919 7772
rect 9861 7763 9919 7769
rect 10778 7760 10784 7772
rect 10836 7760 10842 7812
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 11204 7772 11914 7800
rect 11204 7760 11210 7772
rect 5592 7704 5948 7732
rect 5997 7735 6055 7741
rect 5592 7692 5598 7704
rect 5997 7701 6009 7735
rect 6043 7732 6055 7735
rect 6270 7732 6276 7744
rect 6043 7704 6276 7732
rect 6043 7701 6055 7704
rect 5997 7695 6055 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 6733 7735 6791 7741
rect 6733 7701 6745 7735
rect 6779 7732 6791 7735
rect 7282 7732 7288 7744
rect 6779 7704 7288 7732
rect 6779 7701 6791 7704
rect 6733 7695 6791 7701
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 8110 7692 8116 7744
rect 8168 7732 8174 7744
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 8168 7704 9321 7732
rect 8168 7692 8174 7704
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9309 7695 9367 7701
rect 9677 7735 9735 7741
rect 9677 7701 9689 7735
rect 9723 7732 9735 7735
rect 10061 7735 10119 7741
rect 10061 7732 10073 7735
rect 9723 7704 10073 7732
rect 9723 7701 9735 7704
rect 9677 7695 9735 7701
rect 10061 7701 10073 7704
rect 10107 7701 10119 7735
rect 10061 7695 10119 7701
rect 10229 7735 10287 7741
rect 10229 7701 10241 7735
rect 10275 7732 10287 7735
rect 10318 7732 10324 7744
rect 10275 7704 10324 7732
rect 10275 7701 10287 7704
rect 10229 7695 10287 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 11808 7732 11836 7772
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 14384 7800 14412 7831
rect 13872 7772 14412 7800
rect 14476 7800 14504 7831
rect 15102 7828 15108 7880
rect 15160 7828 15166 7880
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15378 7868 15384 7880
rect 15335 7840 15384 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 19058 7868 19064 7880
rect 15988 7840 19064 7868
rect 15988 7828 15994 7840
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 20622 7868 20628 7880
rect 19392 7840 20628 7868
rect 19392 7828 19398 7840
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 20824 7877 20852 7908
rect 21910 7896 21916 7908
rect 21968 7896 21974 7948
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 23201 7939 23259 7945
rect 22152 7908 23060 7936
rect 22152 7896 22158 7908
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7837 20867 7871
rect 20809 7831 20867 7837
rect 21082 7828 21088 7880
rect 21140 7828 21146 7880
rect 21174 7828 21180 7880
rect 21232 7868 21238 7880
rect 22922 7868 22928 7880
rect 21232 7840 22928 7868
rect 21232 7828 21238 7840
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 23032 7877 23060 7908
rect 23201 7905 23213 7939
rect 23247 7936 23259 7939
rect 23750 7936 23756 7948
rect 23247 7908 23756 7936
rect 23247 7905 23259 7908
rect 23201 7899 23259 7905
rect 23750 7896 23756 7908
rect 23808 7896 23814 7948
rect 24578 7896 24584 7948
rect 24636 7896 24642 7948
rect 24688 7936 24716 8044
rect 25682 8032 25688 8084
rect 25740 8072 25746 8084
rect 25869 8075 25927 8081
rect 25869 8072 25881 8075
rect 25740 8044 25881 8072
rect 25740 8032 25746 8044
rect 25869 8041 25881 8044
rect 25915 8041 25927 8075
rect 25869 8035 25927 8041
rect 26970 8032 26976 8084
rect 27028 8072 27034 8084
rect 27246 8072 27252 8084
rect 27028 8044 27252 8072
rect 27028 8032 27034 8044
rect 27246 8032 27252 8044
rect 27304 8032 27310 8084
rect 29822 8032 29828 8084
rect 29880 8032 29886 8084
rect 30098 8032 30104 8084
rect 30156 8032 30162 8084
rect 33870 8032 33876 8084
rect 33928 8072 33934 8084
rect 35069 8075 35127 8081
rect 35069 8072 35081 8075
rect 33928 8044 35081 8072
rect 33928 8032 33934 8044
rect 35069 8041 35081 8044
rect 35115 8041 35127 8075
rect 35069 8035 35127 8041
rect 35342 8032 35348 8084
rect 35400 8032 35406 8084
rect 26142 7964 26148 8016
rect 26200 8004 26206 8016
rect 26789 8007 26847 8013
rect 26789 8004 26801 8007
rect 26200 7976 26801 8004
rect 26200 7964 26206 7976
rect 26789 7973 26801 7976
rect 26835 7973 26847 8007
rect 26789 7967 26847 7973
rect 24765 7939 24823 7945
rect 24765 7936 24777 7939
rect 24688 7908 24777 7936
rect 24765 7905 24777 7908
rect 24811 7905 24823 7939
rect 26881 7939 26939 7945
rect 24765 7899 24823 7905
rect 25424 7908 25912 7936
rect 23017 7871 23075 7877
rect 23017 7837 23029 7871
rect 23063 7837 23075 7871
rect 23017 7831 23075 7837
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 24489 7871 24547 7877
rect 24489 7837 24501 7871
rect 24535 7837 24547 7871
rect 24489 7831 24547 7837
rect 15013 7803 15071 7809
rect 14476 7772 14964 7800
rect 13872 7760 13878 7772
rect 12894 7732 12900 7744
rect 11808 7704 12900 7732
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 14737 7735 14795 7741
rect 14737 7732 14749 7735
rect 13412 7704 14749 7732
rect 13412 7692 13418 7704
rect 14737 7701 14749 7704
rect 14783 7701 14795 7735
rect 14936 7732 14964 7772
rect 15013 7769 15025 7803
rect 15059 7800 15071 7803
rect 15562 7800 15568 7812
rect 15059 7772 15568 7800
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 15562 7760 15568 7772
rect 15620 7760 15626 7812
rect 15746 7760 15752 7812
rect 15804 7800 15810 7812
rect 16942 7800 16948 7812
rect 15804 7772 16948 7800
rect 15804 7760 15810 7772
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 18690 7760 18696 7812
rect 18748 7800 18754 7812
rect 19242 7800 19248 7812
rect 18748 7772 19248 7800
rect 18748 7760 18754 7772
rect 19242 7760 19248 7772
rect 19300 7760 19306 7812
rect 19702 7760 19708 7812
rect 19760 7800 19766 7812
rect 19760 7772 21036 7800
rect 19760 7760 19766 7772
rect 20530 7732 20536 7744
rect 14936 7704 20536 7732
rect 14737 7695 14795 7701
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 20625 7735 20683 7741
rect 20625 7701 20637 7735
rect 20671 7732 20683 7735
rect 20714 7732 20720 7744
rect 20671 7704 20720 7732
rect 20671 7701 20683 7704
rect 20625 7695 20683 7701
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 21008 7741 21036 7772
rect 20993 7735 21051 7741
rect 20993 7701 21005 7735
rect 21039 7732 21051 7735
rect 22462 7732 22468 7744
rect 21039 7704 22468 7732
rect 21039 7701 21051 7704
rect 20993 7695 21051 7701
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 22741 7735 22799 7741
rect 22741 7701 22753 7735
rect 22787 7732 22799 7735
rect 23014 7732 23020 7744
rect 22787 7704 23020 7732
rect 22787 7701 22799 7704
rect 22741 7695 22799 7701
rect 23014 7692 23020 7704
rect 23072 7692 23078 7744
rect 24504 7732 24532 7831
rect 24596 7800 24624 7896
rect 24670 7828 24676 7880
rect 24728 7828 24734 7880
rect 25314 7828 25320 7880
rect 25372 7828 25378 7880
rect 25424 7812 25452 7908
rect 25498 7828 25504 7880
rect 25556 7828 25562 7880
rect 25682 7828 25688 7880
rect 25740 7828 25746 7880
rect 25774 7828 25780 7880
rect 25832 7828 25838 7880
rect 25884 7877 25912 7908
rect 26881 7905 26893 7939
rect 26927 7936 26939 7939
rect 26970 7936 26976 7948
rect 26927 7908 26976 7936
rect 26927 7905 26939 7908
rect 26881 7899 26939 7905
rect 26970 7896 26976 7908
rect 27028 7896 27034 7948
rect 27798 7896 27804 7948
rect 27856 7896 27862 7948
rect 28000 7908 28212 7936
rect 25869 7871 25927 7877
rect 25869 7837 25881 7871
rect 25915 7837 25927 7871
rect 25869 7831 25927 7837
rect 26050 7828 26056 7880
rect 26108 7828 26114 7880
rect 26329 7871 26387 7877
rect 26329 7868 26341 7871
rect 26153 7840 26341 7868
rect 25222 7800 25228 7812
rect 24596 7772 25228 7800
rect 25222 7760 25228 7772
rect 25280 7760 25286 7812
rect 25406 7760 25412 7812
rect 25464 7760 25470 7812
rect 24854 7732 24860 7744
rect 24504 7704 24860 7732
rect 24854 7692 24860 7704
rect 24912 7692 24918 7744
rect 24946 7692 24952 7744
rect 25004 7692 25010 7744
rect 25038 7692 25044 7744
rect 25096 7732 25102 7744
rect 25133 7735 25191 7741
rect 25133 7732 25145 7735
rect 25096 7704 25145 7732
rect 25096 7692 25102 7704
rect 25133 7701 25145 7704
rect 25179 7701 25191 7735
rect 25240 7732 25268 7760
rect 26153 7732 26181 7840
rect 26329 7837 26341 7840
rect 26375 7837 26387 7871
rect 26329 7831 26387 7837
rect 26421 7871 26479 7877
rect 26421 7837 26433 7871
rect 26467 7868 26479 7871
rect 26510 7868 26516 7880
rect 26467 7840 26516 7868
rect 26467 7837 26479 7840
rect 26421 7831 26479 7837
rect 26510 7828 26516 7840
rect 26568 7828 26574 7880
rect 27246 7828 27252 7880
rect 27304 7868 27310 7880
rect 27433 7871 27491 7877
rect 27433 7868 27445 7871
rect 27304 7840 27445 7868
rect 27304 7828 27310 7840
rect 27433 7837 27445 7840
rect 27479 7837 27491 7871
rect 27433 7831 27491 7837
rect 27709 7871 27767 7877
rect 27709 7837 27721 7871
rect 27755 7837 27767 7871
rect 27709 7831 27767 7837
rect 26602 7760 26608 7812
rect 26660 7800 26666 7812
rect 27341 7803 27399 7809
rect 27341 7800 27353 7803
rect 26660 7772 27353 7800
rect 26660 7760 26666 7772
rect 27341 7769 27353 7772
rect 27387 7769 27399 7803
rect 27724 7800 27752 7831
rect 27890 7828 27896 7880
rect 27948 7828 27954 7880
rect 28000 7800 28028 7908
rect 28077 7871 28135 7877
rect 28077 7837 28089 7871
rect 28123 7837 28135 7871
rect 28077 7831 28135 7837
rect 27724 7772 28028 7800
rect 27341 7763 27399 7769
rect 25240 7704 26181 7732
rect 25133 7695 25191 7701
rect 26786 7692 26792 7744
rect 26844 7732 26850 7744
rect 28092 7732 28120 7831
rect 28184 7800 28212 7908
rect 28534 7896 28540 7948
rect 28592 7896 28598 7948
rect 29840 7936 29868 8032
rect 30009 8007 30067 8013
rect 30009 7973 30021 8007
rect 30055 8004 30067 8007
rect 30282 8004 30288 8016
rect 30055 7976 30288 8004
rect 30055 7973 30067 7976
rect 30009 7967 30067 7973
rect 30282 7964 30288 7976
rect 30340 7964 30346 8016
rect 30374 7964 30380 8016
rect 30432 8004 30438 8016
rect 30469 8007 30527 8013
rect 30469 8004 30481 8007
rect 30432 7976 30481 8004
rect 30432 7964 30438 7976
rect 30469 7973 30481 7976
rect 30515 8004 30527 8007
rect 32214 8004 32220 8016
rect 30515 7976 32220 8004
rect 30515 7973 30527 7976
rect 30469 7967 30527 7973
rect 32214 7964 32220 7976
rect 32272 7964 32278 8016
rect 34790 7964 34796 8016
rect 34848 8004 34854 8016
rect 35161 8007 35219 8013
rect 35161 8004 35173 8007
rect 34848 7976 35173 8004
rect 34848 7964 34854 7976
rect 35161 7973 35173 7976
rect 35207 7973 35219 8007
rect 35161 7967 35219 7973
rect 28644 7908 29868 7936
rect 29917 7939 29975 7945
rect 28644 7877 28672 7908
rect 29917 7905 29929 7939
rect 29963 7936 29975 7939
rect 30834 7936 30840 7948
rect 29963 7908 30840 7936
rect 29963 7905 29975 7908
rect 29917 7899 29975 7905
rect 30834 7896 30840 7908
rect 30892 7896 30898 7948
rect 35253 7939 35311 7945
rect 35253 7905 35265 7939
rect 35299 7936 35311 7939
rect 35434 7936 35440 7948
rect 35299 7908 35440 7936
rect 35299 7905 35311 7908
rect 35253 7899 35311 7905
rect 35434 7896 35440 7908
rect 35492 7896 35498 7948
rect 28629 7871 28687 7877
rect 28629 7837 28641 7871
rect 28675 7837 28687 7871
rect 28629 7831 28687 7837
rect 28718 7828 28724 7880
rect 28776 7868 28782 7880
rect 30561 7871 30619 7877
rect 28776 7840 30328 7868
rect 28776 7828 28782 7840
rect 29822 7800 29828 7812
rect 28184 7772 29828 7800
rect 29822 7760 29828 7772
rect 29880 7760 29886 7812
rect 30300 7800 30328 7840
rect 30561 7837 30573 7871
rect 30607 7837 30619 7871
rect 30561 7831 30619 7837
rect 30576 7800 30604 7831
rect 30926 7828 30932 7880
rect 30984 7828 30990 7880
rect 31113 7871 31171 7877
rect 31113 7837 31125 7871
rect 31159 7868 31171 7871
rect 32858 7868 32864 7880
rect 31159 7840 32864 7868
rect 31159 7837 31171 7840
rect 31113 7831 31171 7837
rect 32858 7828 32864 7840
rect 32916 7828 32922 7880
rect 33410 7828 33416 7880
rect 33468 7868 33474 7880
rect 34701 7871 34759 7877
rect 34701 7868 34713 7871
rect 33468 7840 34713 7868
rect 33468 7828 33474 7840
rect 34701 7837 34713 7840
rect 34747 7837 34759 7871
rect 34701 7831 34759 7837
rect 31018 7800 31024 7812
rect 30300 7772 31024 7800
rect 31018 7760 31024 7772
rect 31076 7800 31082 7812
rect 31846 7800 31852 7812
rect 31076 7772 31852 7800
rect 31076 7760 31082 7772
rect 31846 7760 31852 7772
rect 31904 7760 31910 7812
rect 29270 7732 29276 7744
rect 26844 7704 29276 7732
rect 26844 7692 26850 7704
rect 29270 7692 29276 7704
rect 29328 7692 29334 7744
rect 30650 7692 30656 7744
rect 30708 7692 30714 7744
rect 1104 7642 36432 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 36432 7642
rect 1104 7568 36432 7590
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 4338 7528 4344 7540
rect 2271 7500 4344 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4614 7528 4620 7540
rect 4479 7500 4620 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5258 7528 5264 7540
rect 5215 7500 5264 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 5997 7531 6055 7537
rect 5997 7528 6009 7531
rect 5868 7500 6009 7528
rect 5868 7488 5874 7500
rect 5997 7497 6009 7500
rect 6043 7528 6055 7531
rect 6730 7528 6736 7540
rect 6043 7500 6736 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7466 7488 7472 7540
rect 7524 7528 7530 7540
rect 8481 7531 8539 7537
rect 8481 7528 8493 7531
rect 7524 7500 8493 7528
rect 7524 7488 7530 7500
rect 8481 7497 8493 7500
rect 8527 7497 8539 7531
rect 8481 7491 8539 7497
rect 8938 7488 8944 7540
rect 8996 7528 9002 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8996 7500 9137 7528
rect 8996 7488 9002 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 10502 7528 10508 7540
rect 9125 7491 9183 7497
rect 9508 7500 10508 7528
rect 2958 7420 2964 7472
rect 3016 7420 3022 7472
rect 7006 7460 7012 7472
rect 3988 7432 7012 7460
rect 3988 7401 4016 7432
rect 7006 7420 7012 7432
rect 7064 7460 7070 7472
rect 8386 7460 8392 7472
rect 7064 7432 8392 7460
rect 7064 7420 7070 7432
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 4522 7352 4528 7404
rect 4580 7352 4586 7404
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 5316 7364 5365 7392
rect 5316 7352 5322 7364
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5442 7352 5448 7404
rect 5500 7352 5506 7404
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 4709 7327 4767 7333
rect 3743 7296 4108 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 4080 7265 4108 7296
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 4798 7324 4804 7336
rect 4755 7296 4804 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 5460 7324 5488 7352
rect 5224 7296 5488 7324
rect 5224 7284 5230 7296
rect 4065 7259 4123 7265
rect 4065 7225 4077 7259
rect 4111 7225 4123 7259
rect 4065 7219 4123 7225
rect 5552 7188 5580 7355
rect 5736 7256 5764 7355
rect 5828 7324 5856 7355
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 7190 7352 7196 7404
rect 7248 7352 7254 7404
rect 7760 7401 7788 7432
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 8754 7420 8760 7472
rect 8812 7420 8818 7472
rect 8846 7420 8852 7472
rect 8904 7420 8910 7472
rect 9398 7420 9404 7472
rect 9456 7460 9462 7472
rect 9508 7469 9536 7500
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 10597 7531 10655 7537
rect 10597 7497 10609 7531
rect 10643 7528 10655 7531
rect 10870 7528 10876 7540
rect 10643 7500 10876 7528
rect 10643 7497 10655 7500
rect 10597 7491 10655 7497
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 12710 7528 12716 7540
rect 11900 7500 12716 7528
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 9456 7432 9505 7460
rect 9456 7420 9462 7432
rect 9493 7429 9505 7432
rect 9539 7429 9551 7463
rect 9493 7423 9551 7429
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 9824 7432 10272 7460
rect 9824 7420 9830 7432
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 9030 7352 9036 7404
rect 9088 7352 9094 7404
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9582 7392 9588 7404
rect 9355 7364 9588 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 5994 7324 6000 7336
rect 5828 7296 6000 7324
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 6362 7284 6368 7336
rect 6420 7284 6426 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6472 7296 6929 7324
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 5736 7228 6193 7256
rect 6181 7225 6193 7228
rect 6227 7225 6239 7259
rect 6181 7219 6239 7225
rect 5994 7188 6000 7200
rect 5552 7160 6000 7188
rect 5994 7148 6000 7160
rect 6052 7188 6058 7200
rect 6472 7188 6500 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 9324 7324 9352 7355
rect 9582 7352 9588 7364
rect 9640 7392 9646 7404
rect 9861 7395 9919 7401
rect 9640 7352 9674 7392
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10042 7392 10048 7404
rect 9907 7364 10048 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10244 7401 10272 7432
rect 10318 7420 10324 7472
rect 10376 7460 10382 7472
rect 11900 7469 11928 7500
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 13446 7528 13452 7540
rect 13004 7500 13452 7528
rect 11885 7463 11943 7469
rect 10376 7432 10548 7460
rect 10376 7420 10382 7432
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 7984 7296 9352 7324
rect 7984 7284 7990 7296
rect 6638 7216 6644 7268
rect 6696 7216 6702 7268
rect 7009 7259 7067 7265
rect 7009 7225 7021 7259
rect 7055 7256 7067 7259
rect 8570 7256 8576 7268
rect 7055 7228 8576 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 9646 7256 9674 7352
rect 10152 7256 10180 7355
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 10520 7401 10548 7432
rect 11885 7429 11897 7463
rect 11931 7429 11943 7463
rect 11885 7423 11943 7429
rect 11977 7463 12035 7469
rect 11977 7429 11989 7463
rect 12023 7460 12035 7463
rect 12618 7460 12624 7472
rect 12023 7432 12624 7460
rect 12023 7429 12035 7432
rect 11977 7423 12035 7429
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 13004 7460 13032 7500
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 14093 7531 14151 7537
rect 14093 7497 14105 7531
rect 14139 7528 14151 7531
rect 14182 7528 14188 7540
rect 14139 7500 14188 7528
rect 14139 7497 14151 7500
rect 14093 7491 14151 7497
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 15657 7531 15715 7537
rect 15657 7497 15669 7531
rect 15703 7528 15715 7531
rect 15746 7528 15752 7540
rect 15703 7500 15752 7528
rect 15703 7497 15715 7500
rect 15657 7491 15715 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16666 7488 16672 7540
rect 16724 7488 16730 7540
rect 18138 7488 18144 7540
rect 18196 7488 18202 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 18874 7528 18880 7540
rect 18656 7500 18880 7528
rect 18656 7488 18662 7500
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 19518 7528 19524 7540
rect 19076 7500 19524 7528
rect 14369 7463 14427 7469
rect 12952 7432 13110 7460
rect 12952 7420 12958 7432
rect 14369 7429 14381 7463
rect 14415 7460 14427 7463
rect 14550 7460 14556 7472
rect 14415 7432 14556 7460
rect 14415 7429 14427 7432
rect 14369 7423 14427 7429
rect 14550 7420 14556 7432
rect 14608 7420 14614 7472
rect 14734 7420 14740 7472
rect 14792 7420 14798 7472
rect 15194 7420 15200 7472
rect 15252 7460 15258 7472
rect 17310 7460 17316 7472
rect 15252 7432 17316 7460
rect 15252 7420 15258 7432
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7392 10931 7395
rect 11422 7392 11428 7404
rect 10919 7364 11428 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11422 7352 11428 7364
rect 11480 7352 11486 7404
rect 11606 7352 11612 7404
rect 11664 7352 11670 7404
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 12101 7395 12159 7401
rect 12101 7361 12113 7395
rect 12147 7392 12159 7395
rect 12250 7392 12256 7404
rect 12147 7364 12256 7392
rect 12147 7361 12159 7364
rect 12101 7355 12159 7361
rect 10778 7284 10784 7336
rect 10836 7284 10842 7336
rect 10962 7284 10968 7336
rect 11020 7284 11026 7336
rect 11054 7284 11060 7336
rect 11112 7284 11118 7336
rect 11716 7324 11744 7355
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14752 7392 14780 7420
rect 14332 7364 14780 7392
rect 15473 7395 15531 7401
rect 14332 7352 14338 7364
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16482 7392 16488 7404
rect 15795 7364 16488 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 11790 7324 11796 7336
rect 11716 7296 11796 7324
rect 11716 7256 11744 7296
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 12176 7296 12357 7324
rect 9646 7228 10088 7256
rect 10152 7228 11744 7256
rect 6052 7160 6500 7188
rect 6052 7148 6058 7160
rect 6822 7148 6828 7200
rect 6880 7148 6886 7200
rect 7377 7191 7435 7197
rect 7377 7157 7389 7191
rect 7423 7188 7435 7191
rect 8202 7188 8208 7200
rect 7423 7160 8208 7188
rect 7423 7157 7435 7160
rect 7377 7151 7435 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 9766 7148 9772 7200
rect 9824 7148 9830 7200
rect 9950 7148 9956 7200
rect 10008 7148 10014 7200
rect 10060 7188 10088 7228
rect 10226 7188 10232 7200
rect 10060 7160 10232 7188
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 11698 7188 11704 7200
rect 10376 7160 11704 7188
rect 10376 7148 10382 7160
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12176 7188 12204 7296
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 12618 7284 12624 7336
rect 12676 7284 12682 7336
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 14642 7324 14648 7336
rect 12768 7296 14648 7324
rect 12768 7284 12774 7296
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 15488 7256 15516 7355
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16868 7401 16896 7432
rect 17310 7420 17316 7432
rect 17368 7420 17374 7472
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 18104 7432 18736 7460
rect 18104 7420 18110 7432
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17126 7352 17132 7404
rect 17184 7352 17190 7404
rect 18230 7352 18236 7404
rect 18288 7392 18294 7404
rect 18708 7401 18736 7432
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18288 7364 18613 7392
rect 18288 7352 18294 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7361 18751 7395
rect 18693 7355 18751 7361
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 19076 7392 19104 7500
rect 19518 7488 19524 7500
rect 19576 7528 19582 7540
rect 20257 7531 20315 7537
rect 19576 7500 20024 7528
rect 19576 7488 19582 7500
rect 19426 7420 19432 7472
rect 19484 7460 19490 7472
rect 19702 7460 19708 7472
rect 19484 7432 19708 7460
rect 19484 7420 19490 7432
rect 19702 7420 19708 7432
rect 19760 7420 19766 7472
rect 19905 7463 19963 7469
rect 19905 7460 19917 7463
rect 19904 7429 19917 7460
rect 19951 7429 19963 7463
rect 19996 7460 20024 7500
rect 20257 7497 20269 7531
rect 20303 7528 20315 7531
rect 20438 7528 20444 7540
rect 20303 7500 20444 7528
rect 20303 7497 20315 7500
rect 20257 7491 20315 7497
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 24946 7528 24952 7540
rect 20588 7500 22094 7528
rect 20588 7488 20594 7500
rect 21082 7460 21088 7472
rect 19996 7432 21088 7460
rect 19904 7423 19963 7429
rect 18923 7364 19104 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 19150 7352 19156 7404
rect 19208 7352 19214 7404
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 19904 7392 19932 7423
rect 21082 7420 21088 7432
rect 21140 7420 21146 7472
rect 21821 7463 21879 7469
rect 21821 7429 21833 7463
rect 21867 7460 21879 7463
rect 21910 7460 21916 7472
rect 21867 7432 21916 7460
rect 21867 7429 21879 7432
rect 21821 7423 21879 7429
rect 21910 7420 21916 7432
rect 21968 7420 21974 7472
rect 22066 7460 22094 7500
rect 22940 7500 24952 7528
rect 22066 7432 22784 7460
rect 19300 7364 19932 7392
rect 19300 7352 19306 7364
rect 17037 7327 17095 7333
rect 17037 7293 17049 7327
rect 17083 7324 17095 7327
rect 17218 7324 17224 7336
rect 17083 7296 17224 7324
rect 17083 7293 17095 7296
rect 17037 7287 17095 7293
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 19168 7324 19196 7352
rect 18432 7296 19196 7324
rect 19904 7324 19932 7364
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 20622 7392 20628 7404
rect 20487 7364 20628 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 20772 7364 20944 7392
rect 20772 7352 20778 7364
rect 20916 7324 20944 7364
rect 21634 7352 21640 7404
rect 21692 7352 21698 7404
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 22370 7392 22376 7404
rect 22327 7364 22376 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 22462 7352 22468 7404
rect 22520 7352 22526 7404
rect 19904 7296 20852 7324
rect 20916 7296 22094 7324
rect 18432 7265 18460 7296
rect 18417 7259 18475 7265
rect 18417 7256 18429 7259
rect 15488 7228 18429 7256
rect 18417 7225 18429 7228
rect 18463 7225 18475 7259
rect 18417 7219 18475 7225
rect 18509 7259 18567 7265
rect 18509 7225 18521 7259
rect 18555 7256 18567 7259
rect 19150 7256 19156 7268
rect 18555 7228 19156 7256
rect 18555 7225 18567 7228
rect 18509 7219 18567 7225
rect 19150 7216 19156 7228
rect 19208 7216 19214 7268
rect 20714 7256 20720 7268
rect 19260 7228 20720 7256
rect 12124 7160 12204 7188
rect 12124 7148 12130 7160
rect 12250 7148 12256 7200
rect 12308 7148 12314 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 15473 7191 15531 7197
rect 15473 7188 15485 7191
rect 15436 7160 15485 7188
rect 15436 7148 15442 7160
rect 15473 7157 15485 7160
rect 15519 7157 15531 7191
rect 15473 7151 15531 7157
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 17129 7191 17187 7197
rect 17129 7188 17141 7191
rect 16632 7160 17141 7188
rect 16632 7148 16638 7160
rect 17129 7157 17141 7160
rect 17175 7188 17187 7191
rect 19260 7188 19288 7228
rect 20714 7216 20720 7228
rect 20772 7216 20778 7268
rect 17175 7160 19288 7188
rect 17175 7157 17187 7160
rect 17129 7151 17187 7157
rect 19886 7148 19892 7200
rect 19944 7148 19950 7200
rect 20070 7148 20076 7200
rect 20128 7148 20134 7200
rect 20824 7188 20852 7296
rect 22066 7268 22094 7296
rect 22066 7228 22100 7268
rect 22094 7216 22100 7228
rect 22152 7216 22158 7268
rect 22189 7259 22247 7265
rect 22189 7225 22201 7259
rect 22235 7225 22247 7259
rect 22480 7256 22508 7352
rect 22756 7324 22784 7432
rect 22830 7352 22836 7404
rect 22888 7352 22894 7404
rect 22940 7401 22968 7500
rect 24946 7488 24952 7500
rect 25004 7488 25010 7540
rect 26234 7488 26240 7540
rect 26292 7528 26298 7540
rect 27430 7528 27436 7540
rect 26292 7500 27436 7528
rect 26292 7488 26298 7500
rect 27430 7488 27436 7500
rect 27488 7528 27494 7540
rect 27801 7531 27859 7537
rect 27801 7528 27813 7531
rect 27488 7500 27813 7528
rect 27488 7488 27494 7500
rect 27801 7497 27813 7500
rect 27847 7497 27859 7531
rect 27801 7491 27859 7497
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 30837 7531 30895 7537
rect 30837 7528 30849 7531
rect 27948 7500 30849 7528
rect 27948 7488 27954 7500
rect 30837 7497 30849 7500
rect 30883 7528 30895 7531
rect 30926 7528 30932 7540
rect 30883 7500 30932 7528
rect 30883 7497 30895 7500
rect 30837 7491 30895 7497
rect 30926 7488 30932 7500
rect 30984 7488 30990 7540
rect 31294 7488 31300 7540
rect 31352 7528 31358 7540
rect 31757 7531 31815 7537
rect 31757 7528 31769 7531
rect 31352 7500 31769 7528
rect 31352 7488 31358 7500
rect 31757 7497 31769 7500
rect 31803 7497 31815 7531
rect 31757 7491 31815 7497
rect 25038 7460 25044 7472
rect 23124 7432 25044 7460
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7361 22983 7395
rect 22925 7355 22983 7361
rect 23014 7352 23020 7404
rect 23072 7352 23078 7404
rect 23124 7401 23152 7432
rect 25038 7420 25044 7432
rect 25096 7420 25102 7472
rect 25682 7460 25688 7472
rect 25148 7432 25688 7460
rect 25148 7401 25176 7432
rect 25682 7420 25688 7432
rect 25740 7460 25746 7472
rect 28074 7460 28080 7472
rect 25740 7432 28080 7460
rect 25740 7420 25746 7432
rect 23109 7395 23167 7401
rect 23109 7361 23121 7395
rect 23155 7361 23167 7395
rect 23109 7355 23167 7361
rect 24949 7395 25007 7401
rect 24949 7361 24961 7395
rect 24995 7361 25007 7395
rect 24949 7355 25007 7361
rect 25133 7395 25191 7401
rect 25133 7361 25145 7395
rect 25179 7361 25191 7395
rect 25133 7355 25191 7361
rect 24964 7324 24992 7355
rect 25222 7352 25228 7404
rect 25280 7392 25286 7404
rect 25501 7395 25559 7401
rect 25501 7392 25513 7395
rect 25280 7364 25513 7392
rect 25280 7352 25286 7364
rect 25501 7361 25513 7364
rect 25547 7392 25559 7395
rect 25590 7392 25596 7404
rect 25547 7364 25596 7392
rect 25547 7361 25559 7364
rect 25501 7355 25559 7361
rect 25590 7352 25596 7364
rect 25648 7352 25654 7404
rect 25777 7395 25835 7401
rect 25777 7361 25789 7395
rect 25823 7392 25835 7395
rect 26142 7392 26148 7404
rect 25823 7364 26148 7392
rect 25823 7361 25835 7364
rect 25777 7355 25835 7361
rect 26142 7352 26148 7364
rect 26200 7352 26206 7404
rect 27724 7401 27752 7432
rect 28074 7420 28080 7432
rect 28132 7420 28138 7472
rect 30944 7460 30972 7488
rect 30944 7432 31708 7460
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 27890 7352 27896 7404
rect 27948 7352 27954 7404
rect 30834 7352 30840 7404
rect 30892 7392 30898 7404
rect 31021 7395 31079 7401
rect 31021 7392 31033 7395
rect 30892 7364 31033 7392
rect 30892 7352 30898 7364
rect 31021 7361 31033 7364
rect 31067 7392 31079 7395
rect 31067 7364 31340 7392
rect 31067 7361 31079 7364
rect 31021 7355 31079 7361
rect 25406 7324 25412 7336
rect 22756 7296 25412 7324
rect 23658 7256 23664 7268
rect 22480 7228 23664 7256
rect 22189 7219 22247 7225
rect 21453 7191 21511 7197
rect 21453 7188 21465 7191
rect 20824 7160 21465 7188
rect 21453 7157 21465 7160
rect 21499 7188 21511 7191
rect 22204 7188 22232 7219
rect 23658 7216 23664 7228
rect 23716 7216 23722 7268
rect 24946 7216 24952 7268
rect 25004 7216 25010 7268
rect 25332 7265 25360 7296
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 25682 7284 25688 7336
rect 25740 7324 25746 7336
rect 26970 7324 26976 7336
rect 25740 7296 26976 7324
rect 25740 7284 25746 7296
rect 26970 7284 26976 7296
rect 27028 7284 27034 7336
rect 25317 7259 25375 7265
rect 25317 7225 25329 7259
rect 25363 7225 25375 7259
rect 30650 7256 30656 7268
rect 25317 7219 25375 7225
rect 25424 7228 30656 7256
rect 21499 7160 22232 7188
rect 21499 7157 21511 7160
rect 21453 7151 21511 7157
rect 22646 7148 22652 7200
rect 22704 7148 22710 7200
rect 23474 7148 23480 7200
rect 23532 7188 23538 7200
rect 25424 7188 25452 7228
rect 30650 7216 30656 7228
rect 30708 7216 30714 7268
rect 23532 7160 25452 7188
rect 23532 7148 23538 7160
rect 25498 7148 25504 7200
rect 25556 7188 25562 7200
rect 25777 7191 25835 7197
rect 25777 7188 25789 7191
rect 25556 7160 25789 7188
rect 25556 7148 25562 7160
rect 25777 7157 25789 7160
rect 25823 7188 25835 7191
rect 26510 7188 26516 7200
rect 25823 7160 26516 7188
rect 25823 7157 25835 7160
rect 25777 7151 25835 7157
rect 26510 7148 26516 7160
rect 26568 7148 26574 7200
rect 27062 7148 27068 7200
rect 27120 7188 27126 7200
rect 27522 7188 27528 7200
rect 27120 7160 27528 7188
rect 27120 7148 27126 7160
rect 27522 7148 27528 7160
rect 27580 7148 27586 7200
rect 30834 7148 30840 7200
rect 30892 7188 30898 7200
rect 31021 7191 31079 7197
rect 31021 7188 31033 7191
rect 30892 7160 31033 7188
rect 30892 7148 30898 7160
rect 31021 7157 31033 7160
rect 31067 7157 31079 7191
rect 31312 7188 31340 7364
rect 31386 7352 31392 7404
rect 31444 7352 31450 7404
rect 31680 7401 31708 7432
rect 33042 7420 33048 7472
rect 33100 7420 33106 7472
rect 31665 7395 31723 7401
rect 31665 7361 31677 7395
rect 31711 7361 31723 7395
rect 31665 7355 31723 7361
rect 31846 7352 31852 7404
rect 31904 7392 31910 7404
rect 32309 7395 32367 7401
rect 32309 7392 32321 7395
rect 31904 7364 32321 7392
rect 31904 7352 31910 7364
rect 32309 7361 32321 7364
rect 32355 7361 32367 7395
rect 32309 7355 32367 7361
rect 32858 7352 32864 7404
rect 32916 7352 32922 7404
rect 31481 7327 31539 7333
rect 31481 7293 31493 7327
rect 31527 7293 31539 7327
rect 31481 7287 31539 7293
rect 31496 7256 31524 7287
rect 31662 7256 31668 7268
rect 31496 7228 31668 7256
rect 31662 7216 31668 7228
rect 31720 7216 31726 7268
rect 31478 7188 31484 7200
rect 31312 7160 31484 7188
rect 31021 7151 31079 7157
rect 31478 7148 31484 7160
rect 31536 7188 31542 7200
rect 32490 7188 32496 7200
rect 31536 7160 32496 7188
rect 31536 7148 31542 7160
rect 32490 7148 32496 7160
rect 32548 7148 32554 7200
rect 1104 7098 36432 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 36432 7098
rect 1104 7024 36432 7046
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 3970 6984 3976 6996
rect 3016 6956 3976 6984
rect 3016 6944 3022 6956
rect 3970 6944 3976 6956
rect 4028 6944 4034 6996
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 4614 6984 4620 6996
rect 4571 6956 4620 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 5166 6984 5172 6996
rect 4856 6956 5172 6984
rect 4856 6944 4862 6956
rect 5166 6944 5172 6956
rect 5224 6984 5230 6996
rect 5902 6984 5908 6996
rect 5224 6956 5908 6984
rect 5224 6944 5230 6956
rect 4706 6916 4712 6928
rect 4172 6888 4712 6916
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4172 6848 4200 6888
rect 4706 6876 4712 6888
rect 4764 6876 4770 6928
rect 5828 6916 5856 6956
rect 5902 6944 5908 6956
rect 5960 6984 5966 6996
rect 5960 6956 7052 6984
rect 5960 6944 5966 6956
rect 4908 6888 5672 6916
rect 4908 6857 4936 6888
rect 5644 6860 5672 6888
rect 5736 6888 5856 6916
rect 4111 6820 4200 6848
rect 4249 6851 4307 6857
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4617 6851 4675 6857
rect 4617 6848 4629 6851
rect 4295 6820 4629 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4617 6817 4629 6820
rect 4663 6817 4675 6851
rect 4893 6851 4951 6857
rect 4893 6848 4905 6851
rect 4617 6811 4675 6817
rect 4724 6820 4905 6848
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3568 6752 4169 6780
rect 3568 6740 3574 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4338 6740 4344 6792
rect 4396 6740 4402 6792
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 4724 6780 4752 6820
rect 4893 6817 4905 6820
rect 4939 6817 4951 6851
rect 4893 6811 4951 6817
rect 4985 6851 5043 6857
rect 4985 6817 4997 6851
rect 5031 6848 5043 6851
rect 5031 6820 5580 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 5552 6792 5580 6820
rect 5626 6808 5632 6860
rect 5684 6808 5690 6860
rect 4488 6752 4752 6780
rect 4488 6740 4494 6752
rect 4798 6740 4804 6792
rect 4856 6740 4862 6792
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 5092 6712 5120 6743
rect 4304 6684 5120 6712
rect 5276 6712 5304 6743
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 5736 6789 5764 6888
rect 6730 6876 6736 6928
rect 6788 6916 6794 6928
rect 7024 6916 7052 6956
rect 8570 6944 8576 6996
rect 8628 6944 8634 6996
rect 9756 6987 9814 6993
rect 9756 6953 9768 6987
rect 9802 6984 9814 6987
rect 9950 6984 9956 6996
rect 9802 6956 9956 6984
rect 9802 6953 9814 6956
rect 9756 6947 9814 6953
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 10468 6956 11008 6984
rect 10468 6944 10474 6956
rect 6788 6888 6960 6916
rect 7024 6888 7880 6916
rect 6788 6876 6794 6888
rect 6932 6857 6960 6888
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 5859 6820 6837 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 6918 6851 6976 6857
rect 6918 6817 6930 6851
rect 6964 6817 6976 6851
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6918 6811 6976 6817
rect 7006 6817 7021 6848
rect 7055 6817 7067 6851
rect 7852 6848 7880 6888
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 10980 6916 11008 6956
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11609 6987 11667 6993
rect 11609 6984 11621 6987
rect 11112 6956 11621 6984
rect 11112 6944 11118 6956
rect 11609 6953 11621 6956
rect 11655 6953 11667 6987
rect 11609 6947 11667 6953
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 12989 6987 13047 6993
rect 12989 6984 13001 6987
rect 12676 6956 13001 6984
rect 12676 6944 12682 6956
rect 12989 6953 13001 6956
rect 13035 6953 13047 6987
rect 12989 6947 13047 6953
rect 13354 6944 13360 6996
rect 13412 6944 13418 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13872 6956 14105 6984
rect 13872 6944 13878 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 17773 6987 17831 6993
rect 17773 6984 17785 6987
rect 17276 6956 17785 6984
rect 17276 6944 17282 6956
rect 17773 6953 17785 6956
rect 17819 6984 17831 6987
rect 17862 6984 17868 6996
rect 17819 6956 17868 6984
rect 17819 6953 17831 6956
rect 17773 6947 17831 6953
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 17957 6987 18015 6993
rect 17957 6953 17969 6987
rect 18003 6984 18015 6987
rect 19886 6984 19892 6996
rect 18003 6956 19892 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 19886 6944 19892 6956
rect 19944 6944 19950 6996
rect 20714 6944 20720 6996
rect 20772 6984 20778 6996
rect 21634 6984 21640 6996
rect 20772 6956 21640 6984
rect 20772 6944 20778 6956
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 22094 6944 22100 6996
rect 22152 6984 22158 6996
rect 25314 6984 25320 6996
rect 22152 6956 25320 6984
rect 22152 6944 22158 6956
rect 25314 6944 25320 6956
rect 25372 6984 25378 6996
rect 25866 6984 25872 6996
rect 25372 6956 25872 6984
rect 25372 6944 25378 6956
rect 25866 6944 25872 6956
rect 25924 6944 25930 6996
rect 26418 6944 26424 6996
rect 26476 6984 26482 6996
rect 27065 6987 27123 6993
rect 27065 6984 27077 6987
rect 26476 6956 27077 6984
rect 26476 6944 26482 6956
rect 27065 6953 27077 6956
rect 27111 6953 27123 6987
rect 27065 6947 27123 6953
rect 13538 6916 13544 6928
rect 8260 6888 9628 6916
rect 10980 6888 13544 6916
rect 8260 6876 8266 6888
rect 7852 6820 8064 6848
rect 7006 6811 7067 6817
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6749 5779 6783
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 5721 6743 5779 6749
rect 6012 6752 6101 6780
rect 5442 6712 5448 6724
rect 5276 6684 5448 6712
rect 4304 6672 4310 6684
rect 5092 6644 5120 6684
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 5902 6672 5908 6724
rect 5960 6672 5966 6724
rect 6012 6644 6040 6752
rect 6089 6749 6101 6752
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 6328 6752 6377 6780
rect 6328 6740 6334 6752
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 6546 6740 6552 6792
rect 6604 6780 6610 6792
rect 7006 6780 7034 6811
rect 6604 6752 7034 6780
rect 6604 6740 6610 6752
rect 7006 6712 7034 6752
rect 7094 6783 7152 6789
rect 7094 6749 7106 6783
rect 7140 6774 7152 6783
rect 7466 6780 7472 6792
rect 7299 6774 7472 6780
rect 7140 6752 7472 6774
rect 7140 6749 7327 6752
rect 7094 6746 7327 6749
rect 7094 6743 7152 6746
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7650 6740 7656 6792
rect 7708 6740 7714 6792
rect 7926 6740 7932 6792
rect 7984 6740 7990 6792
rect 8036 6780 8064 6820
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 9490 6848 9496 6860
rect 8444 6820 9496 6848
rect 8444 6808 8450 6820
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9600 6848 9628 6888
rect 13538 6876 13544 6888
rect 13596 6876 13602 6928
rect 18233 6919 18291 6925
rect 18233 6916 18245 6919
rect 17696 6888 18245 6916
rect 10318 6848 10324 6860
rect 9600 6820 10324 6848
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 10962 6848 10968 6860
rect 10468 6820 10968 6848
rect 10468 6808 10474 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11514 6808 11520 6860
rect 11572 6848 11578 6860
rect 13814 6848 13820 6860
rect 11572 6820 12434 6848
rect 11572 6808 11578 6820
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8036 6752 8493 6780
rect 8481 6749 8493 6752
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6780 8723 6783
rect 8846 6780 8852 6792
rect 8711 6752 8852 6780
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 8680 6712 8708 6743
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 7006 6684 8708 6712
rect 8956 6712 8984 6743
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11793 6783 11851 6789
rect 11793 6780 11805 6783
rect 11112 6752 11805 6780
rect 11112 6740 11118 6752
rect 11793 6749 11805 6752
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 12158 6780 12164 6792
rect 12115 6752 12164 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 8956 6684 10088 6712
rect 5092 6616 6040 6644
rect 6273 6647 6331 6653
rect 6273 6613 6285 6647
rect 6319 6644 6331 6647
rect 6546 6644 6552 6656
rect 6319 6616 6552 6644
rect 6319 6613 6331 6616
rect 6273 6607 6331 6613
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 6641 6647 6699 6653
rect 6641 6613 6653 6647
rect 6687 6644 6699 6647
rect 7190 6644 7196 6656
rect 6687 6616 7196 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7466 6644 7472 6656
rect 7331 6616 7472 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 9030 6644 9036 6656
rect 8536 6616 9036 6644
rect 8536 6604 8542 6616
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 9309 6647 9367 6653
rect 9309 6613 9321 6647
rect 9355 6644 9367 6647
rect 9950 6644 9956 6656
rect 9355 6616 9956 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10060 6644 10088 6684
rect 10226 6672 10232 6724
rect 10284 6672 10290 6724
rect 11238 6672 11244 6724
rect 11296 6712 11302 6724
rect 11882 6712 11888 6724
rect 11296 6684 11888 6712
rect 11296 6672 11302 6684
rect 11882 6672 11888 6684
rect 11940 6712 11946 6724
rect 11992 6712 12020 6743
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 12406 6780 12434 6820
rect 12820 6820 13820 6848
rect 12820 6780 12848 6820
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 13924 6820 14473 6848
rect 12406 6752 12848 6780
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 12986 6780 12992 6792
rect 12943 6752 12992 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13170 6740 13176 6792
rect 13228 6740 13234 6792
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 13924 6789 13952 6820
rect 14461 6817 14473 6820
rect 14507 6848 14519 6851
rect 17126 6848 17132 6860
rect 14507 6820 17132 6848
rect 14507 6817 14519 6820
rect 14461 6811 14519 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 17696 6848 17724 6888
rect 18233 6885 18245 6888
rect 18279 6885 18291 6919
rect 18785 6919 18843 6925
rect 18785 6916 18797 6919
rect 18233 6879 18291 6885
rect 18524 6888 18797 6916
rect 17368 6820 17724 6848
rect 17368 6808 17374 6820
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 18524 6848 18552 6888
rect 18785 6885 18797 6888
rect 18831 6885 18843 6919
rect 18785 6879 18843 6885
rect 19521 6919 19579 6925
rect 19521 6885 19533 6919
rect 19567 6916 19579 6919
rect 20070 6916 20076 6928
rect 19567 6888 20076 6916
rect 19567 6885 19579 6888
rect 19521 6879 19579 6885
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 24210 6876 24216 6928
rect 24268 6916 24274 6928
rect 25774 6916 25780 6928
rect 24268 6888 25780 6916
rect 24268 6876 24274 6888
rect 25774 6876 25780 6888
rect 25832 6876 25838 6928
rect 27080 6916 27108 6947
rect 27522 6944 27528 6996
rect 27580 6944 27586 6996
rect 32585 6987 32643 6993
rect 32585 6953 32597 6987
rect 32631 6984 32643 6987
rect 32858 6984 32864 6996
rect 32631 6956 32864 6984
rect 32631 6953 32643 6956
rect 32585 6947 32643 6953
rect 32858 6944 32864 6956
rect 32916 6944 32922 6996
rect 28810 6916 28816 6928
rect 27080 6888 28816 6916
rect 28810 6876 28816 6888
rect 28868 6876 28874 6928
rect 32769 6919 32827 6925
rect 32769 6885 32781 6919
rect 32815 6885 32827 6919
rect 34790 6916 34796 6928
rect 32769 6879 32827 6885
rect 34348 6888 34796 6916
rect 17920 6820 18552 6848
rect 17920 6808 17926 6820
rect 18598 6808 18604 6860
rect 18656 6808 18662 6860
rect 18693 6851 18751 6857
rect 18693 6817 18705 6851
rect 18739 6817 18751 6851
rect 18693 6811 18751 6817
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 12434 6712 12440 6724
rect 11940 6684 12440 6712
rect 11940 6672 11946 6684
rect 12434 6672 12440 6684
rect 12492 6712 12498 6724
rect 13541 6715 13599 6721
rect 13541 6712 13553 6715
rect 12492 6684 13553 6712
rect 12492 6672 12498 6684
rect 13541 6681 13553 6684
rect 13587 6681 13599 6715
rect 13740 6712 13768 6743
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14292 6712 14320 6740
rect 13740 6684 14320 6712
rect 14568 6712 14596 6743
rect 18506 6740 18512 6792
rect 18564 6740 18570 6792
rect 18708 6780 18736 6811
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 19613 6851 19671 6857
rect 19613 6848 19625 6851
rect 18932 6820 19625 6848
rect 18932 6808 18938 6820
rect 19613 6817 19625 6820
rect 19659 6817 19671 6851
rect 19613 6811 19671 6817
rect 22002 6808 22008 6860
rect 22060 6848 22066 6860
rect 24118 6848 24124 6860
rect 22060 6820 24124 6848
rect 22060 6808 22066 6820
rect 24118 6808 24124 6820
rect 24176 6848 24182 6860
rect 25866 6848 25872 6860
rect 24176 6820 25872 6848
rect 24176 6808 24182 6820
rect 25866 6808 25872 6820
rect 25924 6808 25930 6860
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 26384 6820 27568 6848
rect 26384 6808 26390 6820
rect 18616 6752 18736 6780
rect 18969 6783 19027 6789
rect 17218 6712 17224 6724
rect 14568 6684 17224 6712
rect 13541 6675 13599 6681
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 18046 6712 18052 6724
rect 17328 6684 18052 6712
rect 10410 6644 10416 6656
rect 10060 6616 10416 6644
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 12253 6647 12311 6653
rect 12253 6644 12265 6647
rect 11204 6616 12265 6644
rect 11204 6604 11210 6616
rect 12253 6613 12265 6616
rect 12299 6613 12311 6647
rect 12253 6607 12311 6613
rect 13354 6604 13360 6656
rect 13412 6644 13418 6656
rect 13906 6644 13912 6656
rect 13412 6616 13912 6644
rect 13412 6604 13418 6616
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 17328 6644 17356 6684
rect 18046 6672 18052 6684
rect 18104 6712 18110 6724
rect 18141 6715 18199 6721
rect 18141 6712 18153 6715
rect 18104 6684 18153 6712
rect 18104 6672 18110 6684
rect 18141 6681 18153 6684
rect 18187 6681 18199 6715
rect 18141 6675 18199 6681
rect 18230 6672 18236 6724
rect 18288 6712 18294 6724
rect 18616 6712 18644 6752
rect 18969 6749 18981 6783
rect 19015 6780 19027 6783
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19015 6752 19441 6780
rect 19015 6749 19027 6752
rect 18969 6743 19027 6749
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 18288 6684 18644 6712
rect 18288 6672 18294 6684
rect 18874 6672 18880 6724
rect 18932 6712 18938 6724
rect 19444 6712 19472 6743
rect 19702 6740 19708 6792
rect 19760 6780 19766 6792
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 19760 6752 19901 6780
rect 19760 6740 19766 6752
rect 19889 6749 19901 6752
rect 19935 6749 19947 6783
rect 19889 6743 19947 6749
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6780 20315 6783
rect 20438 6780 20444 6792
rect 20303 6752 20444 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 20438 6740 20444 6752
rect 20496 6740 20502 6792
rect 20530 6740 20536 6792
rect 20588 6780 20594 6792
rect 20588 6752 27476 6780
rect 20588 6740 20594 6752
rect 21450 6712 21456 6724
rect 18932 6684 19380 6712
rect 19444 6684 21456 6712
rect 18932 6672 18938 6684
rect 14700 6616 17356 6644
rect 17957 6647 18015 6653
rect 14700 6604 14706 6616
rect 17957 6613 17969 6647
rect 18003 6644 18015 6647
rect 18690 6644 18696 6656
rect 18003 6616 18696 6644
rect 18003 6613 18015 6616
rect 17957 6607 18015 6613
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19242 6604 19248 6656
rect 19300 6604 19306 6656
rect 19352 6644 19380 6684
rect 21450 6672 21456 6684
rect 21508 6672 21514 6724
rect 22922 6672 22928 6724
rect 22980 6712 22986 6724
rect 26878 6712 26884 6724
rect 22980 6684 26884 6712
rect 22980 6672 22986 6684
rect 26878 6672 26884 6684
rect 26936 6672 26942 6724
rect 19610 6644 19616 6656
rect 19352 6616 19616 6644
rect 19610 6604 19616 6616
rect 19668 6604 19674 6656
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 21542 6644 21548 6656
rect 20864 6616 21548 6644
rect 20864 6604 20870 6616
rect 21542 6604 21548 6616
rect 21600 6644 21606 6656
rect 25406 6644 25412 6656
rect 21600 6616 25412 6644
rect 21600 6604 21606 6616
rect 25406 6604 25412 6616
rect 25464 6604 25470 6656
rect 26234 6604 26240 6656
rect 26292 6644 26298 6656
rect 27062 6644 27068 6656
rect 27120 6653 27126 6656
rect 27120 6647 27144 6653
rect 26292 6616 27068 6644
rect 26292 6604 26298 6616
rect 27062 6604 27068 6616
rect 27132 6613 27144 6647
rect 27120 6607 27144 6613
rect 27120 6604 27126 6607
rect 27246 6604 27252 6656
rect 27304 6604 27310 6656
rect 27338 6604 27344 6656
rect 27396 6604 27402 6656
rect 27448 6644 27476 6752
rect 27540 6721 27568 6820
rect 29914 6808 29920 6860
rect 29972 6808 29978 6860
rect 32490 6808 32496 6860
rect 32548 6848 32554 6860
rect 32677 6851 32735 6857
rect 32677 6848 32689 6851
rect 32548 6820 32689 6848
rect 32548 6808 32554 6820
rect 32677 6817 32689 6820
rect 32723 6817 32735 6851
rect 32784 6848 32812 6879
rect 33870 6848 33876 6860
rect 32784 6820 33876 6848
rect 32677 6811 32735 6817
rect 33870 6808 33876 6820
rect 33928 6808 33934 6860
rect 29822 6740 29828 6792
rect 29880 6740 29886 6792
rect 30009 6783 30067 6789
rect 30009 6749 30021 6783
rect 30055 6780 30067 6783
rect 32858 6780 32864 6792
rect 30055 6774 31754 6780
rect 31864 6774 32864 6780
rect 30055 6752 32864 6774
rect 30055 6749 30067 6752
rect 30009 6743 30067 6749
rect 31726 6746 31892 6752
rect 32858 6740 32864 6752
rect 32916 6740 32922 6792
rect 33137 6783 33195 6789
rect 33137 6749 33149 6783
rect 33183 6749 33195 6783
rect 33137 6743 33195 6749
rect 33229 6783 33287 6789
rect 33229 6749 33241 6783
rect 33275 6780 33287 6783
rect 33410 6780 33416 6792
rect 33275 6752 33416 6780
rect 33275 6749 33287 6752
rect 33229 6743 33287 6749
rect 27509 6715 27568 6721
rect 27509 6681 27521 6715
rect 27555 6684 27568 6715
rect 27555 6681 27567 6684
rect 27509 6675 27567 6681
rect 27614 6672 27620 6724
rect 27672 6712 27678 6724
rect 27709 6715 27767 6721
rect 27709 6712 27721 6715
rect 27672 6684 27721 6712
rect 27672 6672 27678 6684
rect 27709 6681 27721 6684
rect 27755 6681 27767 6715
rect 27709 6675 27767 6681
rect 31386 6672 31392 6724
rect 31444 6712 31450 6724
rect 33152 6712 33180 6743
rect 33410 6740 33416 6752
rect 33468 6740 33474 6792
rect 34348 6712 34376 6888
rect 34790 6876 34796 6888
rect 34848 6876 34854 6928
rect 31444 6684 34376 6712
rect 31444 6672 31450 6684
rect 29086 6644 29092 6656
rect 27448 6616 29092 6644
rect 29086 6604 29092 6616
rect 29144 6644 29150 6656
rect 30558 6644 30564 6656
rect 29144 6616 30564 6644
rect 29144 6604 29150 6616
rect 30558 6604 30564 6616
rect 30616 6604 30622 6656
rect 31662 6604 31668 6656
rect 31720 6644 31726 6656
rect 33870 6644 33876 6656
rect 31720 6616 33876 6644
rect 31720 6604 31726 6616
rect 33870 6604 33876 6616
rect 33928 6604 33934 6656
rect 1104 6554 36432 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 36432 6554
rect 1104 6480 36432 6502
rect 4338 6400 4344 6452
rect 4396 6400 4402 6452
rect 5077 6443 5135 6449
rect 5077 6409 5089 6443
rect 5123 6440 5135 6443
rect 5258 6440 5264 6452
rect 5123 6412 5264 6440
rect 5123 6409 5135 6412
rect 5077 6403 5135 6409
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5350 6400 5356 6452
rect 5408 6400 5414 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5902 6440 5908 6452
rect 5592 6412 5908 6440
rect 5592 6400 5598 6412
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 6236 6412 6469 6440
rect 6236 6400 6242 6412
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 6457 6403 6515 6409
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 7650 6440 7656 6452
rect 6880 6412 7656 6440
rect 6880 6400 6886 6412
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 8754 6400 8760 6452
rect 8812 6400 8818 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 11333 6443 11391 6449
rect 10008 6412 11192 6440
rect 10008 6400 10014 6412
rect 5169 6375 5227 6381
rect 5169 6372 5181 6375
rect 4172 6344 5181 6372
rect 4172 6316 4200 6344
rect 5169 6341 5181 6344
rect 5215 6341 5227 6375
rect 5169 6335 5227 6341
rect 5368 6344 6316 6372
rect 4154 6264 4160 6316
rect 4212 6264 4218 6316
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4338 6304 4344 6316
rect 4295 6276 4344 6304
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 4614 6304 4620 6316
rect 4479 6276 4620 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 4890 6304 4896 6316
rect 4755 6276 4896 6304
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5368 6313 5396 6344
rect 6288 6316 6316 6344
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 7285 6375 7343 6381
rect 7285 6372 7297 6375
rect 7248 6344 7297 6372
rect 7248 6332 7254 6344
rect 7285 6341 7297 6344
rect 7331 6341 7343 6375
rect 7285 6335 7343 6341
rect 7742 6332 7748 6384
rect 7800 6332 7806 6384
rect 9033 6375 9091 6381
rect 9033 6341 9045 6375
rect 9079 6372 9091 6375
rect 9766 6372 9772 6384
rect 9079 6344 9772 6372
rect 9079 6341 9091 6344
rect 9033 6335 9091 6341
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 11164 6372 11192 6412
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11514 6440 11520 6452
rect 11379 6412 11520 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 13170 6440 13176 6452
rect 12299 6412 13176 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13538 6400 13544 6452
rect 13596 6400 13602 6452
rect 13630 6400 13636 6452
rect 13688 6440 13694 6452
rect 13725 6443 13783 6449
rect 13725 6440 13737 6443
rect 13688 6412 13737 6440
rect 13688 6400 13694 6412
rect 13725 6409 13737 6412
rect 13771 6409 13783 6443
rect 13725 6403 13783 6409
rect 14090 6400 14096 6452
rect 14148 6400 14154 6452
rect 17310 6440 17316 6452
rect 14200 6412 17316 6440
rect 12066 6372 12072 6384
rect 11164 6344 12072 6372
rect 12066 6332 12072 6344
rect 12124 6372 12130 6384
rect 12897 6375 12955 6381
rect 12897 6372 12909 6375
rect 12124 6344 12909 6372
rect 12124 6332 12130 6344
rect 12897 6341 12909 6344
rect 12943 6341 12955 6375
rect 14200 6372 14228 6412
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 17678 6440 17684 6452
rect 17460 6412 17684 6440
rect 17460 6400 17466 6412
rect 17678 6400 17684 6412
rect 17736 6440 17742 6452
rect 18141 6443 18199 6449
rect 17736 6412 18000 6440
rect 17736 6400 17742 6412
rect 15102 6372 15108 6384
rect 12897 6335 12955 6341
rect 13096 6344 14228 6372
rect 14292 6344 15108 6372
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 5491 6276 5764 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6236 4859 6239
rect 5258 6236 5264 6248
rect 4847 6208 5264 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 5626 6196 5632 6248
rect 5684 6196 5690 6248
rect 5736 6236 5764 6276
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6328 6276 6377 6304
rect 6328 6264 6334 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 6564 6236 6592 6264
rect 5736 6208 6592 6236
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8720 6208 9137 6236
rect 8720 6196 8726 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9324 6236 9352 6267
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9548 6276 9597 6304
rect 9548 6264 9554 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 11606 6304 11612 6316
rect 10994 6276 11612 6304
rect 9585 6267 9643 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6304 12403 6307
rect 12434 6304 12440 6316
rect 12391 6276 12440 6304
rect 12391 6273 12403 6276
rect 12345 6267 12403 6273
rect 9861 6239 9919 6245
rect 9324 6208 9628 6236
rect 9125 6199 9183 6205
rect 9600 6180 9628 6208
rect 9861 6205 9873 6239
rect 9907 6236 9919 6239
rect 10870 6236 10876 6248
rect 9907 6208 10876 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 12176 6236 12204 6267
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6273 12863 6307
rect 12805 6267 12863 6273
rect 12710 6236 12716 6248
rect 10980 6208 12204 6236
rect 12268 6208 12716 6236
rect 10980 6180 11008 6208
rect 9582 6128 9588 6180
rect 9640 6128 9646 6180
rect 10962 6128 10968 6180
rect 11020 6128 11026 6180
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5442 6100 5448 6112
rect 4948 6072 5448 6100
rect 4948 6060 4954 6072
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 7432 6072 9045 6100
rect 7432 6060 7438 6072
rect 9033 6069 9045 6072
rect 9079 6100 9091 6103
rect 9398 6100 9404 6112
rect 9079 6072 9404 6100
rect 9079 6069 9091 6072
rect 9033 6063 9091 6069
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 9493 6103 9551 6109
rect 9493 6069 9505 6103
rect 9539 6100 9551 6103
rect 10042 6100 10048 6112
rect 9539 6072 10048 6100
rect 9539 6069 9551 6072
rect 9493 6063 9551 6069
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 12268 6100 12296 6208
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 12820 6236 12848 6267
rect 12894 6236 12900 6248
rect 12820 6208 12900 6236
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 13096 6245 13124 6344
rect 13262 6264 13268 6316
rect 13320 6264 13326 6316
rect 13814 6264 13820 6316
rect 13872 6264 13878 6316
rect 14292 6313 14320 6344
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 15197 6375 15255 6381
rect 15197 6341 15209 6375
rect 15243 6372 15255 6375
rect 15413 6375 15471 6381
rect 15243 6344 15332 6372
rect 15243 6341 15255 6344
rect 15197 6335 15255 6341
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 13081 6239 13139 6245
rect 13081 6205 13093 6239
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6236 13599 6239
rect 13722 6236 13728 6248
rect 13587 6208 13728 6236
rect 13587 6205 13599 6208
rect 13541 6199 13599 6205
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 14384 6236 14412 6267
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 15304 6304 15332 6344
rect 15413 6341 15425 6375
rect 15459 6372 15471 6375
rect 16206 6372 16212 6384
rect 15459 6344 16212 6372
rect 15459 6341 15471 6344
rect 15413 6335 15471 6341
rect 16206 6332 16212 6344
rect 16264 6332 16270 6384
rect 16942 6332 16948 6384
rect 17000 6372 17006 6384
rect 17972 6381 18000 6412
rect 18141 6409 18153 6443
rect 18187 6440 18199 6443
rect 18322 6440 18328 6452
rect 18187 6412 18328 6440
rect 18187 6409 18199 6412
rect 18141 6403 18199 6409
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 19610 6440 19616 6452
rect 18432 6412 19616 6440
rect 17773 6375 17831 6381
rect 17773 6372 17785 6375
rect 17000 6344 17785 6372
rect 17000 6332 17006 6344
rect 17773 6341 17785 6344
rect 17819 6372 17831 6375
rect 17972 6375 18031 6381
rect 17819 6344 17908 6372
rect 17972 6344 17985 6375
rect 17819 6341 17831 6344
rect 17773 6335 17831 6341
rect 17880 6316 17908 6344
rect 17973 6341 17985 6344
rect 18019 6372 18031 6375
rect 18432 6372 18460 6412
rect 19610 6400 19616 6412
rect 19668 6440 19674 6452
rect 20530 6440 20536 6452
rect 19668 6412 20536 6440
rect 19668 6400 19674 6412
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 21361 6443 21419 6449
rect 21361 6409 21373 6443
rect 21407 6440 21419 6443
rect 21450 6440 21456 6452
rect 21407 6412 21456 6440
rect 21407 6409 21419 6412
rect 21361 6403 21419 6409
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 21634 6400 21640 6452
rect 21692 6440 21698 6452
rect 23569 6443 23627 6449
rect 23569 6440 23581 6443
rect 21692 6412 23581 6440
rect 21692 6400 21698 6412
rect 23569 6409 23581 6412
rect 23615 6409 23627 6443
rect 23569 6403 23627 6409
rect 23750 6400 23756 6452
rect 23808 6440 23814 6452
rect 23937 6443 23995 6449
rect 23937 6440 23949 6443
rect 23808 6412 23949 6440
rect 23808 6400 23814 6412
rect 23937 6409 23949 6412
rect 23983 6440 23995 6443
rect 24670 6440 24676 6452
rect 23983 6412 24676 6440
rect 23983 6409 23995 6412
rect 23937 6403 23995 6409
rect 24670 6400 24676 6412
rect 24728 6440 24734 6452
rect 24765 6443 24823 6449
rect 24765 6440 24777 6443
rect 24728 6412 24777 6440
rect 24728 6400 24734 6412
rect 24765 6409 24777 6412
rect 24811 6409 24823 6443
rect 24765 6403 24823 6409
rect 25866 6400 25872 6452
rect 25924 6440 25930 6452
rect 26253 6443 26311 6449
rect 26253 6440 26265 6443
rect 25924 6412 26265 6440
rect 25924 6400 25930 6412
rect 26253 6409 26265 6412
rect 26299 6409 26311 6443
rect 26253 6403 26311 6409
rect 26421 6443 26479 6449
rect 26421 6409 26433 6443
rect 26467 6440 26479 6443
rect 26467 6412 28120 6440
rect 26467 6409 26479 6412
rect 26421 6403 26479 6409
rect 19334 6372 19340 6384
rect 18019 6344 18460 6372
rect 18524 6344 18828 6372
rect 18019 6341 18031 6344
rect 17973 6335 18031 6341
rect 15654 6304 15660 6316
rect 15304 6276 15660 6304
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18524 6304 18552 6344
rect 17920 6276 18552 6304
rect 18601 6307 18659 6313
rect 17920 6264 17926 6276
rect 18601 6273 18613 6307
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 16298 6236 16304 6248
rect 14384 6208 16304 6236
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 17126 6196 17132 6248
rect 17184 6236 17190 6248
rect 18230 6236 18236 6248
rect 17184 6208 18236 6236
rect 17184 6196 17190 6208
rect 18230 6196 18236 6208
rect 18288 6236 18294 6248
rect 18325 6239 18383 6245
rect 18325 6236 18337 6239
rect 18288 6208 18337 6236
rect 18288 6196 18294 6208
rect 18325 6205 18337 6208
rect 18371 6205 18383 6239
rect 18616 6236 18644 6267
rect 18690 6264 18696 6316
rect 18748 6264 18754 6316
rect 18800 6313 18828 6344
rect 18892 6344 19340 6372
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 18892 6236 18920 6344
rect 19334 6332 19340 6344
rect 19392 6332 19398 6384
rect 20993 6375 21051 6381
rect 20993 6341 21005 6375
rect 21039 6372 21051 6375
rect 21082 6372 21088 6384
rect 21039 6344 21088 6372
rect 21039 6341 21051 6344
rect 20993 6335 21051 6341
rect 21082 6332 21088 6344
rect 21140 6332 21146 6384
rect 21209 6375 21267 6381
rect 21209 6341 21221 6375
rect 21255 6372 21267 6375
rect 21542 6372 21548 6384
rect 21255 6344 21548 6372
rect 21255 6341 21267 6344
rect 21209 6335 21267 6341
rect 21542 6332 21548 6344
rect 21600 6332 21606 6384
rect 21818 6332 21824 6384
rect 21876 6372 21882 6384
rect 21876 6344 23888 6372
rect 21876 6332 21882 6344
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19702 6304 19708 6316
rect 19024 6276 19708 6304
rect 19024 6264 19030 6276
rect 19702 6264 19708 6276
rect 19760 6304 19766 6316
rect 20898 6304 20904 6316
rect 19760 6276 20904 6304
rect 19760 6264 19766 6276
rect 20898 6264 20904 6276
rect 20956 6264 20962 6316
rect 21100 6304 21128 6332
rect 23106 6304 23112 6316
rect 21100 6276 23112 6304
rect 23106 6264 23112 6276
rect 23164 6264 23170 6316
rect 23860 6313 23888 6344
rect 24026 6332 24032 6384
rect 24084 6332 24090 6384
rect 25038 6372 25044 6384
rect 24320 6344 25044 6372
rect 23845 6307 23903 6313
rect 23845 6273 23857 6307
rect 23891 6304 23903 6307
rect 24118 6304 24124 6316
rect 23891 6276 24124 6304
rect 23891 6273 23903 6276
rect 23845 6267 23903 6273
rect 24118 6264 24124 6276
rect 24176 6264 24182 6316
rect 24320 6313 24348 6344
rect 25038 6332 25044 6344
rect 25096 6372 25102 6384
rect 25096 6344 25636 6372
rect 25096 6332 25102 6344
rect 25608 6316 25636 6344
rect 26050 6332 26056 6384
rect 26108 6332 26114 6384
rect 27246 6332 27252 6384
rect 27304 6372 27310 6384
rect 27304 6344 27752 6372
rect 27304 6332 27310 6344
rect 24305 6307 24363 6313
rect 24305 6273 24317 6307
rect 24351 6273 24363 6307
rect 24305 6267 24363 6273
rect 24670 6264 24676 6316
rect 24728 6313 24734 6316
rect 24728 6304 24737 6313
rect 24857 6307 24915 6313
rect 24728 6276 24773 6304
rect 24728 6267 24737 6276
rect 24857 6273 24869 6307
rect 24903 6304 24915 6307
rect 25317 6307 25375 6313
rect 25317 6304 25329 6307
rect 24903 6276 25329 6304
rect 24903 6273 24915 6276
rect 24857 6267 24915 6273
rect 25317 6273 25329 6276
rect 25363 6273 25375 6307
rect 25317 6267 25375 6273
rect 24728 6264 24734 6267
rect 22738 6236 22744 6248
rect 18616 6208 18920 6236
rect 19306 6208 22744 6236
rect 18325 6199 18383 6205
rect 12342 6128 12348 6180
rect 12400 6168 12406 6180
rect 13357 6171 13415 6177
rect 13357 6168 13369 6171
rect 12400 6140 13369 6168
rect 12400 6128 12406 6140
rect 13357 6137 13369 6140
rect 13403 6137 13415 6171
rect 13357 6131 13415 6137
rect 13906 6128 13912 6180
rect 13964 6168 13970 6180
rect 15746 6168 15752 6180
rect 13964 6140 15752 6168
rect 13964 6128 13970 6140
rect 15746 6128 15752 6140
rect 15804 6128 15810 6180
rect 15838 6128 15844 6180
rect 15896 6168 15902 6180
rect 19306 6168 19334 6208
rect 22738 6196 22744 6208
rect 22796 6196 22802 6248
rect 15896 6140 19334 6168
rect 24949 6171 25007 6177
rect 15896 6128 15902 6140
rect 24949 6137 24961 6171
rect 24995 6137 25007 6171
rect 25332 6168 25360 6267
rect 25498 6264 25504 6316
rect 25556 6264 25562 6316
rect 25590 6264 25596 6316
rect 25648 6304 25654 6316
rect 25777 6307 25835 6313
rect 25777 6304 25789 6307
rect 25648 6276 25789 6304
rect 25648 6264 25654 6276
rect 25777 6273 25789 6276
rect 25823 6273 25835 6307
rect 25777 6267 25835 6273
rect 27338 6264 27344 6316
rect 27396 6264 27402 6316
rect 27724 6313 27752 6344
rect 28092 6313 28120 6412
rect 28810 6400 28816 6452
rect 28868 6440 28874 6452
rect 29457 6443 29515 6449
rect 29457 6440 29469 6443
rect 28868 6412 29469 6440
rect 28868 6400 28874 6412
rect 29457 6409 29469 6412
rect 29503 6409 29515 6443
rect 29457 6403 29515 6409
rect 29917 6443 29975 6449
rect 29917 6409 29929 6443
rect 29963 6440 29975 6443
rect 30926 6440 30932 6452
rect 29963 6412 30932 6440
rect 29963 6409 29975 6412
rect 29917 6403 29975 6409
rect 30926 6400 30932 6412
rect 30984 6400 30990 6452
rect 33318 6400 33324 6452
rect 33376 6400 33382 6452
rect 33597 6443 33655 6449
rect 33597 6409 33609 6443
rect 33643 6440 33655 6443
rect 33870 6440 33876 6452
rect 33643 6412 33876 6440
rect 33643 6409 33655 6412
rect 33597 6403 33655 6409
rect 33870 6400 33876 6412
rect 33928 6400 33934 6452
rect 29825 6375 29883 6381
rect 29825 6341 29837 6375
rect 29871 6372 29883 6375
rect 30098 6372 30104 6384
rect 29871 6344 30104 6372
rect 29871 6341 29883 6344
rect 29825 6335 29883 6341
rect 30098 6332 30104 6344
rect 30156 6332 30162 6384
rect 31662 6372 31668 6384
rect 30576 6344 31668 6372
rect 30576 6316 30604 6344
rect 31662 6332 31668 6344
rect 31720 6372 31726 6384
rect 32217 6375 32275 6381
rect 32217 6372 32229 6375
rect 31720 6344 32229 6372
rect 31720 6332 31726 6344
rect 32217 6341 32229 6344
rect 32263 6341 32275 6375
rect 32217 6335 32275 6341
rect 32306 6332 32312 6384
rect 32364 6332 32370 6384
rect 34057 6375 34115 6381
rect 34057 6372 34069 6375
rect 33428 6344 34069 6372
rect 33428 6316 33456 6344
rect 34057 6341 34069 6344
rect 34103 6341 34115 6375
rect 34057 6335 34115 6341
rect 27709 6307 27767 6313
rect 27709 6273 27721 6307
rect 27755 6273 27767 6307
rect 27709 6267 27767 6273
rect 28077 6307 28135 6313
rect 28077 6273 28089 6307
rect 28123 6273 28135 6307
rect 28445 6307 28503 6313
rect 28445 6304 28457 6307
rect 28077 6267 28135 6273
rect 28184 6276 28457 6304
rect 25406 6196 25412 6248
rect 25464 6236 25470 6248
rect 27249 6239 27307 6245
rect 27249 6236 27261 6239
rect 25464 6208 27261 6236
rect 25464 6196 25470 6208
rect 27249 6205 27261 6208
rect 27295 6205 27307 6239
rect 27249 6199 27307 6205
rect 26142 6168 26148 6180
rect 25332 6140 26148 6168
rect 24949 6131 25007 6137
rect 11572 6072 12296 6100
rect 11572 6060 11578 6072
rect 12434 6060 12440 6112
rect 12492 6060 12498 6112
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 15286 6100 15292 6112
rect 14599 6072 15292 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 15378 6060 15384 6112
rect 15436 6060 15442 6112
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 15528 6072 15577 6100
rect 15528 6060 15534 6072
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 15565 6063 15623 6069
rect 17957 6103 18015 6109
rect 17957 6069 17969 6103
rect 18003 6100 18015 6103
rect 18966 6100 18972 6112
rect 18003 6072 18972 6100
rect 18003 6069 18015 6072
rect 17957 6063 18015 6069
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 21177 6103 21235 6109
rect 21177 6100 21189 6103
rect 20772 6072 21189 6100
rect 20772 6060 20778 6072
rect 21177 6069 21189 6072
rect 21223 6100 21235 6103
rect 21634 6100 21640 6112
rect 21223 6072 21640 6100
rect 21223 6069 21235 6072
rect 21177 6063 21235 6069
rect 21634 6060 21640 6072
rect 21692 6100 21698 6112
rect 22370 6100 22376 6112
rect 21692 6072 22376 6100
rect 21692 6060 21698 6072
rect 22370 6060 22376 6072
rect 22428 6060 22434 6112
rect 24213 6103 24271 6109
rect 24213 6069 24225 6103
rect 24259 6100 24271 6103
rect 24578 6100 24584 6112
rect 24259 6072 24584 6100
rect 24259 6069 24271 6072
rect 24213 6063 24271 6069
rect 24578 6060 24584 6072
rect 24636 6060 24642 6112
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 24964 6100 24992 6131
rect 26142 6128 26148 6140
rect 26200 6128 26206 6180
rect 26786 6128 26792 6180
rect 26844 6168 26850 6180
rect 28184 6168 28212 6276
rect 28445 6273 28457 6276
rect 28491 6304 28503 6307
rect 28626 6304 28632 6316
rect 28491 6276 28632 6304
rect 28491 6273 28503 6276
rect 28445 6267 28503 6273
rect 28626 6264 28632 6276
rect 28684 6264 28690 6316
rect 29181 6307 29239 6313
rect 29181 6273 29193 6307
rect 29227 6304 29239 6307
rect 29227 6276 29592 6304
rect 29227 6273 29239 6276
rect 29181 6267 29239 6273
rect 28902 6196 28908 6248
rect 28960 6236 28966 6248
rect 29273 6239 29331 6245
rect 29273 6236 29285 6239
rect 28960 6208 29285 6236
rect 28960 6196 28966 6208
rect 29273 6205 29285 6208
rect 29319 6205 29331 6239
rect 29564 6236 29592 6276
rect 29730 6264 29736 6316
rect 29788 6304 29794 6316
rect 30009 6307 30067 6313
rect 30009 6304 30021 6307
rect 29788 6276 30021 6304
rect 29788 6264 29794 6276
rect 30009 6273 30021 6276
rect 30055 6304 30067 6307
rect 30282 6304 30288 6316
rect 30055 6276 30288 6304
rect 30055 6273 30067 6276
rect 30009 6267 30067 6273
rect 30282 6264 30288 6276
rect 30340 6264 30346 6316
rect 30558 6264 30564 6316
rect 30616 6264 30622 6316
rect 30834 6264 30840 6316
rect 30892 6264 30898 6316
rect 30926 6264 30932 6316
rect 30984 6304 30990 6316
rect 31205 6307 31263 6313
rect 31205 6304 31217 6307
rect 30984 6276 31217 6304
rect 30984 6264 30990 6276
rect 31205 6273 31217 6276
rect 31251 6304 31263 6307
rect 31386 6304 31392 6316
rect 31251 6276 31392 6304
rect 31251 6273 31263 6276
rect 31205 6267 31263 6273
rect 31386 6264 31392 6276
rect 31444 6264 31450 6316
rect 32677 6307 32735 6313
rect 32677 6273 32689 6307
rect 32723 6273 32735 6307
rect 32677 6267 32735 6273
rect 32769 6307 32827 6313
rect 32769 6273 32781 6307
rect 32815 6304 32827 6307
rect 32858 6304 32864 6316
rect 32815 6276 32864 6304
rect 32815 6273 32827 6276
rect 32769 6267 32827 6273
rect 29914 6236 29920 6248
rect 29564 6208 29920 6236
rect 29273 6199 29331 6205
rect 29914 6196 29920 6208
rect 29972 6196 29978 6248
rect 30469 6239 30527 6245
rect 30469 6205 30481 6239
rect 30515 6236 30527 6239
rect 30742 6236 30748 6248
rect 30515 6208 30748 6236
rect 30515 6205 30527 6208
rect 30469 6199 30527 6205
rect 30742 6196 30748 6208
rect 30800 6196 30806 6248
rect 32214 6196 32220 6248
rect 32272 6236 32278 6248
rect 32692 6236 32720 6267
rect 32858 6264 32864 6276
rect 32916 6304 32922 6316
rect 33229 6307 33287 6313
rect 32916 6276 33180 6304
rect 32916 6264 32922 6276
rect 33152 6236 33180 6276
rect 33229 6273 33241 6307
rect 33275 6304 33287 6307
rect 33410 6304 33416 6316
rect 33275 6276 33416 6304
rect 33275 6273 33287 6276
rect 33229 6267 33287 6273
rect 33410 6264 33416 6276
rect 33468 6264 33474 6316
rect 33505 6307 33563 6313
rect 33505 6273 33517 6307
rect 33551 6304 33563 6307
rect 34606 6304 34612 6316
rect 33551 6276 34612 6304
rect 33551 6273 33563 6276
rect 33505 6267 33563 6273
rect 33520 6236 33548 6267
rect 34606 6264 34612 6276
rect 34664 6264 34670 6316
rect 32272 6208 32812 6236
rect 33152 6208 33548 6236
rect 32272 6196 32278 6208
rect 26844 6140 28212 6168
rect 26844 6128 26850 6140
rect 29638 6128 29644 6180
rect 29696 6168 29702 6180
rect 30193 6171 30251 6177
rect 30193 6168 30205 6171
rect 29696 6140 30205 6168
rect 29696 6128 29702 6140
rect 30193 6137 30205 6140
rect 30239 6168 30251 6171
rect 31478 6168 31484 6180
rect 30239 6140 31484 6168
rect 30239 6137 30251 6140
rect 30193 6131 30251 6137
rect 31478 6128 31484 6140
rect 31536 6128 31542 6180
rect 32784 6168 32812 6208
rect 34057 6171 34115 6177
rect 34057 6168 34069 6171
rect 32784 6140 34069 6168
rect 34057 6137 34069 6140
rect 34103 6168 34115 6171
rect 34238 6168 34244 6180
rect 34103 6140 34244 6168
rect 34103 6137 34115 6140
rect 34057 6131 34115 6137
rect 34238 6128 34244 6140
rect 34296 6128 34302 6180
rect 25682 6100 25688 6112
rect 24728 6072 25688 6100
rect 24728 6060 24734 6072
rect 25682 6060 25688 6072
rect 25740 6060 25746 6112
rect 26234 6060 26240 6112
rect 26292 6060 26298 6112
rect 26510 6060 26516 6112
rect 26568 6100 26574 6112
rect 28350 6100 28356 6112
rect 26568 6072 28356 6100
rect 26568 6060 26574 6072
rect 28350 6060 28356 6072
rect 28408 6060 28414 6112
rect 1104 6010 36432 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 36432 6010
rect 1104 5936 36432 5958
rect 5258 5856 5264 5908
rect 5316 5856 5322 5908
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 7340 5868 7573 5896
rect 7340 5856 7346 5868
rect 7561 5865 7573 5868
rect 7607 5865 7619 5899
rect 7561 5859 7619 5865
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 10836 5868 10885 5896
rect 10836 5856 10842 5868
rect 10873 5865 10885 5868
rect 10919 5865 10931 5899
rect 10873 5859 10931 5865
rect 12056 5899 12114 5905
rect 12056 5865 12068 5899
rect 12102 5896 12114 5899
rect 12434 5896 12440 5908
rect 12102 5868 12440 5896
rect 12102 5865 12114 5868
rect 12056 5859 12114 5865
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 16206 5856 16212 5908
rect 16264 5856 16270 5908
rect 16298 5856 16304 5908
rect 16356 5896 16362 5908
rect 17313 5899 17371 5905
rect 17313 5896 17325 5899
rect 16356 5868 17325 5896
rect 16356 5856 16362 5868
rect 17313 5865 17325 5868
rect 17359 5865 17371 5899
rect 17313 5859 17371 5865
rect 17497 5899 17555 5905
rect 17497 5865 17509 5899
rect 17543 5896 17555 5899
rect 20714 5896 20720 5908
rect 17543 5868 20720 5896
rect 17543 5865 17555 5868
rect 17497 5859 17555 5865
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 20809 5899 20867 5905
rect 20809 5865 20821 5899
rect 20855 5896 20867 5899
rect 20898 5896 20904 5908
rect 20855 5868 20904 5896
rect 20855 5865 20867 5868
rect 20809 5859 20867 5865
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 20993 5899 21051 5905
rect 20993 5865 21005 5899
rect 21039 5896 21051 5899
rect 21266 5896 21272 5908
rect 21039 5868 21272 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 21376 5868 22692 5896
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8168 5800 9720 5828
rect 8168 5788 8174 5800
rect 5626 5760 5632 5772
rect 5184 5732 5632 5760
rect 5184 5701 5212 5732
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 7098 5720 7104 5772
rect 7156 5760 7162 5772
rect 7156 5732 7788 5760
rect 7156 5720 7162 5732
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 5350 5652 5356 5704
rect 5408 5652 5414 5704
rect 6362 5652 6368 5704
rect 6420 5692 6426 5704
rect 7760 5701 7788 5732
rect 9582 5720 9588 5772
rect 9640 5720 9646 5772
rect 9692 5760 9720 5800
rect 9950 5788 9956 5840
rect 10008 5828 10014 5840
rect 10137 5831 10195 5837
rect 10137 5828 10149 5831
rect 10008 5800 10149 5828
rect 10008 5788 10014 5800
rect 10137 5797 10149 5800
rect 10183 5797 10195 5831
rect 10137 5791 10195 5797
rect 13817 5831 13875 5837
rect 13817 5797 13829 5831
rect 13863 5828 13875 5831
rect 13906 5828 13912 5840
rect 13863 5800 13912 5828
rect 13863 5797 13875 5800
rect 13817 5791 13875 5797
rect 13906 5788 13912 5800
rect 13964 5828 13970 5840
rect 21376 5828 21404 5868
rect 13964 5800 21404 5828
rect 21453 5831 21511 5837
rect 13964 5788 13970 5800
rect 21453 5797 21465 5831
rect 21499 5828 21511 5831
rect 22554 5828 22560 5840
rect 21499 5800 22560 5828
rect 21499 5797 21511 5800
rect 21453 5791 21511 5797
rect 22554 5788 22560 5800
rect 22612 5788 22618 5840
rect 22664 5828 22692 5868
rect 22738 5856 22744 5908
rect 22796 5896 22802 5908
rect 22833 5899 22891 5905
rect 22833 5896 22845 5899
rect 22796 5868 22845 5896
rect 22796 5856 22802 5868
rect 22833 5865 22845 5868
rect 22879 5865 22891 5899
rect 22833 5859 22891 5865
rect 24578 5856 24584 5908
rect 24636 5896 24642 5908
rect 25498 5896 25504 5908
rect 24636 5868 25504 5896
rect 24636 5856 24642 5868
rect 25498 5856 25504 5868
rect 25556 5856 25562 5908
rect 27893 5899 27951 5905
rect 27893 5896 27905 5899
rect 27172 5868 27905 5896
rect 26786 5828 26792 5840
rect 22664 5800 26792 5828
rect 26786 5788 26792 5800
rect 26844 5788 26850 5840
rect 27172 5828 27200 5868
rect 27893 5865 27905 5868
rect 27939 5896 27951 5899
rect 30374 5896 30380 5908
rect 27939 5868 30380 5896
rect 27939 5865 27951 5868
rect 27893 5859 27951 5865
rect 30374 5856 30380 5868
rect 30432 5856 30438 5908
rect 30558 5856 30564 5908
rect 30616 5896 30622 5908
rect 31113 5899 31171 5905
rect 31113 5896 31125 5899
rect 30616 5868 31125 5896
rect 30616 5856 30622 5868
rect 31113 5865 31125 5868
rect 31159 5865 31171 5899
rect 31113 5859 31171 5865
rect 31938 5856 31944 5908
rect 31996 5856 32002 5908
rect 27126 5800 27200 5828
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 9692 5732 11529 5760
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 11790 5720 11796 5772
rect 11848 5720 11854 5772
rect 12710 5720 12716 5772
rect 12768 5760 12774 5772
rect 19242 5760 19248 5772
rect 12768 5732 13768 5760
rect 12768 5720 12774 5732
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 6420 5664 7573 5692
rect 6420 5652 6426 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 8570 5652 8576 5704
rect 8628 5652 8634 5704
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 13740 5701 13768 5732
rect 13832 5732 19248 5760
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 9539 5664 10977 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10137 5627 10195 5633
rect 10137 5624 10149 5627
rect 10100 5596 10149 5624
rect 10100 5584 10106 5596
rect 10137 5593 10149 5596
rect 10183 5593 10195 5627
rect 10137 5587 10195 5593
rect 10597 5627 10655 5633
rect 10597 5593 10609 5627
rect 10643 5624 10655 5627
rect 10870 5624 10876 5636
rect 10643 5596 10876 5624
rect 10643 5593 10655 5596
rect 10597 5587 10655 5593
rect 10870 5584 10876 5596
rect 10928 5624 10934 5636
rect 11330 5624 11336 5636
rect 10928 5596 11336 5624
rect 10928 5584 10934 5596
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 11606 5584 11612 5636
rect 11664 5624 11670 5636
rect 12526 5624 12532 5636
rect 11664 5596 12532 5624
rect 11664 5584 11670 5596
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 13832 5624 13860 5732
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 24489 5763 24547 5769
rect 24489 5760 24501 5763
rect 19536 5732 20116 5760
rect 13998 5652 14004 5704
rect 14056 5692 14062 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 14056 5664 14105 5692
rect 14056 5652 14062 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 14792 5664 15025 5692
rect 14792 5652 14798 5664
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15194 5652 15200 5704
rect 15252 5652 15258 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 13464 5596 13860 5624
rect 15304 5624 15332 5655
rect 15470 5652 15476 5704
rect 15528 5652 15534 5704
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5692 15623 5695
rect 15654 5692 15660 5704
rect 15611 5664 15660 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 16209 5695 16267 5701
rect 16209 5661 16221 5695
rect 16255 5692 16267 5695
rect 16390 5692 16396 5704
rect 16255 5664 16396 5692
rect 16255 5661 16267 5664
rect 16209 5655 16267 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16482 5652 16488 5704
rect 16540 5652 16546 5704
rect 19426 5692 19432 5704
rect 17328 5664 19432 5692
rect 15838 5624 15844 5636
rect 15304 5596 15844 5624
rect 8386 5516 8392 5568
rect 8444 5556 8450 5568
rect 8662 5556 8668 5568
rect 8444 5528 8668 5556
rect 8444 5516 8450 5528
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 9033 5559 9091 5565
rect 9033 5525 9045 5559
rect 9079 5556 9091 5559
rect 9306 5556 9312 5568
rect 9079 5528 9312 5556
rect 9079 5525 9091 5528
rect 9033 5519 9091 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 10689 5559 10747 5565
rect 10689 5525 10701 5559
rect 10735 5556 10747 5559
rect 10778 5556 10784 5568
rect 10735 5528 10784 5556
rect 10735 5525 10747 5528
rect 10689 5519 10747 5525
rect 10778 5516 10784 5528
rect 10836 5556 10842 5568
rect 13464 5556 13492 5596
rect 15838 5584 15844 5596
rect 15896 5584 15902 5636
rect 17328 5624 17356 5664
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 16408 5596 17356 5624
rect 10836 5528 13492 5556
rect 10836 5516 10842 5528
rect 13538 5516 13544 5568
rect 13596 5516 13602 5568
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 14737 5559 14795 5565
rect 14737 5556 14749 5559
rect 14608 5528 14749 5556
rect 14608 5516 14614 5528
rect 14737 5525 14749 5528
rect 14783 5525 14795 5559
rect 14737 5519 14795 5525
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 16408 5565 16436 5596
rect 17402 5584 17408 5636
rect 17460 5633 17466 5636
rect 17460 5627 17523 5633
rect 17460 5593 17477 5627
rect 17511 5593 17523 5627
rect 17460 5587 17523 5593
rect 17681 5627 17739 5633
rect 17681 5593 17693 5627
rect 17727 5593 17739 5627
rect 17681 5587 17739 5593
rect 17460 5584 17466 5587
rect 16393 5559 16451 5565
rect 16393 5556 16405 5559
rect 15620 5528 16405 5556
rect 15620 5516 15626 5528
rect 16393 5525 16405 5528
rect 16439 5525 16451 5559
rect 17696 5556 17724 5587
rect 17954 5584 17960 5636
rect 18012 5624 18018 5636
rect 19536 5624 19564 5732
rect 19610 5652 19616 5704
rect 19668 5652 19674 5704
rect 19702 5652 19708 5704
rect 19760 5652 19766 5704
rect 19978 5701 19984 5704
rect 19935 5695 19984 5701
rect 19935 5661 19947 5695
rect 19981 5661 19984 5695
rect 19935 5655 19984 5661
rect 19978 5652 19984 5655
rect 20036 5652 20042 5704
rect 20088 5701 20116 5732
rect 21376 5732 24501 5760
rect 20073 5695 20131 5701
rect 20073 5661 20085 5695
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 18012 5596 19564 5624
rect 19797 5627 19855 5633
rect 18012 5584 18018 5596
rect 19797 5593 19809 5627
rect 19843 5593 19855 5627
rect 20088 5624 20116 5655
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 21376 5701 21404 5732
rect 24489 5729 24501 5732
rect 24535 5729 24547 5763
rect 24489 5723 24547 5729
rect 24670 5720 24676 5772
rect 24728 5720 24734 5772
rect 24857 5763 24915 5769
rect 24857 5729 24869 5763
rect 24903 5760 24915 5763
rect 25038 5760 25044 5772
rect 24903 5732 25044 5760
rect 24903 5729 24915 5732
rect 24857 5723 24915 5729
rect 21085 5695 21143 5701
rect 21085 5692 21097 5695
rect 20312 5664 21097 5692
rect 20312 5652 20318 5664
rect 21085 5661 21097 5664
rect 21131 5661 21143 5695
rect 21085 5655 21143 5661
rect 21361 5695 21419 5701
rect 21361 5661 21373 5695
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 20625 5627 20683 5633
rect 20625 5624 20637 5627
rect 20088 5596 20637 5624
rect 19797 5587 19855 5593
rect 20625 5593 20637 5596
rect 20671 5624 20683 5627
rect 20714 5624 20720 5636
rect 20671 5596 20720 5624
rect 20671 5593 20683 5596
rect 20625 5587 20683 5593
rect 18046 5556 18052 5568
rect 17696 5528 18052 5556
rect 16393 5519 16451 5525
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19429 5559 19487 5565
rect 19429 5556 19441 5559
rect 19392 5528 19441 5556
rect 19392 5516 19398 5528
rect 19429 5525 19441 5528
rect 19475 5525 19487 5559
rect 19429 5519 19487 5525
rect 19518 5516 19524 5568
rect 19576 5556 19582 5568
rect 19812 5556 19840 5587
rect 20714 5584 20720 5596
rect 20772 5584 20778 5636
rect 20841 5627 20899 5633
rect 20841 5593 20853 5627
rect 20887 5624 20899 5627
rect 21376 5624 21404 5655
rect 21542 5652 21548 5704
rect 21600 5652 21606 5704
rect 21634 5652 21640 5704
rect 21692 5652 21698 5704
rect 21818 5652 21824 5704
rect 21876 5652 21882 5704
rect 22830 5652 22836 5704
rect 22888 5652 22894 5704
rect 23385 5695 23443 5701
rect 23385 5661 23397 5695
rect 23431 5692 23443 5695
rect 23566 5692 23572 5704
rect 23431 5664 23572 5692
rect 23431 5661 23443 5664
rect 23385 5655 23443 5661
rect 23566 5652 23572 5664
rect 23624 5652 23630 5704
rect 23750 5652 23756 5704
rect 23808 5652 23814 5704
rect 24213 5695 24271 5701
rect 24213 5661 24225 5695
rect 24259 5661 24271 5695
rect 24213 5655 24271 5661
rect 20887 5596 21404 5624
rect 20887 5593 20899 5596
rect 20841 5587 20899 5593
rect 19576 5528 19840 5556
rect 21560 5556 21588 5652
rect 24228 5624 24256 5655
rect 24578 5652 24584 5704
rect 24636 5692 24642 5704
rect 24765 5695 24823 5701
rect 24765 5692 24777 5695
rect 24636 5664 24777 5692
rect 24636 5652 24642 5664
rect 24765 5661 24777 5664
rect 24811 5661 24823 5695
rect 24765 5655 24823 5661
rect 24872 5624 24900 5723
rect 25038 5720 25044 5732
rect 25096 5760 25102 5772
rect 26421 5763 26479 5769
rect 26421 5760 26433 5763
rect 25096 5732 26433 5760
rect 25096 5720 25102 5732
rect 26421 5729 26433 5732
rect 26467 5729 26479 5763
rect 27126 5760 27154 5800
rect 27246 5788 27252 5840
rect 27304 5828 27310 5840
rect 27982 5828 27988 5840
rect 27304 5800 27988 5828
rect 27304 5788 27310 5800
rect 27982 5788 27988 5800
rect 28040 5828 28046 5840
rect 30190 5828 30196 5840
rect 28040 5800 29040 5828
rect 28040 5788 28046 5800
rect 28445 5763 28503 5769
rect 28445 5760 28457 5763
rect 26421 5723 26479 5729
rect 27080 5732 27154 5760
rect 27816 5732 28457 5760
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5692 25007 5695
rect 26142 5692 26148 5704
rect 24995 5664 26148 5692
rect 24995 5661 25007 5664
rect 24949 5655 25007 5661
rect 26142 5652 26148 5664
rect 26200 5692 26206 5704
rect 26881 5695 26939 5701
rect 26881 5692 26893 5695
rect 26200 5664 26893 5692
rect 26200 5652 26206 5664
rect 26881 5661 26893 5664
rect 26927 5661 26939 5695
rect 26881 5655 26939 5661
rect 24228 5596 24900 5624
rect 26513 5627 26571 5633
rect 26513 5593 26525 5627
rect 26559 5593 26571 5627
rect 26513 5587 26571 5593
rect 23934 5556 23940 5568
rect 21560 5528 23940 5556
rect 19576 5516 19582 5528
rect 23934 5516 23940 5528
rect 23992 5516 23998 5568
rect 26326 5516 26332 5568
rect 26384 5556 26390 5568
rect 26528 5556 26556 5587
rect 26384 5528 26556 5556
rect 26896 5556 26924 5655
rect 26970 5652 26976 5704
rect 27028 5652 27034 5704
rect 27080 5701 27108 5732
rect 27816 5701 27844 5732
rect 28445 5729 28457 5732
rect 28491 5760 28503 5763
rect 28902 5760 28908 5772
rect 28491 5732 28908 5760
rect 28491 5729 28503 5732
rect 28445 5723 28503 5729
rect 28902 5720 28908 5732
rect 28960 5720 28966 5772
rect 29012 5760 29040 5800
rect 29840 5800 30196 5828
rect 29730 5760 29736 5772
rect 29012 5732 29736 5760
rect 27065 5695 27123 5701
rect 27065 5661 27077 5695
rect 27111 5661 27123 5695
rect 27065 5655 27123 5661
rect 27433 5695 27491 5701
rect 27433 5661 27445 5695
rect 27479 5661 27491 5695
rect 27433 5655 27491 5661
rect 27801 5695 27859 5701
rect 27801 5661 27813 5695
rect 27847 5661 27859 5695
rect 27801 5655 27859 5661
rect 27448 5624 27476 5655
rect 27982 5652 27988 5704
rect 28040 5652 28046 5704
rect 28813 5695 28871 5701
rect 28092 5664 28580 5692
rect 28092 5624 28120 5664
rect 28350 5633 28356 5636
rect 27080 5596 28120 5624
rect 28328 5627 28356 5633
rect 27080 5556 27108 5596
rect 28328 5593 28340 5627
rect 28328 5587 28356 5593
rect 28350 5584 28356 5587
rect 28408 5584 28414 5636
rect 28552 5633 28580 5664
rect 28813 5661 28825 5695
rect 28859 5692 28871 5695
rect 29012 5692 29040 5732
rect 29730 5720 29736 5732
rect 29788 5720 29794 5772
rect 29840 5769 29868 5800
rect 30190 5788 30196 5800
rect 30248 5788 30254 5840
rect 30650 5788 30656 5840
rect 30708 5788 30714 5840
rect 30834 5788 30840 5840
rect 30892 5828 30898 5840
rect 31021 5831 31079 5837
rect 31021 5828 31033 5831
rect 30892 5800 31033 5828
rect 30892 5788 30898 5800
rect 31021 5797 31033 5800
rect 31067 5797 31079 5831
rect 31021 5791 31079 5797
rect 29825 5763 29883 5769
rect 29825 5729 29837 5763
rect 29871 5729 29883 5763
rect 30852 5760 30880 5788
rect 29825 5723 29883 5729
rect 30208 5732 30880 5760
rect 28859 5664 29040 5692
rect 28859 5661 28871 5664
rect 28813 5655 28871 5661
rect 29638 5652 29644 5704
rect 29696 5652 29702 5704
rect 30208 5701 30236 5732
rect 30926 5720 30932 5772
rect 30984 5720 30990 5772
rect 31036 5760 31064 5791
rect 31478 5788 31484 5840
rect 31536 5788 31542 5840
rect 32122 5760 32128 5772
rect 31036 5732 31708 5760
rect 30193 5695 30251 5701
rect 30193 5661 30205 5695
rect 30239 5661 30251 5695
rect 30193 5655 30251 5661
rect 30285 5695 30343 5701
rect 30285 5661 30297 5695
rect 30331 5692 30343 5695
rect 30558 5692 30564 5704
rect 30331 5664 30564 5692
rect 30331 5661 30343 5664
rect 30285 5655 30343 5661
rect 30558 5652 30564 5664
rect 30616 5652 30622 5704
rect 28537 5627 28595 5633
rect 28537 5593 28549 5627
rect 28583 5624 28595 5627
rect 30098 5624 30104 5636
rect 28583 5596 30104 5624
rect 28583 5593 28595 5596
rect 28537 5587 28595 5593
rect 30098 5584 30104 5596
rect 30156 5584 30162 5636
rect 30377 5627 30435 5633
rect 30377 5593 30389 5627
rect 30423 5624 30435 5627
rect 30944 5624 30972 5720
rect 31573 5695 31631 5701
rect 31573 5661 31585 5695
rect 31619 5661 31631 5695
rect 31573 5655 31631 5661
rect 30423 5596 30972 5624
rect 30423 5593 30435 5596
rect 30377 5587 30435 5593
rect 26896 5528 27108 5556
rect 26384 5516 26390 5528
rect 27338 5516 27344 5568
rect 27396 5556 27402 5568
rect 27617 5559 27675 5565
rect 27617 5556 27629 5559
rect 27396 5528 27629 5556
rect 27396 5516 27402 5528
rect 27617 5525 27629 5528
rect 27663 5525 27675 5559
rect 27617 5519 27675 5525
rect 28166 5516 28172 5568
rect 28224 5516 28230 5568
rect 29546 5516 29552 5568
rect 29604 5556 29610 5568
rect 31588 5556 31616 5655
rect 31680 5624 31708 5732
rect 31772 5732 32128 5760
rect 31772 5701 31800 5732
rect 32122 5720 32128 5732
rect 32180 5760 32186 5772
rect 32401 5763 32459 5769
rect 32401 5760 32413 5763
rect 32180 5732 32413 5760
rect 32180 5720 32186 5732
rect 32401 5729 32413 5732
rect 32447 5729 32459 5763
rect 32401 5723 32459 5729
rect 31757 5695 31815 5701
rect 31757 5661 31769 5695
rect 31803 5661 31815 5695
rect 31757 5655 31815 5661
rect 32214 5652 32220 5704
rect 32272 5652 32278 5704
rect 32858 5652 32864 5704
rect 32916 5652 32922 5704
rect 32953 5695 33011 5701
rect 32953 5661 32965 5695
rect 32999 5692 33011 5695
rect 33870 5692 33876 5704
rect 32999 5664 33876 5692
rect 32999 5661 33011 5664
rect 32953 5655 33011 5661
rect 33870 5652 33876 5664
rect 33928 5652 33934 5704
rect 32769 5627 32827 5633
rect 32769 5624 32781 5627
rect 31680 5596 32781 5624
rect 32769 5593 32781 5596
rect 32815 5624 32827 5627
rect 33410 5624 33416 5636
rect 32815 5596 33416 5624
rect 32815 5593 32827 5596
rect 32769 5587 32827 5593
rect 33410 5584 33416 5596
rect 33468 5584 33474 5636
rect 29604 5528 31616 5556
rect 29604 5516 29610 5528
rect 1104 5466 36432 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 36432 5466
rect 1104 5392 36432 5414
rect 8110 5312 8116 5364
rect 8168 5312 8174 5364
rect 11698 5352 11704 5364
rect 10244 5324 11704 5352
rect 7742 5244 7748 5296
rect 7800 5284 7806 5296
rect 7800 5270 8418 5284
rect 7800 5256 8432 5270
rect 7800 5244 7806 5256
rect 8404 5148 8432 5256
rect 9306 5244 9312 5296
rect 9364 5284 9370 5296
rect 10244 5293 10272 5324
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 11848 5324 14320 5352
rect 11848 5312 11854 5324
rect 9585 5287 9643 5293
rect 9585 5284 9597 5287
rect 9364 5256 9597 5284
rect 9364 5244 9370 5256
rect 9585 5253 9597 5256
rect 9631 5253 9643 5287
rect 10229 5287 10287 5293
rect 10229 5284 10241 5287
rect 9585 5247 9643 5253
rect 9876 5256 10241 5284
rect 9876 5225 9904 5256
rect 10229 5253 10241 5256
rect 10275 5253 10287 5287
rect 10229 5247 10287 5253
rect 11054 5244 11060 5296
rect 11112 5244 11118 5296
rect 11238 5244 11244 5296
rect 11296 5244 11302 5296
rect 11882 5284 11888 5296
rect 11532 5256 11888 5284
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10192 5188 10977 5216
rect 10192 5176 10198 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 11256 5216 11284 5244
rect 10965 5179 11023 5185
rect 11072 5188 11284 5216
rect 10226 5148 10232 5160
rect 8404 5120 10232 5148
rect 9876 5092 9904 5120
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 9858 5040 9864 5092
rect 9916 5040 9922 5092
rect 10980 5080 11008 5179
rect 11072 5157 11100 5188
rect 11330 5176 11336 5228
rect 11388 5176 11394 5228
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 11532 5225 11560 5256
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 12802 5244 12808 5296
rect 12860 5244 12866 5296
rect 13078 5244 13084 5296
rect 13136 5284 13142 5296
rect 14182 5284 14188 5296
rect 13136 5256 14188 5284
rect 13136 5244 13142 5256
rect 14182 5244 14188 5256
rect 14240 5244 14246 5296
rect 14292 5293 14320 5324
rect 19150 5312 19156 5364
rect 19208 5352 19214 5364
rect 19521 5355 19579 5361
rect 19521 5352 19533 5355
rect 19208 5324 19533 5352
rect 19208 5312 19214 5324
rect 19521 5321 19533 5324
rect 19567 5321 19579 5355
rect 19521 5315 19579 5321
rect 22002 5312 22008 5364
rect 22060 5352 22066 5364
rect 24302 5352 24308 5364
rect 22060 5324 24308 5352
rect 22060 5312 22066 5324
rect 14274 5287 14332 5293
rect 14274 5253 14286 5287
rect 14320 5253 14332 5287
rect 14274 5247 14332 5253
rect 14366 5244 14372 5296
rect 14424 5284 14430 5296
rect 15654 5284 15660 5296
rect 14424 5256 15660 5284
rect 14424 5244 14430 5256
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 19242 5244 19248 5296
rect 19300 5284 19306 5296
rect 19673 5287 19731 5293
rect 19673 5284 19685 5287
rect 19300 5256 19685 5284
rect 19300 5244 19306 5256
rect 19673 5253 19685 5256
rect 19719 5253 19731 5287
rect 19673 5247 19731 5253
rect 19889 5287 19947 5293
rect 19889 5253 19901 5287
rect 19935 5284 19947 5287
rect 21726 5284 21732 5296
rect 19935 5256 21732 5284
rect 19935 5253 19947 5256
rect 19889 5247 19947 5253
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11480 5188 11529 5216
rect 11480 5176 11486 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 15197 5219 15255 5225
rect 15197 5216 15209 5219
rect 11517 5179 11575 5185
rect 13832 5188 15209 5216
rect 13832 5160 13860 5188
rect 15197 5185 15209 5188
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 19061 5219 19119 5225
rect 19061 5216 19073 5219
rect 18564 5188 19073 5216
rect 18564 5176 18570 5188
rect 19061 5185 19073 5188
rect 19107 5185 19119 5219
rect 19061 5179 19119 5185
rect 19150 5176 19156 5228
rect 19208 5176 19214 5228
rect 11057 5151 11115 5157
rect 11057 5117 11069 5151
rect 11103 5117 11115 5151
rect 11057 5111 11115 5117
rect 11238 5108 11244 5160
rect 11296 5148 11302 5160
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 11296 5120 11805 5148
rect 11296 5108 11302 5120
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 11882 5108 11888 5160
rect 11940 5148 11946 5160
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 11940 5120 13461 5148
rect 11940 5108 11946 5120
rect 13449 5117 13461 5120
rect 13495 5148 13507 5151
rect 13814 5148 13820 5160
rect 13495 5120 13820 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 15010 5108 15016 5160
rect 15068 5108 15074 5160
rect 15286 5108 15292 5160
rect 15344 5148 15350 5160
rect 19904 5148 19932 5247
rect 21726 5244 21732 5256
rect 21784 5244 21790 5296
rect 22112 5293 22140 5324
rect 24302 5312 24308 5324
rect 24360 5312 24366 5364
rect 22097 5287 22155 5293
rect 22097 5253 22109 5287
rect 22143 5253 22155 5287
rect 22097 5247 22155 5253
rect 21174 5176 21180 5228
rect 21232 5216 21238 5228
rect 21913 5219 21971 5225
rect 21913 5216 21925 5219
rect 21232 5188 21925 5216
rect 21232 5176 21238 5188
rect 21913 5185 21925 5188
rect 21959 5185 21971 5219
rect 21913 5179 21971 5185
rect 22186 5176 22192 5228
rect 22244 5176 22250 5228
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 22462 5216 22468 5228
rect 22327 5188 22468 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 22925 5219 22983 5225
rect 22925 5185 22937 5219
rect 22971 5216 22983 5219
rect 24026 5216 24032 5228
rect 22971 5188 24032 5216
rect 22971 5185 22983 5188
rect 22925 5179 22983 5185
rect 24026 5176 24032 5188
rect 24084 5176 24090 5228
rect 26878 5176 26884 5228
rect 26936 5216 26942 5228
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 26936 5188 27169 5216
rect 26936 5176 26942 5188
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5216 27399 5219
rect 27430 5216 27436 5228
rect 27387 5188 27436 5216
rect 27387 5185 27399 5188
rect 27341 5179 27399 5185
rect 27430 5176 27436 5188
rect 27488 5216 27494 5228
rect 29822 5216 29828 5228
rect 27488 5188 29828 5216
rect 27488 5176 27494 5188
rect 29822 5176 29828 5188
rect 29880 5216 29886 5228
rect 30193 5219 30251 5225
rect 30193 5216 30205 5219
rect 29880 5188 30205 5216
rect 29880 5176 29886 5188
rect 30193 5185 30205 5188
rect 30239 5185 30251 5219
rect 30193 5179 30251 5185
rect 30377 5219 30435 5225
rect 30377 5185 30389 5219
rect 30423 5216 30435 5219
rect 30650 5216 30656 5228
rect 30423 5188 30656 5216
rect 30423 5185 30435 5188
rect 30377 5179 30435 5185
rect 30650 5176 30656 5188
rect 30708 5176 30714 5228
rect 15344 5120 19932 5148
rect 15344 5108 15350 5120
rect 13906 5080 13912 5092
rect 10980 5052 11652 5080
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 11241 5015 11299 5021
rect 11241 5012 11253 5015
rect 10836 4984 11253 5012
rect 10836 4972 10842 4984
rect 11241 4981 11253 4984
rect 11287 4981 11299 5015
rect 11624 5012 11652 5052
rect 12912 5052 13912 5080
rect 11790 5012 11796 5024
rect 11624 4984 11796 5012
rect 11241 4975 11299 4981
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12912 5012 12940 5052
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 19429 5083 19487 5089
rect 19429 5049 19441 5083
rect 19475 5080 19487 5083
rect 20162 5080 20168 5092
rect 19475 5052 20168 5080
rect 19475 5049 19487 5052
rect 19429 5043 19487 5049
rect 20162 5040 20168 5052
rect 20220 5040 20226 5092
rect 21082 5040 21088 5092
rect 21140 5080 21146 5092
rect 21634 5080 21640 5092
rect 21140 5052 21640 5080
rect 21140 5040 21146 5052
rect 21634 5040 21640 5052
rect 21692 5080 21698 5092
rect 22649 5083 22707 5089
rect 22649 5080 22661 5083
rect 21692 5052 22661 5080
rect 21692 5040 21698 5052
rect 22649 5049 22661 5052
rect 22695 5049 22707 5083
rect 22649 5043 22707 5049
rect 30374 5040 30380 5092
rect 30432 5040 30438 5092
rect 11940 4984 12940 5012
rect 11940 4972 11946 4984
rect 12986 4972 12992 5024
rect 13044 5012 13050 5024
rect 13265 5015 13323 5021
rect 13265 5012 13277 5015
rect 13044 4984 13277 5012
rect 13044 4972 13050 4984
rect 13265 4981 13277 4984
rect 13311 5012 13323 5015
rect 13538 5012 13544 5024
rect 13311 4984 13544 5012
rect 13311 4981 13323 4984
rect 13265 4975 13323 4981
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 14366 4972 14372 5024
rect 14424 4972 14430 5024
rect 19245 5015 19303 5021
rect 19245 4981 19257 5015
rect 19291 5012 19303 5015
rect 19334 5012 19340 5024
rect 19291 4984 19340 5012
rect 19291 4981 19303 4984
rect 19245 4975 19303 4981
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 19702 4972 19708 5024
rect 19760 4972 19766 5024
rect 22465 5015 22523 5021
rect 22465 4981 22477 5015
rect 22511 5012 22523 5015
rect 22554 5012 22560 5024
rect 22511 4984 22560 5012
rect 22511 4981 22523 4984
rect 22465 4975 22523 4981
rect 22554 4972 22560 4984
rect 22612 4972 22618 5024
rect 26970 4972 26976 5024
rect 27028 4972 27034 5024
rect 27338 4972 27344 5024
rect 27396 4972 27402 5024
rect 1104 4922 36432 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 36432 4922
rect 1104 4848 36432 4870
rect 11238 4768 11244 4820
rect 11296 4808 11302 4820
rect 11517 4811 11575 4817
rect 11517 4808 11529 4811
rect 11296 4780 11529 4808
rect 11296 4768 11302 4780
rect 11517 4777 11529 4780
rect 11563 4777 11575 4811
rect 11517 4771 11575 4777
rect 11606 4768 11612 4820
rect 11664 4808 11670 4820
rect 11701 4811 11759 4817
rect 11701 4808 11713 4811
rect 11664 4780 11713 4808
rect 11664 4768 11670 4780
rect 11701 4777 11713 4780
rect 11747 4777 11759 4811
rect 15286 4808 15292 4820
rect 11701 4771 11759 4777
rect 13188 4780 15292 4808
rect 10980 4712 11284 4740
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9950 4672 9956 4684
rect 8803 4644 9956 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10980 4681 11008 4712
rect 11256 4684 11284 4712
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11882 4740 11888 4752
rect 11388 4712 11888 4740
rect 11388 4700 11394 4712
rect 11882 4700 11888 4712
rect 11940 4700 11946 4752
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 11146 4672 11152 4684
rect 11103 4644 11152 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 11238 4632 11244 4684
rect 11296 4632 11302 4684
rect 12158 4672 12164 4684
rect 11808 4644 12164 4672
rect 11808 4616 11836 4644
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12342 4632 12348 4684
rect 12400 4672 12406 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 12400 4644 12449 4672
rect 12400 4632 12406 4644
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 12437 4635 12495 4641
rect 8018 4564 8024 4616
rect 8076 4604 8082 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 8076 4576 8125 4604
rect 8076 4564 8082 4576
rect 8113 4573 8125 4576
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 11698 4604 11704 4616
rect 10735 4576 11704 4604
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 8128 4468 8156 4567
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11790 4564 11796 4616
rect 11848 4564 11854 4616
rect 12066 4564 12072 4616
rect 12124 4604 12130 4616
rect 13188 4613 13216 4780
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 15654 4768 15660 4820
rect 15712 4808 15718 4820
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 15712 4780 16313 4808
rect 15712 4768 15718 4780
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 16301 4771 16359 4777
rect 17402 4768 17408 4820
rect 17460 4808 17466 4820
rect 17460 4780 18460 4808
rect 17460 4768 17466 4780
rect 14366 4740 14372 4752
rect 13280 4712 14372 4740
rect 13280 4681 13308 4712
rect 14366 4700 14372 4712
rect 14424 4700 14430 4752
rect 14645 4743 14703 4749
rect 14645 4709 14657 4743
rect 14691 4740 14703 4743
rect 15930 4740 15936 4752
rect 14691 4712 15936 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 15930 4700 15936 4712
rect 15988 4700 15994 4752
rect 17494 4740 17500 4752
rect 16592 4712 17500 4740
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 13354 4632 13360 4684
rect 13412 4632 13418 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 14384 4644 15485 4672
rect 12253 4607 12311 4613
rect 12253 4604 12265 4607
rect 12124 4576 12265 4604
rect 12124 4564 12130 4576
rect 12253 4573 12265 4576
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 13630 4564 13636 4616
rect 13688 4564 13694 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 14384 4613 14412 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 15473 4635 15531 4641
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 15804 4644 16160 4672
rect 15804 4632 15810 4644
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 14737 4607 14795 4613
rect 14737 4604 14749 4607
rect 14369 4567 14427 4573
rect 14476 4576 14749 4604
rect 9858 4496 9864 4548
rect 9916 4496 9922 4548
rect 10134 4496 10140 4548
rect 10192 4536 10198 4548
rect 10413 4539 10471 4545
rect 10413 4536 10425 4539
rect 10192 4508 10425 4536
rect 10192 4496 10198 4508
rect 10413 4505 10425 4508
rect 10459 4505 10471 4539
rect 10413 4499 10471 4505
rect 10962 4496 10968 4548
rect 11020 4536 11026 4548
rect 14292 4536 14320 4564
rect 14476 4536 14504 4576
rect 14737 4573 14749 4576
rect 14783 4573 14795 4607
rect 15838 4604 15844 4616
rect 14737 4567 14795 4573
rect 15304 4576 15844 4604
rect 11020 4508 13860 4536
rect 14292 4508 14504 4536
rect 14645 4539 14703 4545
rect 11020 4496 11026 4508
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 8128 4440 8953 4468
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 8941 4431 8999 4437
rect 11149 4471 11207 4477
rect 11149 4437 11161 4471
rect 11195 4468 11207 4471
rect 11790 4468 11796 4480
rect 11195 4440 11796 4468
rect 11195 4437 11207 4440
rect 11149 4431 11207 4437
rect 11790 4428 11796 4440
rect 11848 4428 11854 4480
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 11974 4468 11980 4480
rect 11931 4440 11980 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 12342 4428 12348 4480
rect 12400 4428 12406 4480
rect 12802 4428 12808 4480
rect 12860 4428 12866 4480
rect 13832 4477 13860 4508
rect 14645 4505 14657 4539
rect 14691 4536 14703 4539
rect 15304 4536 15332 4576
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 16022 4564 16028 4616
rect 16080 4564 16086 4616
rect 16132 4604 16160 4644
rect 16592 4613 16620 4712
rect 17494 4700 17500 4712
rect 17552 4700 17558 4752
rect 17865 4743 17923 4749
rect 17865 4709 17877 4743
rect 17911 4740 17923 4743
rect 18230 4740 18236 4752
rect 17911 4712 18236 4740
rect 17911 4709 17923 4712
rect 17865 4703 17923 4709
rect 18230 4700 18236 4712
rect 18288 4700 18294 4752
rect 18432 4740 18460 4780
rect 18506 4768 18512 4820
rect 18564 4768 18570 4820
rect 20714 4768 20720 4820
rect 20772 4808 20778 4820
rect 21082 4808 21088 4820
rect 20772 4780 21088 4808
rect 20772 4768 20778 4780
rect 21082 4768 21088 4780
rect 21140 4808 21146 4820
rect 21453 4811 21511 4817
rect 21453 4808 21465 4811
rect 21140 4780 21465 4808
rect 21140 4768 21146 4780
rect 21453 4777 21465 4780
rect 21499 4808 21511 4811
rect 22186 4808 22192 4820
rect 21499 4780 22192 4808
rect 21499 4777 21511 4780
rect 21453 4771 21511 4777
rect 22186 4768 22192 4780
rect 22244 4768 22250 4820
rect 23106 4768 23112 4820
rect 23164 4808 23170 4820
rect 23937 4811 23995 4817
rect 23937 4808 23949 4811
rect 23164 4780 23949 4808
rect 23164 4768 23170 4780
rect 23937 4777 23949 4780
rect 23983 4808 23995 4811
rect 24394 4808 24400 4820
rect 23983 4780 24400 4808
rect 23983 4777 23995 4780
rect 23937 4771 23995 4777
rect 24394 4768 24400 4780
rect 24452 4768 24458 4820
rect 25406 4768 25412 4820
rect 25464 4808 25470 4820
rect 34514 4808 34520 4820
rect 25464 4780 34520 4808
rect 25464 4768 25470 4780
rect 34514 4768 34520 4780
rect 34572 4768 34578 4820
rect 21266 4740 21272 4752
rect 18432 4712 21272 4740
rect 21266 4700 21272 4712
rect 21324 4700 21330 4752
rect 21358 4700 21364 4752
rect 21416 4740 21422 4752
rect 21726 4740 21732 4752
rect 21416 4712 21732 4740
rect 21416 4700 21422 4712
rect 21726 4700 21732 4712
rect 21784 4740 21790 4752
rect 23201 4743 23259 4749
rect 23201 4740 23213 4743
rect 21784 4712 23213 4740
rect 21784 4700 21790 4712
rect 23201 4709 23213 4712
rect 23247 4709 23259 4743
rect 23201 4703 23259 4709
rect 17034 4632 17040 4684
rect 17092 4672 17098 4684
rect 17092 4644 18184 4672
rect 17092 4632 17098 4644
rect 16577 4607 16635 4613
rect 16132 4576 16528 4604
rect 14691 4508 15332 4536
rect 15381 4539 15439 4545
rect 14691 4505 14703 4508
rect 14645 4499 14703 4505
rect 15381 4505 15393 4539
rect 15427 4536 15439 4539
rect 16114 4536 16120 4548
rect 15427 4508 16120 4536
rect 15427 4505 15439 4508
rect 15381 4499 15439 4505
rect 16114 4496 16120 4508
rect 16172 4496 16178 4548
rect 16500 4536 16528 4576
rect 16577 4573 16589 4607
rect 16623 4573 16635 4607
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 16577 4567 16635 4573
rect 16684 4576 17601 4604
rect 16684 4536 16712 4576
rect 17589 4573 17601 4576
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 17954 4564 17960 4616
rect 18012 4564 18018 4616
rect 18156 4613 18184 4644
rect 22646 4632 22652 4684
rect 22704 4632 22710 4684
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 18414 4604 18420 4616
rect 18371 4576 18420 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 21634 4564 21640 4616
rect 21692 4564 21698 4616
rect 21818 4564 21824 4616
rect 21876 4564 21882 4616
rect 22278 4564 22284 4616
rect 22336 4564 22342 4616
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4604 23075 4607
rect 23934 4604 23940 4616
rect 23063 4576 23940 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 23934 4564 23940 4576
rect 23992 4564 23998 4616
rect 16500 4508 16712 4536
rect 16850 4496 16856 4548
rect 16908 4536 16914 4548
rect 17129 4539 17187 4545
rect 17129 4536 17141 4539
rect 16908 4508 17141 4536
rect 16908 4496 16914 4508
rect 17129 4505 17141 4508
rect 17175 4505 17187 4539
rect 17129 4499 17187 4505
rect 17313 4539 17371 4545
rect 17313 4505 17325 4539
rect 17359 4536 17371 4539
rect 17402 4536 17408 4548
rect 17359 4508 17408 4536
rect 17359 4505 17371 4508
rect 17313 4499 17371 4505
rect 13817 4471 13875 4477
rect 13817 4437 13829 4471
rect 13863 4437 13875 4471
rect 13817 4431 13875 4437
rect 14185 4471 14243 4477
rect 14185 4437 14197 4471
rect 14231 4468 14243 4471
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 14231 4440 14473 4468
rect 14231 4437 14243 4440
rect 14185 4431 14243 4437
rect 14461 4437 14473 4440
rect 14507 4468 14519 4471
rect 16206 4468 16212 4480
rect 14507 4440 16212 4468
rect 14507 4437 14519 4440
rect 14461 4431 14519 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 17144 4468 17172 4499
rect 17402 4496 17408 4508
rect 17460 4496 17466 4548
rect 17865 4539 17923 4545
rect 17604 4508 17816 4536
rect 17604 4468 17632 4508
rect 17144 4440 17632 4468
rect 17678 4428 17684 4480
rect 17736 4428 17742 4480
rect 17788 4468 17816 4508
rect 17865 4505 17877 4539
rect 17911 4536 17923 4539
rect 18046 4536 18052 4548
rect 17911 4508 18052 4536
rect 17911 4505 17923 4508
rect 17865 4499 17923 4505
rect 18046 4496 18052 4508
rect 18104 4496 18110 4548
rect 18233 4539 18291 4545
rect 18233 4505 18245 4539
rect 18279 4536 18291 4539
rect 21358 4536 21364 4548
rect 18279 4508 21364 4536
rect 18279 4505 18291 4508
rect 18233 4499 18291 4505
rect 21358 4496 21364 4508
rect 21416 4496 21422 4548
rect 23842 4496 23848 4548
rect 23900 4496 23906 4548
rect 21821 4471 21879 4477
rect 21821 4468 21833 4471
rect 17788 4440 21833 4468
rect 21821 4437 21833 4440
rect 21867 4437 21879 4471
rect 21821 4431 21879 4437
rect 1104 4378 36432 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 36432 4378
rect 1104 4304 36432 4326
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 10689 4267 10747 4273
rect 10689 4264 10701 4267
rect 9824 4236 10701 4264
rect 9824 4224 9830 4236
rect 10689 4233 10701 4236
rect 10735 4233 10747 4267
rect 10689 4227 10747 4233
rect 10778 4224 10784 4276
rect 10836 4264 10842 4276
rect 13630 4264 13636 4276
rect 10836 4236 13636 4264
rect 10836 4224 10842 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 15565 4267 15623 4273
rect 15565 4233 15577 4267
rect 15611 4264 15623 4267
rect 16022 4264 16028 4276
rect 15611 4236 16028 4264
rect 15611 4233 15623 4236
rect 15565 4227 15623 4233
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 18414 4224 18420 4276
rect 18472 4224 18478 4276
rect 21637 4267 21695 4273
rect 21637 4233 21649 4267
rect 21683 4233 21695 4267
rect 21637 4227 21695 4233
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 9861 4199 9919 4205
rect 9861 4196 9873 4199
rect 9732 4168 9873 4196
rect 9732 4156 9738 4168
rect 9861 4165 9873 4168
rect 9907 4165 9919 4199
rect 12158 4196 12164 4208
rect 9861 4159 9919 4165
rect 11624 4168 12164 4196
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10152 4100 11008 4128
rect 8662 4020 8668 4072
rect 8720 4020 8726 4072
rect 8846 4020 8852 4072
rect 8904 4020 8910 4072
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 9582 4060 9588 4072
rect 9272 4032 9588 4060
rect 9272 4020 9278 4032
rect 9582 4020 9588 4032
rect 9640 4060 9646 4072
rect 10152 4069 10180 4100
rect 10980 4069 11008 4100
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11112 4100 11529 4128
rect 11112 4088 11118 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9640 4032 10149 4060
rect 9640 4020 9646 4032
rect 10137 4029 10149 4032
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11238 4060 11244 4072
rect 11011 4032 11244 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 9401 3995 9459 4001
rect 9401 3961 9413 3995
rect 9447 3992 9459 3995
rect 10796 3992 10824 4023
rect 11238 4020 11244 4032
rect 11296 4060 11302 4072
rect 11624 4060 11652 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 12710 4156 12716 4208
rect 12768 4156 12774 4208
rect 13446 4156 13452 4208
rect 13504 4196 13510 4208
rect 14366 4196 14372 4208
rect 13504 4168 14372 4196
rect 13504 4156 13510 4168
rect 14366 4156 14372 4168
rect 14424 4196 14430 4208
rect 21652 4196 21680 4227
rect 14424 4168 14582 4196
rect 15856 4168 16436 4196
rect 14424 4156 14430 4168
rect 15856 4140 15884 4168
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 11756 4100 11805 4128
rect 11756 4088 11762 4100
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 13814 4088 13820 4140
rect 13872 4088 13878 4140
rect 15838 4088 15844 4140
rect 15896 4088 15902 4140
rect 16114 4088 16120 4140
rect 16172 4088 16178 4140
rect 16206 4088 16212 4140
rect 16264 4128 16270 4140
rect 16301 4131 16359 4137
rect 16301 4128 16313 4131
rect 16264 4100 16313 4128
rect 16264 4088 16270 4100
rect 16301 4097 16313 4100
rect 16347 4097 16359 4131
rect 16408 4128 16436 4168
rect 17972 4168 18184 4196
rect 21652 4168 21772 4196
rect 17972 4128 18000 4168
rect 16408 4100 18000 4128
rect 16301 4091 16359 4097
rect 18046 4088 18052 4140
rect 18104 4088 18110 4140
rect 18156 4137 18184 4168
rect 18141 4131 18199 4137
rect 18141 4097 18153 4131
rect 18187 4097 18199 4131
rect 18141 4091 18199 4097
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 11296 4032 11652 4060
rect 12069 4063 12127 4069
rect 11296 4020 11302 4032
rect 12069 4029 12081 4063
rect 12115 4060 12127 4063
rect 12802 4060 12808 4072
rect 12115 4032 12808 4060
rect 12115 4029 12127 4032
rect 12069 4023 12127 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 14458 4060 14464 4072
rect 14139 4032 14464 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 14458 4020 14464 4032
rect 14516 4020 14522 4072
rect 15378 4020 15384 4072
rect 15436 4060 15442 4072
rect 15654 4060 15660 4072
rect 15436 4032 15660 4060
rect 15436 4020 15442 4032
rect 15654 4020 15660 4032
rect 15712 4060 15718 4072
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15712 4032 15945 4060
rect 15712 4020 15718 4032
rect 15933 4029 15945 4032
rect 15979 4029 15991 4063
rect 15933 4023 15991 4029
rect 16025 4063 16083 4069
rect 16025 4029 16037 4063
rect 16071 4060 16083 4063
rect 16390 4060 16396 4072
rect 16071 4032 16396 4060
rect 16071 4029 16083 4032
rect 16025 4023 16083 4029
rect 9447 3964 10824 3992
rect 15948 3992 15976 4023
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16482 4020 16488 4072
rect 16540 4060 16546 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16540 4032 16681 4060
rect 16540 4020 16546 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 17405 4063 17463 4069
rect 17405 4060 17417 4063
rect 17184 4032 17417 4060
rect 17184 4020 17190 4032
rect 17405 4029 17417 4032
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 17678 4020 17684 4072
rect 17736 4060 17742 4072
rect 18340 4060 18368 4091
rect 18598 4088 18604 4140
rect 18656 4088 18662 4140
rect 19245 4131 19303 4137
rect 19245 4097 19257 4131
rect 19291 4128 19303 4131
rect 20990 4128 20996 4140
rect 19291 4100 20996 4128
rect 19291 4097 19303 4100
rect 19245 4091 19303 4097
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 21082 4088 21088 4140
rect 21140 4088 21146 4140
rect 21269 4131 21327 4137
rect 21269 4097 21281 4131
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 21284 4060 21312 4091
rect 21358 4088 21364 4140
rect 21416 4088 21422 4140
rect 21450 4088 21456 4140
rect 21508 4088 21514 4140
rect 21744 4128 21772 4168
rect 24302 4156 24308 4208
rect 24360 4156 24366 4208
rect 24394 4156 24400 4208
rect 24452 4156 24458 4208
rect 21744 4100 21864 4128
rect 21542 4060 21548 4072
rect 17736 4032 18368 4060
rect 18524 4032 21220 4060
rect 21284 4032 21548 4060
rect 17736 4020 17742 4032
rect 18524 3992 18552 4032
rect 15948 3964 18552 3992
rect 9447 3961 9459 3964
rect 9401 3955 9459 3961
rect 18598 3952 18604 4004
rect 18656 3992 18662 4004
rect 19061 3995 19119 4001
rect 19061 3992 19073 3995
rect 18656 3964 19073 3992
rect 18656 3952 18662 3964
rect 19061 3961 19073 3964
rect 19107 3961 19119 3995
rect 21192 3992 21220 4032
rect 21542 4020 21548 4032
rect 21600 4020 21606 4072
rect 21836 4060 21864 4100
rect 23566 4088 23572 4140
rect 23624 4088 23630 4140
rect 24118 4088 24124 4140
rect 24176 4088 24182 4140
rect 24489 4131 24547 4137
rect 24489 4097 24501 4131
rect 24535 4097 24547 4131
rect 24489 4091 24547 4097
rect 21836 4032 22140 4060
rect 21450 3992 21456 4004
rect 21192 3964 21456 3992
rect 19061 3955 19119 3961
rect 21450 3952 21456 3964
rect 21508 3992 21514 4004
rect 22112 3992 22140 4032
rect 22186 4020 22192 4072
rect 22244 4020 22250 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 22296 4032 22477 4060
rect 22296 3992 22324 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24504 3992 24532 4091
rect 25314 4088 25320 4140
rect 25372 4088 25378 4140
rect 25685 4131 25743 4137
rect 25685 4097 25697 4131
rect 25731 4128 25743 4131
rect 26050 4128 26056 4140
rect 25731 4100 26056 4128
rect 25731 4097 25743 4100
rect 25685 4091 25743 4097
rect 26050 4088 26056 4100
rect 26108 4088 26114 4140
rect 28626 4088 28632 4140
rect 28684 4088 28690 4140
rect 28997 4131 29055 4137
rect 28997 4097 29009 4131
rect 29043 4128 29055 4131
rect 29086 4128 29092 4140
rect 29043 4100 29092 4128
rect 29043 4097 29055 4100
rect 28997 4091 29055 4097
rect 29086 4088 29092 4100
rect 29144 4088 29150 4140
rect 27430 3992 27436 4004
rect 21508 3964 22048 3992
rect 22112 3964 22324 3992
rect 23492 3964 24532 3992
rect 25700 3964 27436 3992
rect 21508 3952 21514 3964
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8294 3924 8300 3936
rect 8067 3896 8300 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 9493 3927 9551 3933
rect 9493 3893 9505 3927
rect 9539 3924 9551 3927
rect 10134 3924 10140 3936
rect 9539 3896 10140 3924
rect 9539 3893 9551 3896
rect 9493 3887 9551 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10321 3927 10379 3933
rect 10321 3893 10333 3927
rect 10367 3924 10379 3927
rect 10870 3924 10876 3936
rect 10367 3896 10876 3924
rect 10367 3893 10379 3896
rect 10321 3887 10379 3893
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11609 3927 11667 3933
rect 11609 3893 11621 3927
rect 11655 3924 11667 3927
rect 13446 3924 13452 3936
rect 11655 3896 13452 3924
rect 11655 3893 11667 3896
rect 11609 3887 11667 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 13541 3927 13599 3933
rect 13541 3893 13553 3927
rect 13587 3924 13599 3927
rect 14826 3924 14832 3936
rect 13587 3896 14832 3924
rect 13587 3893 13599 3896
rect 13541 3887 13599 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 15746 3884 15752 3936
rect 15804 3924 15810 3936
rect 16206 3924 16212 3936
rect 15804 3896 16212 3924
rect 15804 3884 15810 3896
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 17310 3884 17316 3936
rect 17368 3884 17374 3936
rect 17402 3884 17408 3936
rect 17460 3924 17466 3936
rect 18782 3924 18788 3936
rect 17460 3896 18788 3924
rect 17460 3884 17466 3896
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 21266 3884 21272 3936
rect 21324 3924 21330 3936
rect 21910 3924 21916 3936
rect 21324 3896 21916 3924
rect 21324 3884 21330 3896
rect 21910 3884 21916 3896
rect 21968 3884 21974 3936
rect 22020 3924 22048 3964
rect 22462 3924 22468 3936
rect 22020 3896 22468 3924
rect 22462 3884 22468 3896
rect 22520 3924 22526 3936
rect 23492 3924 23520 3964
rect 22520 3896 23520 3924
rect 22520 3884 22526 3896
rect 23934 3884 23940 3936
rect 23992 3884 23998 3936
rect 24670 3884 24676 3936
rect 24728 3884 24734 3936
rect 25700 3933 25728 3964
rect 27430 3952 27436 3964
rect 27488 3992 27494 4004
rect 27488 3964 28672 3992
rect 27488 3952 27494 3964
rect 25685 3927 25743 3933
rect 25685 3893 25697 3927
rect 25731 3893 25743 3927
rect 25685 3887 25743 3893
rect 25869 3927 25927 3933
rect 25869 3893 25881 3927
rect 25915 3924 25927 3927
rect 26878 3924 26884 3936
rect 25915 3896 26884 3924
rect 25915 3893 25927 3896
rect 25869 3887 25927 3893
rect 26878 3884 26884 3896
rect 26936 3884 26942 3936
rect 27062 3884 27068 3936
rect 27120 3924 27126 3936
rect 28644 3933 28672 3964
rect 28445 3927 28503 3933
rect 28445 3924 28457 3927
rect 27120 3896 28457 3924
rect 27120 3884 27126 3896
rect 28445 3893 28457 3896
rect 28491 3893 28503 3927
rect 28445 3887 28503 3893
rect 28629 3927 28687 3933
rect 28629 3893 28641 3927
rect 28675 3893 28687 3927
rect 28629 3887 28687 3893
rect 1104 3834 36432 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 36432 3834
rect 1104 3760 36432 3782
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9122 3720 9128 3732
rect 8904 3692 9128 3720
rect 8904 3680 8910 3692
rect 9122 3680 9128 3692
rect 9180 3720 9186 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 9180 3692 9413 3720
rect 9180 3680 9186 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 11698 3720 11704 3732
rect 9401 3683 9459 3689
rect 11164 3692 11704 3720
rect 7745 3655 7803 3661
rect 7745 3621 7757 3655
rect 7791 3652 7803 3655
rect 9766 3652 9772 3664
rect 7791 3624 9772 3652
rect 7791 3621 7803 3624
rect 7745 3615 7803 3621
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3553 8263 3587
rect 8205 3547 8263 3553
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8220 3516 8248 3547
rect 8294 3544 8300 3596
rect 8352 3544 8358 3596
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 10778 3584 10784 3596
rect 8536 3556 10784 3584
rect 8536 3544 8542 3556
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 10870 3544 10876 3596
rect 10928 3544 10934 3596
rect 11164 3593 11192 3692
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 11790 3680 11796 3732
rect 11848 3720 11854 3732
rect 12894 3720 12900 3732
rect 11848 3692 12900 3720
rect 11848 3680 11854 3692
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 14458 3720 14464 3732
rect 13955 3692 14464 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 16114 3720 16120 3732
rect 15344 3692 16120 3720
rect 15344 3680 15350 3692
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 19613 3723 19671 3729
rect 19613 3720 19625 3723
rect 19576 3692 19625 3720
rect 19576 3680 19582 3692
rect 19613 3689 19625 3692
rect 19659 3689 19671 3723
rect 19613 3683 19671 3689
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 21545 3723 21603 3729
rect 21545 3720 21557 3723
rect 20680 3692 21557 3720
rect 20680 3680 20686 3692
rect 21545 3689 21557 3692
rect 21591 3689 21603 3723
rect 21545 3683 21603 3689
rect 22066 3692 23612 3720
rect 13173 3655 13231 3661
rect 13173 3621 13185 3655
rect 13219 3652 13231 3655
rect 13998 3652 14004 3664
rect 13219 3624 14004 3652
rect 13219 3621 13231 3624
rect 13173 3615 13231 3621
rect 13998 3612 14004 3624
rect 14056 3612 14062 3664
rect 14093 3655 14151 3661
rect 14093 3621 14105 3655
rect 14139 3652 14151 3655
rect 14182 3652 14188 3664
rect 14139 3624 14188 3652
rect 14139 3621 14151 3624
rect 14093 3615 14151 3621
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 14921 3655 14979 3661
rect 14921 3652 14933 3655
rect 14292 3624 14933 3652
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11238 3584 11244 3596
rect 11195 3556 11244 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11422 3544 11428 3596
rect 11480 3544 11486 3596
rect 13354 3584 13360 3596
rect 12820 3556 13360 3584
rect 7975 3488 8156 3516
rect 8220 3488 8340 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 8128 3460 8156 3488
rect 8110 3408 8116 3460
rect 8168 3408 8174 3460
rect 8312 3448 8340 3488
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 9214 3516 9220 3528
rect 8496 3488 9220 3516
rect 8496 3448 8524 3488
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9306 3476 9312 3528
rect 9364 3476 9370 3528
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 12820 3516 12848 3556
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 14292 3584 14320 3624
rect 14921 3621 14933 3624
rect 14967 3621 14979 3655
rect 14921 3615 14979 3621
rect 17586 3612 17592 3664
rect 17644 3652 17650 3664
rect 20165 3655 20223 3661
rect 20165 3652 20177 3655
rect 17644 3624 20177 3652
rect 17644 3612 17650 3624
rect 20165 3621 20177 3624
rect 20211 3621 20223 3655
rect 20165 3615 20223 3621
rect 21082 3612 21088 3664
rect 21140 3652 21146 3664
rect 22066 3652 22094 3692
rect 21140 3624 22094 3652
rect 21140 3612 21146 3624
rect 22186 3612 22192 3664
rect 22244 3652 22250 3664
rect 23584 3652 23612 3692
rect 24026 3680 24032 3732
rect 24084 3680 24090 3732
rect 26605 3723 26663 3729
rect 26605 3720 26617 3723
rect 24320 3692 26617 3720
rect 24320 3652 24348 3692
rect 26605 3689 26617 3692
rect 26651 3689 26663 3723
rect 26605 3683 26663 3689
rect 27430 3680 27436 3732
rect 27488 3680 27494 3732
rect 35897 3723 35955 3729
rect 35897 3689 35909 3723
rect 35943 3720 35955 3723
rect 35986 3720 35992 3732
rect 35943 3692 35992 3720
rect 35943 3689 35955 3692
rect 35897 3683 35955 3689
rect 35986 3680 35992 3692
rect 36044 3680 36050 3732
rect 22244 3624 22324 3652
rect 23584 3624 24348 3652
rect 22244 3612 22250 3624
rect 13780 3556 14320 3584
rect 13780 3544 13786 3556
rect 14550 3544 14556 3596
rect 14608 3544 14614 3596
rect 14734 3544 14740 3596
rect 14792 3544 14798 3596
rect 15010 3544 15016 3596
rect 15068 3584 15074 3596
rect 15565 3587 15623 3593
rect 15068 3556 15516 3584
rect 15068 3544 15074 3556
rect 12768 3502 12848 3516
rect 12768 3488 12834 3502
rect 12768 3476 12774 3488
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13044 3488 13277 3516
rect 13044 3476 13050 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 13504 3488 14473 3516
rect 13504 3476 13510 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 15197 3519 15255 3525
rect 15197 3485 15209 3519
rect 15243 3516 15255 3519
rect 15378 3516 15384 3528
rect 15243 3488 15384 3516
rect 15243 3485 15255 3488
rect 15197 3479 15255 3485
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15488 3525 15516 3556
rect 15565 3553 15577 3587
rect 15611 3584 15623 3587
rect 15838 3584 15844 3596
rect 15611 3556 15844 3584
rect 15611 3553 15623 3556
rect 15565 3547 15623 3553
rect 15838 3544 15844 3556
rect 15896 3584 15902 3596
rect 16022 3584 16028 3596
rect 15896 3556 16028 3584
rect 15896 3544 15902 3556
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 17310 3544 17316 3596
rect 17368 3544 17374 3596
rect 18230 3544 18236 3596
rect 18288 3544 18294 3596
rect 21174 3584 21180 3596
rect 19812 3556 21180 3584
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 18966 3476 18972 3528
rect 19024 3476 19030 3528
rect 19812 3525 19840 3556
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 21361 3587 21419 3593
rect 21361 3553 21373 3587
rect 21407 3584 21419 3587
rect 21450 3584 21456 3596
rect 21407 3556 21456 3584
rect 21407 3553 21419 3556
rect 21361 3547 21419 3553
rect 21450 3544 21456 3556
rect 21508 3584 21514 3596
rect 22296 3593 22324 3624
rect 26970 3612 26976 3664
rect 27028 3652 27034 3664
rect 27157 3655 27215 3661
rect 27157 3652 27169 3655
rect 27028 3624 27169 3652
rect 27028 3612 27034 3624
rect 27157 3621 27169 3624
rect 27203 3621 27215 3655
rect 27157 3615 27215 3621
rect 22281 3587 22339 3593
rect 21508 3556 22048 3584
rect 21508 3544 21514 3556
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 19889 3519 19947 3525
rect 19889 3485 19901 3519
rect 19935 3485 19947 3519
rect 19889 3479 19947 3485
rect 8312 3420 8524 3448
rect 9140 3420 9628 3448
rect 8754 3340 8760 3392
rect 8812 3340 8818 3392
rect 9140 3389 9168 3420
rect 9125 3383 9183 3389
rect 9125 3349 9137 3383
rect 9171 3349 9183 3383
rect 9600 3380 9628 3420
rect 9858 3408 9864 3460
rect 9916 3408 9922 3460
rect 11701 3451 11759 3457
rect 11701 3417 11713 3451
rect 11747 3417 11759 3451
rect 14182 3448 14188 3460
rect 11701 3411 11759 3417
rect 13188 3420 14188 3448
rect 11606 3380 11612 3392
rect 9600 3352 11612 3380
rect 9125 3343 9183 3349
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 11716 3380 11744 3411
rect 13188 3380 13216 3420
rect 14182 3408 14188 3420
rect 14240 3408 14246 3460
rect 18598 3448 18604 3460
rect 16882 3420 18604 3448
rect 11716 3352 13216 3380
rect 13262 3340 13268 3392
rect 13320 3380 13326 3392
rect 15102 3380 15108 3392
rect 13320 3352 15108 3380
rect 13320 3340 13326 3352
rect 15102 3340 15108 3352
rect 15160 3380 15166 3392
rect 16960 3380 16988 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 19904 3448 19932 3479
rect 20806 3476 20812 3528
rect 20864 3476 20870 3528
rect 21082 3476 21088 3528
rect 21140 3476 21146 3528
rect 21266 3476 21272 3528
rect 21324 3476 21330 3528
rect 21818 3476 21824 3528
rect 21876 3476 21882 3528
rect 22020 3525 22048 3556
rect 22281 3553 22293 3587
rect 22327 3553 22339 3587
rect 22281 3547 22339 3553
rect 22554 3544 22560 3596
rect 22612 3544 22618 3596
rect 23842 3544 23848 3596
rect 23900 3584 23906 3596
rect 24397 3587 24455 3593
rect 24397 3584 24409 3587
rect 23900 3556 24409 3584
rect 23900 3544 23906 3556
rect 24397 3553 24409 3556
rect 24443 3553 24455 3587
rect 24397 3547 24455 3553
rect 24670 3544 24676 3596
rect 24728 3584 24734 3596
rect 25869 3587 25927 3593
rect 25869 3584 25881 3587
rect 24728 3556 25881 3584
rect 24728 3544 24734 3556
rect 25869 3553 25881 3556
rect 25915 3553 25927 3587
rect 28258 3584 28264 3596
rect 25869 3547 25927 3553
rect 26160 3556 28264 3584
rect 26160 3528 26188 3556
rect 28258 3544 28264 3556
rect 28316 3544 28322 3596
rect 21913 3519 21971 3525
rect 21913 3485 21925 3519
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 22005 3519 22063 3525
rect 22005 3485 22017 3519
rect 22051 3485 22063 3519
rect 22005 3479 22063 3485
rect 22189 3519 22247 3525
rect 22189 3485 22201 3519
rect 22235 3516 22247 3519
rect 22235 3488 22324 3516
rect 22235 3485 22247 3488
rect 22189 3479 22247 3485
rect 19576 3420 19932 3448
rect 19576 3408 19582 3420
rect 15160 3352 16988 3380
rect 15160 3340 15166 3352
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 17681 3383 17739 3389
rect 17681 3380 17693 3383
rect 17552 3352 17693 3380
rect 17552 3340 17558 3352
rect 17681 3349 17693 3352
rect 17727 3349 17739 3383
rect 17681 3343 17739 3349
rect 18414 3340 18420 3392
rect 18472 3340 18478 3392
rect 21928 3380 21956 3479
rect 22296 3460 22324 3488
rect 23566 3476 23572 3528
rect 23624 3516 23630 3528
rect 23624 3502 23690 3516
rect 23624 3488 23704 3502
rect 23624 3476 23630 3488
rect 22278 3408 22284 3460
rect 22336 3408 22342 3460
rect 22094 3380 22100 3392
rect 21928 3352 22100 3380
rect 22094 3340 22100 3352
rect 22152 3380 22158 3392
rect 22646 3380 22652 3392
rect 22152 3352 22652 3380
rect 22152 3340 22158 3352
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 23676 3380 23704 3488
rect 26142 3476 26148 3528
rect 26200 3476 26206 3528
rect 26878 3476 26884 3528
rect 26936 3516 26942 3528
rect 26973 3519 27031 3525
rect 26973 3516 26985 3519
rect 26936 3488 26985 3516
rect 26936 3476 26942 3488
rect 26973 3485 26985 3488
rect 27019 3485 27031 3519
rect 26973 3479 27031 3485
rect 27522 3476 27528 3528
rect 27580 3476 27586 3528
rect 27801 3519 27859 3525
rect 27801 3485 27813 3519
rect 27847 3516 27859 3519
rect 28994 3516 29000 3528
rect 27847 3488 29000 3516
rect 27847 3485 27859 3488
rect 27801 3479 27859 3485
rect 28994 3476 29000 3488
rect 29052 3476 29058 3528
rect 36078 3476 36084 3528
rect 36136 3476 36142 3528
rect 25406 3408 25412 3460
rect 25464 3448 25470 3460
rect 26789 3451 26847 3457
rect 25464 3420 25544 3448
rect 25464 3408 25470 3420
rect 25516 3380 25544 3420
rect 26789 3417 26801 3451
rect 26835 3448 26847 3451
rect 26835 3420 27292 3448
rect 26835 3417 26847 3420
rect 26789 3411 26847 3417
rect 23676 3352 25544 3380
rect 26881 3383 26939 3389
rect 26881 3349 26893 3383
rect 26927 3380 26939 3383
rect 27062 3380 27068 3392
rect 26927 3352 27068 3380
rect 26927 3349 26939 3352
rect 26881 3343 26939 3349
rect 27062 3340 27068 3352
rect 27120 3340 27126 3392
rect 27264 3389 27292 3420
rect 27249 3383 27307 3389
rect 27249 3349 27261 3383
rect 27295 3349 27307 3383
rect 27249 3343 27307 3349
rect 1104 3290 36432 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 36432 3290
rect 1104 3216 36432 3238
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 12253 3179 12311 3185
rect 8812 3148 11008 3176
rect 8812 3136 8818 3148
rect 9030 3068 9036 3120
rect 9088 3068 9094 3120
rect 10980 3117 11008 3148
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12986 3176 12992 3188
rect 12299 3148 12992 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 14016 3148 15884 3176
rect 10965 3111 11023 3117
rect 10965 3077 10977 3111
rect 11011 3077 11023 3111
rect 10965 3071 11023 3077
rect 12161 3111 12219 3117
rect 12161 3077 12173 3111
rect 12207 3108 12219 3111
rect 12342 3108 12348 3120
rect 12207 3080 12348 3108
rect 12207 3077 12219 3080
rect 12161 3071 12219 3077
rect 12342 3068 12348 3080
rect 12400 3068 12406 3120
rect 13262 3068 13268 3120
rect 13320 3068 13326 3120
rect 13814 3068 13820 3120
rect 13872 3108 13878 3120
rect 14016 3108 14044 3148
rect 13872 3080 14044 3108
rect 13872 3068 13878 3080
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8294 3040 8300 3052
rect 7883 3012 8300 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8938 3000 8944 3052
rect 8996 3000 9002 3052
rect 9858 3000 9864 3052
rect 9916 3000 9922 3052
rect 11238 3000 11244 3052
rect 11296 3000 11302 3052
rect 12434 3040 12440 3052
rect 12406 3000 12440 3040
rect 12492 3000 12498 3052
rect 14016 3049 14044 3080
rect 15102 3068 15108 3120
rect 15160 3068 15166 3120
rect 15565 3111 15623 3117
rect 15565 3077 15577 3111
rect 15611 3108 15623 3111
rect 15654 3108 15660 3120
rect 15611 3080 15660 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 15654 3068 15660 3080
rect 15712 3068 15718 3120
rect 15856 3108 15884 3148
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 16080 3148 16129 3176
rect 16080 3136 16086 3148
rect 16117 3145 16129 3148
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 16390 3136 16396 3188
rect 16448 3136 16454 3188
rect 16945 3179 17003 3185
rect 16945 3145 16957 3179
rect 16991 3176 17003 3179
rect 18414 3176 18420 3188
rect 16991 3148 18420 3176
rect 16991 3145 17003 3148
rect 16945 3139 17003 3145
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 18782 3136 18788 3188
rect 18840 3176 18846 3188
rect 22094 3176 22100 3188
rect 18840 3148 19932 3176
rect 18840 3136 18846 3148
rect 16666 3108 16672 3120
rect 15856 3080 16672 3108
rect 15856 3049 15884 3080
rect 16666 3068 16672 3080
rect 16724 3108 16730 3120
rect 17586 3108 17592 3120
rect 16724 3080 17592 3108
rect 16724 3068 16730 3080
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 15930 3000 15936 3052
rect 15988 3000 15994 3052
rect 16206 3000 16212 3052
rect 16264 3000 16270 3052
rect 16298 3000 16304 3052
rect 16356 3000 16362 3052
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 17236 3049 17264 3080
rect 17586 3068 17592 3080
rect 17644 3068 17650 3120
rect 19904 3117 19932 3148
rect 20640 3148 22100 3176
rect 19889 3111 19947 3117
rect 19889 3077 19901 3111
rect 19935 3077 19947 3111
rect 19889 3071 19947 3077
rect 20438 3068 20444 3120
rect 20496 3068 20502 3120
rect 20640 3117 20668 3148
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 20625 3111 20683 3117
rect 20625 3077 20637 3111
rect 20671 3077 20683 3111
rect 22186 3108 22192 3120
rect 20625 3071 20683 3077
rect 21836 3080 22192 3108
rect 16485 3043 16543 3049
rect 16485 3040 16497 3043
rect 16448 3012 16497 3040
rect 16448 3000 16454 3012
rect 16485 3009 16497 3012
rect 16531 3040 16543 3043
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16531 3012 16865 3040
rect 16531 3009 16543 3012
rect 16485 3003 16543 3009
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3009 17279 3043
rect 17221 3003 17279 3009
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8478 2972 8484 2984
rect 8067 2944 8484 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2972 8907 2975
rect 9214 2972 9220 2984
rect 8895 2944 9220 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 11517 2975 11575 2981
rect 11517 2972 11529 2975
rect 9364 2944 11529 2972
rect 9364 2932 9370 2944
rect 11517 2941 11529 2944
rect 11563 2972 11575 2975
rect 12406 2972 12434 3000
rect 11563 2944 12434 2972
rect 11563 2941 11575 2944
rect 11517 2935 11575 2941
rect 13722 2932 13728 2984
rect 13780 2932 13786 2984
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14274 2972 14280 2984
rect 14139 2944 14280 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 17144 2972 17172 3003
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 18656 3012 19748 3040
rect 18656 3000 18662 3012
rect 17144 2944 17264 2972
rect 8662 2864 8668 2916
rect 8720 2904 8726 2916
rect 9493 2907 9551 2913
rect 9493 2904 9505 2907
rect 8720 2876 9505 2904
rect 8720 2864 8726 2876
rect 9493 2873 9505 2876
rect 9539 2873 9551 2907
rect 9493 2867 9551 2873
rect 15933 2907 15991 2913
rect 15933 2873 15945 2907
rect 15979 2904 15991 2907
rect 16482 2904 16488 2916
rect 15979 2876 16488 2904
rect 15979 2873 15991 2876
rect 15933 2867 15991 2873
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 17126 2864 17132 2916
rect 17184 2864 17190 2916
rect 7653 2839 7711 2845
rect 7653 2805 7665 2839
rect 7699 2836 7711 2839
rect 8386 2836 8392 2848
rect 7699 2808 8392 2836
rect 7699 2805 7711 2808
rect 7653 2799 7711 2805
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 8938 2836 8944 2848
rect 8619 2808 8944 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 8938 2796 8944 2808
rect 8996 2796 9002 2848
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 9401 2839 9459 2845
rect 9401 2836 9413 2839
rect 9272 2808 9413 2836
rect 9272 2796 9278 2808
rect 9401 2805 9413 2808
rect 9447 2805 9459 2839
rect 9401 2799 9459 2805
rect 12250 2796 12256 2848
rect 12308 2836 12314 2848
rect 14550 2836 14556 2848
rect 12308 2808 14556 2836
rect 12308 2796 12314 2808
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 17236 2836 17264 2944
rect 17494 2932 17500 2984
rect 17552 2932 17558 2984
rect 17862 2932 17868 2984
rect 17920 2972 17926 2984
rect 19613 2975 19671 2981
rect 19613 2972 19625 2975
rect 17920 2944 19625 2972
rect 17920 2932 17926 2944
rect 19613 2941 19625 2944
rect 19659 2941 19671 2975
rect 19720 2972 19748 3012
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 20036 3012 20361 3040
rect 20036 3000 20042 3012
rect 20349 3009 20361 3012
rect 20395 3009 20407 3043
rect 20349 3003 20407 3009
rect 21450 3000 21456 3052
rect 21508 3000 21514 3052
rect 21836 3049 21864 3080
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 23566 3108 23572 3120
rect 23322 3080 23572 3108
rect 23566 3068 23572 3080
rect 23624 3068 23630 3120
rect 34054 3108 34060 3120
rect 24702 3080 34060 3108
rect 34054 3068 34060 3080
rect 34112 3068 34118 3120
rect 21637 3043 21695 3049
rect 21637 3009 21649 3043
rect 21683 3040 21695 3043
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21683 3012 21833 3040
rect 21683 3009 21695 3012
rect 21637 3003 21695 3009
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 25409 3043 25467 3049
rect 25409 3009 25421 3043
rect 25455 3040 25467 3043
rect 26142 3040 26148 3052
rect 25455 3012 26148 3040
rect 25455 3009 25467 3012
rect 25409 3003 25467 3009
rect 26142 3000 26148 3012
rect 26200 3000 26206 3052
rect 20165 2975 20223 2981
rect 20165 2972 20177 2975
rect 19720 2944 20177 2972
rect 19613 2935 19671 2941
rect 20165 2941 20177 2944
rect 20211 2941 20223 2975
rect 21468 2972 21496 3000
rect 22097 2975 22155 2981
rect 22097 2972 22109 2975
rect 21468 2944 22109 2972
rect 20165 2935 20223 2941
rect 22097 2941 22109 2944
rect 22143 2941 22155 2975
rect 22097 2935 22155 2941
rect 25130 2932 25136 2984
rect 25188 2932 25194 2984
rect 21818 2864 21824 2916
rect 21876 2904 21882 2916
rect 21876 2876 21956 2904
rect 21876 2864 21882 2876
rect 17678 2836 17684 2848
rect 17236 2808 17684 2836
rect 17678 2796 17684 2808
rect 17736 2836 17742 2848
rect 18969 2839 19027 2845
rect 18969 2836 18981 2839
rect 17736 2808 18981 2836
rect 17736 2796 17742 2808
rect 18969 2805 18981 2808
rect 19015 2805 19027 2839
rect 18969 2799 19027 2805
rect 19058 2796 19064 2848
rect 19116 2796 19122 2848
rect 20533 2839 20591 2845
rect 20533 2805 20545 2839
rect 20579 2836 20591 2839
rect 20714 2836 20720 2848
rect 20579 2808 20720 2836
rect 20579 2805 20591 2808
rect 20533 2799 20591 2805
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 21266 2796 21272 2848
rect 21324 2796 21330 2848
rect 21928 2836 21956 2876
rect 22554 2836 22560 2848
rect 21928 2808 22560 2836
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 23566 2796 23572 2848
rect 23624 2796 23630 2848
rect 23658 2796 23664 2848
rect 23716 2796 23722 2848
rect 1104 2746 36432 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 36432 2746
rect 1104 2672 36432 2694
rect 7837 2635 7895 2641
rect 7837 2601 7849 2635
rect 7883 2632 7895 2635
rect 10318 2632 10324 2644
rect 7883 2604 10324 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 10778 2632 10784 2644
rect 10735 2604 10784 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 12492 2604 13277 2632
rect 12492 2592 12498 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 13265 2595 13323 2601
rect 13449 2635 13507 2641
rect 13449 2601 13461 2635
rect 13495 2632 13507 2635
rect 13722 2632 13728 2644
rect 13495 2604 13728 2632
rect 13495 2601 13507 2604
rect 13449 2595 13507 2601
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 14826 2592 14832 2644
rect 14884 2632 14890 2644
rect 18417 2635 18475 2641
rect 14884 2604 16528 2632
rect 14884 2592 14890 2604
rect 16209 2567 16267 2573
rect 16209 2533 16221 2567
rect 16255 2564 16267 2567
rect 16298 2564 16304 2576
rect 16255 2536 16304 2564
rect 16255 2533 16267 2536
rect 16209 2527 16267 2533
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8352 2468 8953 2496
rect 8352 2456 8358 2468
rect 8941 2465 8953 2468
rect 8987 2496 8999 2499
rect 11238 2496 11244 2508
rect 8987 2468 11244 2496
rect 8987 2465 8999 2468
rect 8941 2459 8999 2465
rect 11238 2456 11244 2468
rect 11296 2496 11302 2508
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11296 2468 11529 2496
rect 11296 2456 11302 2468
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11517 2459 11575 2465
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 11882 2496 11888 2508
rect 11839 2468 11888 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14461 2499 14519 2505
rect 14461 2496 14473 2499
rect 13872 2468 14473 2496
rect 13872 2456 13878 2468
rect 14461 2465 14473 2468
rect 14507 2465 14519 2499
rect 14461 2459 14519 2465
rect 14737 2499 14795 2505
rect 14737 2465 14749 2499
rect 14783 2496 14795 2499
rect 16393 2499 16451 2505
rect 16393 2496 16405 2499
rect 14783 2468 16405 2496
rect 14783 2465 14795 2468
rect 14737 2459 14795 2465
rect 16393 2465 16405 2468
rect 16439 2465 16451 2499
rect 16393 2459 16451 2465
rect 8018 2388 8024 2440
rect 8076 2388 8082 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8570 2428 8576 2440
rect 8527 2400 8576 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 8404 2360 8432 2391
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10781 2431 10839 2437
rect 10781 2428 10793 2431
rect 10284 2400 10793 2428
rect 10284 2388 10290 2400
rect 10781 2397 10793 2400
rect 10827 2397 10839 2431
rect 10781 2391 10839 2397
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 13538 2388 13544 2440
rect 13596 2388 13602 2440
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 14056 2400 14105 2428
rect 14056 2388 14062 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16500 2428 16528 2604
rect 18417 2601 18429 2635
rect 18463 2632 18475 2635
rect 18966 2632 18972 2644
rect 18463 2604 18972 2632
rect 18463 2601 18475 2604
rect 18417 2595 18475 2601
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 24857 2635 24915 2641
rect 24857 2601 24869 2635
rect 24903 2632 24915 2635
rect 25130 2632 25136 2644
rect 24903 2604 25136 2632
rect 24903 2601 24915 2604
rect 24857 2595 24915 2601
rect 25130 2592 25136 2604
rect 25188 2592 25194 2644
rect 23937 2567 23995 2573
rect 23032 2536 23704 2564
rect 16666 2456 16672 2508
rect 16724 2456 16730 2508
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 19058 2496 19064 2508
rect 16991 2468 19064 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 19058 2456 19064 2468
rect 19116 2456 19122 2508
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 22152 2468 22753 2496
rect 22152 2456 22158 2468
rect 22741 2465 22753 2468
rect 22787 2465 22799 2499
rect 22741 2459 22799 2465
rect 16347 2400 16528 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 20714 2388 20720 2440
rect 20772 2388 20778 2440
rect 21818 2388 21824 2440
rect 21876 2388 21882 2440
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21968 2400 22201 2428
rect 21968 2388 21974 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2428 22615 2431
rect 22646 2428 22652 2440
rect 22603 2400 22652 2428
rect 22603 2397 22615 2400
rect 22557 2391 22615 2397
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 23032 2437 23060 2536
rect 23676 2508 23704 2536
rect 23937 2533 23949 2567
rect 23983 2564 23995 2567
rect 24673 2567 24731 2573
rect 24673 2564 24685 2567
rect 23983 2536 24685 2564
rect 23983 2533 23995 2536
rect 23937 2527 23995 2533
rect 24673 2533 24685 2536
rect 24719 2533 24731 2567
rect 24673 2527 24731 2533
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 23216 2468 23397 2496
rect 23216 2437 23244 2468
rect 23385 2465 23397 2468
rect 23431 2496 23443 2499
rect 23566 2496 23572 2508
rect 23431 2468 23572 2496
rect 23431 2465 23443 2468
rect 23385 2459 23443 2465
rect 23566 2456 23572 2468
rect 23624 2456 23630 2508
rect 23658 2456 23664 2508
rect 23716 2496 23722 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 23716 2468 24409 2496
rect 23716 2456 23722 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 23017 2431 23075 2437
rect 23017 2397 23029 2431
rect 23063 2397 23075 2431
rect 23017 2391 23075 2397
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2397 23259 2431
rect 23201 2391 23259 2397
rect 9122 2360 9128 2372
rect 8404 2332 9128 2360
rect 9122 2320 9128 2332
rect 9180 2320 9186 2372
rect 9214 2320 9220 2372
rect 9272 2320 9278 2372
rect 9858 2320 9864 2372
rect 9916 2320 9922 2372
rect 10612 2332 11100 2360
rect 8202 2252 8208 2304
rect 8260 2252 8266 2304
rect 8665 2295 8723 2301
rect 8665 2261 8677 2295
rect 8711 2292 8723 2295
rect 10612 2292 10640 2332
rect 8711 2264 10640 2292
rect 11072 2292 11100 2332
rect 12526 2320 12532 2372
rect 12584 2320 12590 2372
rect 14366 2320 14372 2372
rect 14424 2360 14430 2372
rect 15194 2360 15200 2372
rect 14424 2332 15200 2360
rect 14424 2320 14430 2332
rect 15194 2320 15200 2332
rect 15252 2320 15258 2372
rect 17402 2360 17408 2372
rect 16040 2332 17408 2360
rect 12158 2292 12164 2304
rect 11072 2264 12164 2292
rect 8711 2261 8723 2264
rect 8665 2255 8723 2261
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 13817 2295 13875 2301
rect 13817 2261 13829 2295
rect 13863 2292 13875 2295
rect 14182 2292 14188 2304
rect 13863 2264 14188 2292
rect 13863 2261 13875 2264
rect 13817 2255 13875 2261
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 14277 2295 14335 2301
rect 14277 2261 14289 2295
rect 14323 2292 14335 2295
rect 15470 2292 15476 2304
rect 14323 2264 15476 2292
rect 14323 2261 14335 2264
rect 14277 2255 14335 2261
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 16040 2292 16068 2332
rect 17402 2320 17408 2332
rect 17460 2320 17466 2372
rect 15620 2264 16068 2292
rect 15620 2252 15626 2264
rect 16482 2252 16488 2304
rect 16540 2292 16546 2304
rect 17862 2292 17868 2304
rect 16540 2264 17868 2292
rect 16540 2252 16546 2264
rect 17862 2252 17868 2264
rect 17920 2252 17926 2304
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 1104 2202 36432 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 36432 2202
rect 1104 2128 36432 2150
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 11606 2088 11612 2100
rect 8260 2060 11612 2088
rect 8260 2048 8266 2060
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16948 37204 17000 37256
rect 17040 37204 17092 37256
rect 21088 37272 21140 37324
rect 25228 37272 25280 37324
rect 22284 37204 22336 37256
rect 22468 37204 22520 37256
rect 23848 37247 23900 37256
rect 23848 37213 23857 37247
rect 23857 37213 23891 37247
rect 23891 37213 23900 37247
rect 23848 37204 23900 37213
rect 29000 37204 29052 37256
rect 29644 37204 29696 37256
rect 16580 37136 16632 37188
rect 17316 37136 17368 37188
rect 18880 37136 18932 37188
rect 22192 37136 22244 37188
rect 17500 37068 17552 37120
rect 18788 37068 18840 37120
rect 20168 37111 20220 37120
rect 20168 37077 20177 37111
rect 20177 37077 20211 37111
rect 20211 37077 20220 37111
rect 20168 37068 20220 37077
rect 21916 37068 21968 37120
rect 23756 37068 23808 37120
rect 29276 37111 29328 37120
rect 29276 37077 29285 37111
rect 29285 37077 29319 37111
rect 29319 37077 29328 37111
rect 29276 37068 29328 37077
rect 29736 37068 29788 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 9680 36796 9732 36848
rect 16120 36864 16172 36916
rect 14832 36728 14884 36780
rect 14924 36771 14976 36780
rect 14924 36737 14933 36771
rect 14933 36737 14967 36771
rect 14967 36737 14976 36771
rect 14924 36728 14976 36737
rect 15292 36728 15344 36780
rect 10692 36660 10744 36712
rect 11060 36703 11112 36712
rect 11060 36669 11069 36703
rect 11069 36669 11103 36703
rect 11103 36669 11112 36703
rect 11060 36660 11112 36669
rect 12624 36703 12676 36712
rect 12624 36669 12633 36703
rect 12633 36669 12667 36703
rect 12667 36669 12676 36703
rect 12624 36660 12676 36669
rect 13268 36660 13320 36712
rect 14096 36660 14148 36712
rect 14740 36703 14792 36712
rect 14740 36669 14749 36703
rect 14749 36669 14783 36703
rect 14783 36669 14792 36703
rect 14740 36660 14792 36669
rect 15844 36771 15896 36780
rect 15844 36737 15853 36771
rect 15853 36737 15887 36771
rect 15887 36737 15896 36771
rect 15844 36728 15896 36737
rect 16580 36796 16632 36848
rect 16488 36771 16540 36780
rect 16488 36737 16497 36771
rect 16497 36737 16531 36771
rect 16531 36737 16540 36771
rect 16488 36728 16540 36737
rect 17776 36796 17828 36848
rect 17500 36771 17552 36780
rect 17500 36737 17509 36771
rect 17509 36737 17543 36771
rect 17543 36737 17552 36771
rect 17500 36728 17552 36737
rect 17592 36771 17644 36780
rect 17592 36737 17627 36771
rect 17627 36737 17644 36771
rect 17592 36728 17644 36737
rect 17224 36660 17276 36712
rect 17868 36660 17920 36712
rect 14280 36592 14332 36644
rect 18236 36771 18288 36780
rect 18236 36737 18245 36771
rect 18245 36737 18279 36771
rect 18279 36737 18288 36771
rect 18236 36728 18288 36737
rect 18144 36660 18196 36712
rect 18328 36703 18380 36712
rect 18328 36669 18337 36703
rect 18337 36669 18371 36703
rect 18371 36669 18380 36703
rect 18328 36660 18380 36669
rect 18420 36703 18472 36712
rect 18420 36669 18429 36703
rect 18429 36669 18463 36703
rect 18463 36669 18472 36703
rect 18420 36660 18472 36669
rect 18788 36728 18840 36780
rect 22560 36864 22612 36916
rect 23296 36796 23348 36848
rect 25780 36796 25832 36848
rect 22100 36728 22152 36780
rect 22468 36728 22520 36780
rect 23848 36771 23900 36780
rect 23848 36737 23857 36771
rect 23857 36737 23891 36771
rect 23891 36737 23900 36771
rect 23848 36728 23900 36737
rect 18696 36660 18748 36712
rect 19616 36703 19668 36712
rect 19616 36669 19625 36703
rect 19625 36669 19659 36703
rect 19659 36669 19668 36703
rect 19616 36660 19668 36669
rect 18604 36592 18656 36644
rect 23480 36660 23532 36712
rect 24400 36660 24452 36712
rect 12716 36524 12768 36576
rect 13636 36524 13688 36576
rect 14188 36524 14240 36576
rect 17132 36567 17184 36576
rect 17132 36533 17141 36567
rect 17141 36533 17175 36567
rect 17175 36533 17184 36567
rect 17132 36524 17184 36533
rect 17960 36524 18012 36576
rect 18144 36524 18196 36576
rect 18328 36524 18380 36576
rect 18788 36567 18840 36576
rect 18788 36533 18797 36567
rect 18797 36533 18831 36567
rect 18831 36533 18840 36567
rect 18788 36524 18840 36533
rect 22192 36524 22244 36576
rect 23204 36524 23256 36576
rect 23388 36524 23440 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 13268 36363 13320 36372
rect 13268 36329 13277 36363
rect 13277 36329 13311 36363
rect 13311 36329 13320 36363
rect 13268 36320 13320 36329
rect 13636 36320 13688 36372
rect 16672 36320 16724 36372
rect 17040 36320 17092 36372
rect 17960 36320 18012 36372
rect 19616 36320 19668 36372
rect 24400 36363 24452 36372
rect 24400 36329 24409 36363
rect 24409 36329 24443 36363
rect 24443 36329 24452 36363
rect 24400 36320 24452 36329
rect 25228 36363 25280 36372
rect 25228 36329 25237 36363
rect 25237 36329 25271 36363
rect 25271 36329 25280 36363
rect 25228 36320 25280 36329
rect 8944 36252 8996 36304
rect 12624 36252 12676 36304
rect 8300 36184 8352 36236
rect 13360 36227 13412 36236
rect 13360 36193 13369 36227
rect 13369 36193 13403 36227
rect 13403 36193 13412 36227
rect 13360 36184 13412 36193
rect 13544 36184 13596 36236
rect 14188 36227 14240 36236
rect 14188 36193 14197 36227
rect 14197 36193 14231 36227
rect 14231 36193 14240 36227
rect 14188 36184 14240 36193
rect 18420 36184 18472 36236
rect 18696 36227 18748 36236
rect 18696 36193 18705 36227
rect 18705 36193 18739 36227
rect 18739 36193 18748 36227
rect 18696 36184 18748 36193
rect 6000 36116 6052 36168
rect 7840 36116 7892 36168
rect 9312 36159 9364 36168
rect 9312 36125 9321 36159
rect 9321 36125 9355 36159
rect 9355 36125 9364 36159
rect 9312 36116 9364 36125
rect 9588 36091 9640 36100
rect 9588 36057 9597 36091
rect 9597 36057 9631 36091
rect 9631 36057 9640 36091
rect 9588 36048 9640 36057
rect 7104 35980 7156 36032
rect 9772 36116 9824 36168
rect 9864 36159 9916 36168
rect 9864 36125 9873 36159
rect 9873 36125 9907 36159
rect 9907 36125 9916 36159
rect 9864 36116 9916 36125
rect 12624 36159 12676 36168
rect 12624 36125 12633 36159
rect 12633 36125 12667 36159
rect 12667 36125 12676 36159
rect 12624 36116 12676 36125
rect 12808 36159 12860 36168
rect 12808 36125 12817 36159
rect 12817 36125 12851 36159
rect 12851 36125 12860 36159
rect 12808 36116 12860 36125
rect 12900 36159 12952 36168
rect 12900 36125 12909 36159
rect 12909 36125 12943 36159
rect 12943 36125 12952 36159
rect 12900 36116 12952 36125
rect 12992 36159 13044 36168
rect 12992 36125 13001 36159
rect 13001 36125 13035 36159
rect 13035 36125 13044 36159
rect 12992 36116 13044 36125
rect 13176 36116 13228 36168
rect 14096 36116 14148 36168
rect 14280 36159 14332 36168
rect 14280 36125 14289 36159
rect 14289 36125 14323 36159
rect 14323 36125 14332 36159
rect 14280 36116 14332 36125
rect 14832 36116 14884 36168
rect 10140 35980 10192 36032
rect 10416 36091 10468 36100
rect 10416 36057 10425 36091
rect 10425 36057 10459 36091
rect 10459 36057 10468 36091
rect 10416 36048 10468 36057
rect 12164 36091 12216 36100
rect 12164 36057 12173 36091
rect 12173 36057 12207 36091
rect 12207 36057 12216 36091
rect 12164 36048 12216 36057
rect 14740 36091 14792 36100
rect 14740 36057 14749 36091
rect 14749 36057 14783 36091
rect 14783 36057 14792 36091
rect 14740 36048 14792 36057
rect 15200 35980 15252 36032
rect 16488 36091 16540 36100
rect 16488 36057 16497 36091
rect 16497 36057 16531 36091
rect 16531 36057 16540 36091
rect 16488 36048 16540 36057
rect 18328 36048 18380 36100
rect 18512 36048 18564 36100
rect 19064 36159 19116 36168
rect 19064 36125 19073 36159
rect 19073 36125 19107 36159
rect 19107 36125 19116 36159
rect 19064 36116 19116 36125
rect 19248 36184 19300 36236
rect 19800 36184 19852 36236
rect 20168 36227 20220 36236
rect 20168 36193 20177 36227
rect 20177 36193 20211 36227
rect 20211 36193 20220 36227
rect 20168 36184 20220 36193
rect 20260 36184 20312 36236
rect 21916 36227 21968 36236
rect 21916 36193 21925 36227
rect 21925 36193 21959 36227
rect 21959 36193 21968 36227
rect 21916 36184 21968 36193
rect 22192 36184 22244 36236
rect 19340 36116 19392 36168
rect 19156 36048 19208 36100
rect 19524 36116 19576 36168
rect 20260 36048 20312 36100
rect 22284 36116 22336 36168
rect 22744 36184 22796 36236
rect 23480 36227 23532 36236
rect 23480 36193 23489 36227
rect 23489 36193 23523 36227
rect 23523 36193 23532 36227
rect 25044 36227 25096 36236
rect 23480 36184 23532 36193
rect 25044 36193 25053 36227
rect 25053 36193 25087 36227
rect 25087 36193 25096 36227
rect 25044 36184 25096 36193
rect 22100 36048 22152 36100
rect 22744 36048 22796 36100
rect 25596 36091 25648 36100
rect 25596 36057 25605 36091
rect 25605 36057 25639 36091
rect 25639 36057 25648 36091
rect 25596 36048 25648 36057
rect 17684 35980 17736 36032
rect 18604 35980 18656 36032
rect 18972 35980 19024 36032
rect 19248 35980 19300 36032
rect 21548 35980 21600 36032
rect 22652 35980 22704 36032
rect 23296 36023 23348 36032
rect 23296 35989 23305 36023
rect 23305 35989 23339 36023
rect 23339 35989 23348 36023
rect 23296 35980 23348 35989
rect 23388 35980 23440 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 8300 35776 8352 35828
rect 7932 35708 7984 35760
rect 6736 35572 6788 35624
rect 8760 35683 8812 35692
rect 8760 35649 8769 35683
rect 8769 35649 8803 35683
rect 8803 35649 8812 35683
rect 8760 35640 8812 35649
rect 8944 35683 8996 35692
rect 8944 35649 8953 35683
rect 8953 35649 8987 35683
rect 8987 35649 8996 35683
rect 8944 35640 8996 35649
rect 9680 35708 9732 35760
rect 10416 35776 10468 35828
rect 11060 35776 11112 35828
rect 12440 35776 12492 35828
rect 12808 35776 12860 35828
rect 12900 35776 12952 35828
rect 15292 35776 15344 35828
rect 15476 35776 15528 35828
rect 7656 35504 7708 35556
rect 6828 35436 6880 35488
rect 8576 35436 8628 35488
rect 8944 35504 8996 35556
rect 9588 35615 9640 35624
rect 9588 35581 9597 35615
rect 9597 35581 9631 35615
rect 9631 35581 9640 35615
rect 9588 35572 9640 35581
rect 9772 35683 9824 35692
rect 9772 35649 9781 35683
rect 9781 35649 9815 35683
rect 9815 35649 9824 35683
rect 9772 35640 9824 35649
rect 10140 35683 10192 35692
rect 10140 35649 10149 35683
rect 10149 35649 10183 35683
rect 10183 35649 10192 35683
rect 10140 35640 10192 35649
rect 10876 35683 10928 35692
rect 10876 35649 10885 35683
rect 10885 35649 10919 35683
rect 10919 35649 10928 35683
rect 10876 35640 10928 35649
rect 10784 35572 10836 35624
rect 10968 35615 11020 35624
rect 10968 35581 10977 35615
rect 10977 35581 11011 35615
rect 11011 35581 11020 35615
rect 10968 35572 11020 35581
rect 11980 35615 12032 35624
rect 11980 35581 11989 35615
rect 11989 35581 12023 35615
rect 12023 35581 12032 35615
rect 11980 35572 12032 35581
rect 11060 35504 11112 35556
rect 11428 35504 11480 35556
rect 13360 35708 13412 35760
rect 16488 35776 16540 35828
rect 18236 35776 18288 35828
rect 22560 35776 22612 35828
rect 12808 35640 12860 35692
rect 12900 35683 12952 35692
rect 12900 35649 12909 35683
rect 12909 35649 12943 35683
rect 12943 35649 12952 35683
rect 12900 35640 12952 35649
rect 12992 35683 13044 35692
rect 12992 35649 13001 35683
rect 13001 35649 13035 35683
rect 13035 35649 13044 35683
rect 12992 35640 13044 35649
rect 13544 35683 13596 35692
rect 13544 35649 13553 35683
rect 13553 35649 13587 35683
rect 13587 35649 13596 35683
rect 13544 35640 13596 35649
rect 13176 35572 13228 35624
rect 13268 35615 13320 35624
rect 13268 35581 13277 35615
rect 13277 35581 13311 35615
rect 13311 35581 13320 35615
rect 13268 35572 13320 35581
rect 14004 35640 14056 35692
rect 14372 35683 14424 35692
rect 14372 35649 14381 35683
rect 14381 35649 14415 35683
rect 14415 35649 14424 35683
rect 14372 35640 14424 35649
rect 13084 35504 13136 35556
rect 10232 35436 10284 35488
rect 11612 35436 11664 35488
rect 13176 35479 13228 35488
rect 13176 35445 13185 35479
rect 13185 35445 13219 35479
rect 13219 35445 13228 35479
rect 13176 35436 13228 35445
rect 13636 35436 13688 35488
rect 14832 35683 14884 35692
rect 14832 35649 14841 35683
rect 14841 35649 14875 35683
rect 14875 35649 14884 35683
rect 14832 35640 14884 35649
rect 14924 35640 14976 35692
rect 15108 35683 15160 35692
rect 15108 35649 15117 35683
rect 15117 35649 15151 35683
rect 15151 35649 15160 35683
rect 15108 35640 15160 35649
rect 15200 35640 15252 35692
rect 16120 35683 16172 35692
rect 16120 35649 16129 35683
rect 16129 35649 16163 35683
rect 16163 35649 16172 35683
rect 16120 35640 16172 35649
rect 16672 35683 16724 35692
rect 16672 35649 16681 35683
rect 16681 35649 16715 35683
rect 16715 35649 16724 35683
rect 16672 35640 16724 35649
rect 17040 35708 17092 35760
rect 18328 35708 18380 35760
rect 18788 35708 18840 35760
rect 15384 35615 15436 35624
rect 15384 35581 15393 35615
rect 15393 35581 15427 35615
rect 15427 35581 15436 35615
rect 15384 35572 15436 35581
rect 14648 35504 14700 35556
rect 16304 35572 16356 35624
rect 16580 35572 16632 35624
rect 17776 35683 17828 35692
rect 17776 35649 17785 35683
rect 17785 35649 17819 35683
rect 17819 35649 17828 35683
rect 17776 35640 17828 35649
rect 18420 35683 18472 35692
rect 18420 35649 18429 35683
rect 18429 35649 18463 35683
rect 18463 35649 18472 35683
rect 18420 35640 18472 35649
rect 20352 35640 20404 35692
rect 17408 35572 17460 35624
rect 17684 35615 17736 35624
rect 17684 35581 17693 35615
rect 17693 35581 17727 35615
rect 17727 35581 17736 35615
rect 17684 35572 17736 35581
rect 17868 35572 17920 35624
rect 21364 35683 21416 35692
rect 21364 35649 21373 35683
rect 21373 35649 21407 35683
rect 21407 35649 21416 35683
rect 21364 35640 21416 35649
rect 23940 35640 23992 35692
rect 24492 35640 24544 35692
rect 24860 35683 24912 35692
rect 24860 35649 24869 35683
rect 24869 35649 24903 35683
rect 24903 35649 24912 35683
rect 24860 35640 24912 35649
rect 21088 35615 21140 35624
rect 21088 35581 21097 35615
rect 21097 35581 21131 35615
rect 21131 35581 21140 35615
rect 21088 35572 21140 35581
rect 22192 35572 22244 35624
rect 22284 35572 22336 35624
rect 22652 35572 22704 35624
rect 23020 35572 23072 35624
rect 26424 35640 26476 35692
rect 25044 35615 25096 35624
rect 25044 35581 25053 35615
rect 25053 35581 25087 35615
rect 25087 35581 25096 35615
rect 25044 35572 25096 35581
rect 13912 35479 13964 35488
rect 13912 35445 13921 35479
rect 13921 35445 13955 35479
rect 13955 35445 13964 35479
rect 13912 35436 13964 35445
rect 14280 35479 14332 35488
rect 14280 35445 14289 35479
rect 14289 35445 14323 35479
rect 14323 35445 14332 35479
rect 14280 35436 14332 35445
rect 16488 35436 16540 35488
rect 16580 35436 16632 35488
rect 21640 35504 21692 35556
rect 19892 35436 19944 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 6000 35275 6052 35284
rect 6000 35241 6009 35275
rect 6009 35241 6043 35275
rect 6043 35241 6052 35275
rect 6000 35232 6052 35241
rect 6736 35275 6788 35284
rect 6736 35241 6745 35275
rect 6745 35241 6779 35275
rect 6779 35241 6788 35275
rect 6736 35232 6788 35241
rect 7840 35275 7892 35284
rect 7840 35241 7849 35275
rect 7849 35241 7883 35275
rect 7883 35241 7892 35275
rect 7840 35232 7892 35241
rect 8208 35232 8260 35284
rect 7380 35164 7432 35216
rect 8760 35232 8812 35284
rect 9312 35275 9364 35284
rect 9312 35241 9321 35275
rect 9321 35241 9355 35275
rect 9355 35241 9364 35275
rect 9312 35232 9364 35241
rect 10876 35232 10928 35284
rect 11980 35275 12032 35284
rect 11980 35241 11989 35275
rect 11989 35241 12023 35275
rect 12023 35241 12032 35275
rect 11980 35232 12032 35241
rect 14372 35232 14424 35284
rect 15108 35232 15160 35284
rect 16304 35232 16356 35284
rect 17408 35232 17460 35284
rect 17776 35232 17828 35284
rect 21640 35232 21692 35284
rect 27068 35232 27120 35284
rect 6828 35096 6880 35148
rect 10968 35164 11020 35216
rect 6092 35071 6144 35080
rect 6092 35037 6101 35071
rect 6101 35037 6135 35071
rect 6135 35037 6144 35071
rect 6092 35028 6144 35037
rect 6276 35071 6328 35080
rect 6276 35037 6285 35071
rect 6285 35037 6319 35071
rect 6319 35037 6328 35071
rect 6276 35028 6328 35037
rect 6368 35071 6420 35080
rect 6368 35037 6377 35071
rect 6377 35037 6411 35071
rect 6411 35037 6420 35071
rect 6368 35028 6420 35037
rect 6460 35071 6512 35080
rect 6460 35037 6469 35071
rect 6469 35037 6503 35071
rect 6503 35037 6512 35071
rect 6460 35028 6512 35037
rect 7104 35071 7156 35080
rect 7104 35037 7113 35071
rect 7113 35037 7147 35071
rect 7147 35037 7156 35071
rect 7104 35028 7156 35037
rect 7288 35028 7340 35080
rect 7656 35071 7708 35080
rect 7656 35037 7665 35071
rect 7665 35037 7699 35071
rect 7699 35037 7708 35071
rect 7656 35028 7708 35037
rect 7932 35071 7984 35080
rect 9036 35096 9088 35148
rect 11336 35139 11388 35148
rect 11336 35105 11345 35139
rect 11345 35105 11379 35139
rect 11379 35105 11388 35139
rect 11336 35096 11388 35105
rect 7932 35037 7947 35071
rect 7947 35037 7981 35071
rect 7981 35037 7984 35071
rect 7932 35028 7984 35037
rect 7012 34892 7064 34944
rect 8576 35071 8628 35080
rect 8576 35037 8585 35071
rect 8585 35037 8619 35071
rect 8619 35037 8628 35071
rect 8576 35028 8628 35037
rect 8944 35071 8996 35080
rect 8944 35037 8953 35071
rect 8953 35037 8987 35071
rect 8987 35037 8996 35071
rect 8944 35028 8996 35037
rect 8852 34960 8904 35012
rect 9588 35028 9640 35080
rect 10232 35071 10284 35080
rect 10232 35037 10241 35071
rect 10241 35037 10275 35071
rect 10275 35037 10284 35071
rect 10232 35028 10284 35037
rect 10692 35028 10744 35080
rect 10968 35028 11020 35080
rect 11428 35028 11480 35080
rect 11520 35071 11572 35080
rect 11520 35037 11529 35071
rect 11529 35037 11563 35071
rect 11563 35037 11572 35071
rect 11520 35028 11572 35037
rect 11612 35071 11664 35080
rect 11612 35037 11621 35071
rect 11621 35037 11655 35071
rect 11655 35037 11664 35071
rect 11612 35028 11664 35037
rect 13636 35164 13688 35216
rect 14188 35164 14240 35216
rect 14924 35164 14976 35216
rect 17592 35164 17644 35216
rect 18696 35164 18748 35216
rect 12900 35096 12952 35148
rect 13176 35096 13228 35148
rect 14004 35096 14056 35148
rect 14556 35096 14608 35148
rect 9864 34960 9916 35012
rect 13912 35028 13964 35080
rect 17316 35096 17368 35148
rect 18420 35096 18472 35148
rect 19616 35096 19668 35148
rect 14096 34960 14148 35012
rect 15016 35028 15068 35080
rect 15384 35071 15436 35080
rect 15384 35037 15393 35071
rect 15393 35037 15427 35071
rect 15427 35037 15436 35071
rect 15384 35028 15436 35037
rect 8760 34935 8812 34944
rect 8760 34901 8769 34935
rect 8769 34901 8803 34935
rect 8803 34901 8812 34935
rect 8760 34892 8812 34901
rect 11060 34892 11112 34944
rect 12164 34892 12216 34944
rect 14004 34892 14056 34944
rect 14188 34892 14240 34944
rect 14648 34892 14700 34944
rect 14740 34935 14792 34944
rect 14740 34901 14749 34935
rect 14749 34901 14783 34935
rect 14783 34901 14792 34935
rect 14740 34892 14792 34901
rect 15292 34935 15344 34944
rect 15292 34901 15301 34935
rect 15301 34901 15335 34935
rect 15335 34901 15344 34935
rect 16304 35028 16356 35080
rect 16488 35071 16540 35080
rect 16488 35037 16497 35071
rect 16497 35037 16531 35071
rect 16531 35037 16540 35071
rect 16488 35028 16540 35037
rect 16856 35028 16908 35080
rect 16764 34960 16816 35012
rect 17868 35028 17920 35080
rect 22284 35096 22336 35148
rect 23848 35096 23900 35148
rect 23020 35071 23072 35080
rect 23020 35037 23029 35071
rect 23029 35037 23063 35071
rect 23063 35037 23072 35071
rect 23020 35028 23072 35037
rect 19616 34960 19668 35012
rect 20168 35003 20220 35012
rect 20168 34969 20177 35003
rect 20177 34969 20211 35003
rect 20211 34969 20220 35003
rect 20168 34960 20220 34969
rect 21548 34960 21600 35012
rect 22560 34960 22612 35012
rect 15292 34892 15344 34901
rect 16396 34935 16448 34944
rect 16396 34901 16405 34935
rect 16405 34901 16439 34935
rect 16439 34901 16448 34935
rect 16396 34892 16448 34901
rect 25320 34960 25372 35012
rect 27528 35071 27580 35080
rect 27528 35037 27537 35071
rect 27537 35037 27571 35071
rect 27571 35037 27580 35071
rect 27528 35028 27580 35037
rect 27804 34960 27856 35012
rect 26608 34892 26660 34944
rect 27344 34892 27396 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 6092 34731 6144 34740
rect 6092 34697 6101 34731
rect 6101 34697 6135 34731
rect 6135 34697 6144 34731
rect 6092 34688 6144 34697
rect 6276 34688 6328 34740
rect 5448 34484 5500 34536
rect 6184 34595 6236 34604
rect 6184 34561 6193 34595
rect 6193 34561 6227 34595
rect 6227 34561 6236 34595
rect 6184 34552 6236 34561
rect 7104 34663 7156 34672
rect 7104 34629 7113 34663
rect 7113 34629 7147 34663
rect 7147 34629 7156 34663
rect 7104 34620 7156 34629
rect 7012 34595 7064 34604
rect 7012 34561 7021 34595
rect 7021 34561 7055 34595
rect 7055 34561 7064 34595
rect 9036 34688 9088 34740
rect 9772 34688 9824 34740
rect 10692 34688 10744 34740
rect 12440 34688 12492 34740
rect 12624 34688 12676 34740
rect 12808 34688 12860 34740
rect 13912 34688 13964 34740
rect 15292 34688 15344 34740
rect 16212 34688 16264 34740
rect 16672 34731 16724 34740
rect 16672 34697 16681 34731
rect 16681 34697 16715 34731
rect 16715 34697 16724 34731
rect 16672 34688 16724 34697
rect 17408 34731 17460 34740
rect 17408 34697 17417 34731
rect 17417 34697 17451 34731
rect 17451 34697 17460 34731
rect 17408 34688 17460 34697
rect 19248 34688 19300 34740
rect 7012 34552 7064 34561
rect 7288 34595 7340 34604
rect 7288 34561 7297 34595
rect 7297 34561 7331 34595
rect 7331 34561 7340 34595
rect 7288 34552 7340 34561
rect 7380 34595 7432 34604
rect 7380 34561 7389 34595
rect 7389 34561 7423 34595
rect 7423 34561 7432 34595
rect 7380 34552 7432 34561
rect 7472 34595 7524 34604
rect 7472 34561 7481 34595
rect 7481 34561 7515 34595
rect 7515 34561 7524 34595
rect 7472 34552 7524 34561
rect 7656 34595 7708 34604
rect 7656 34561 7665 34595
rect 7665 34561 7699 34595
rect 7699 34561 7708 34595
rect 7656 34552 7708 34561
rect 7104 34484 7156 34536
rect 7840 34484 7892 34536
rect 8208 34595 8260 34604
rect 8208 34561 8217 34595
rect 8217 34561 8251 34595
rect 8251 34561 8260 34595
rect 8208 34552 8260 34561
rect 9312 34620 9364 34672
rect 9404 34620 9456 34672
rect 8576 34552 8628 34604
rect 8944 34552 8996 34604
rect 9864 34595 9916 34604
rect 9864 34561 9873 34595
rect 9873 34561 9907 34595
rect 9907 34561 9916 34595
rect 9864 34552 9916 34561
rect 11336 34552 11388 34604
rect 12164 34552 12216 34604
rect 12440 34552 12492 34604
rect 12532 34595 12584 34604
rect 12532 34561 12541 34595
rect 12541 34561 12575 34595
rect 12575 34561 12584 34595
rect 12532 34552 12584 34561
rect 14280 34620 14332 34672
rect 14740 34620 14792 34672
rect 8852 34527 8904 34536
rect 8852 34493 8861 34527
rect 8861 34493 8895 34527
rect 8895 34493 8904 34527
rect 8852 34484 8904 34493
rect 11980 34484 12032 34536
rect 13268 34552 13320 34604
rect 13636 34552 13688 34604
rect 15200 34552 15252 34604
rect 15844 34552 15896 34604
rect 19892 34663 19944 34672
rect 19892 34629 19901 34663
rect 19901 34629 19935 34663
rect 19935 34629 19944 34663
rect 19892 34620 19944 34629
rect 22100 34688 22152 34740
rect 22560 34688 22612 34740
rect 20352 34620 20404 34672
rect 21640 34663 21692 34672
rect 21640 34629 21649 34663
rect 21649 34629 21683 34663
rect 21683 34629 21692 34663
rect 21640 34620 21692 34629
rect 23572 34688 23624 34740
rect 23848 34688 23900 34740
rect 25412 34688 25464 34740
rect 27436 34688 27488 34740
rect 24124 34620 24176 34672
rect 25136 34620 25188 34672
rect 29000 34620 29052 34672
rect 17224 34552 17276 34604
rect 17500 34595 17552 34604
rect 17500 34561 17509 34595
rect 17509 34561 17543 34595
rect 17543 34561 17552 34595
rect 17500 34552 17552 34561
rect 13544 34484 13596 34536
rect 14372 34484 14424 34536
rect 14924 34484 14976 34536
rect 7932 34416 7984 34468
rect 14004 34416 14056 34468
rect 15016 34416 15068 34468
rect 15568 34527 15620 34536
rect 15568 34493 15577 34527
rect 15577 34493 15611 34527
rect 15611 34493 15620 34527
rect 15568 34484 15620 34493
rect 15660 34527 15712 34536
rect 15660 34493 15669 34527
rect 15669 34493 15703 34527
rect 15703 34493 15712 34527
rect 15660 34484 15712 34493
rect 15752 34484 15804 34536
rect 16488 34484 16540 34536
rect 16212 34416 16264 34468
rect 16304 34459 16356 34468
rect 16304 34425 16313 34459
rect 16313 34425 16347 34459
rect 16347 34425 16356 34459
rect 16304 34416 16356 34425
rect 16396 34416 16448 34468
rect 17040 34527 17092 34536
rect 17040 34493 17049 34527
rect 17049 34493 17083 34527
rect 17083 34493 17092 34527
rect 18052 34595 18104 34604
rect 18052 34561 18061 34595
rect 18061 34561 18095 34595
rect 18095 34561 18104 34595
rect 18052 34552 18104 34561
rect 18420 34595 18472 34604
rect 18420 34561 18429 34595
rect 18429 34561 18463 34595
rect 18463 34561 18472 34595
rect 18420 34552 18472 34561
rect 19156 34595 19208 34604
rect 19156 34561 19165 34595
rect 19165 34561 19199 34595
rect 19199 34561 19208 34595
rect 19156 34552 19208 34561
rect 19432 34595 19484 34604
rect 17040 34484 17092 34493
rect 18880 34484 18932 34536
rect 18604 34416 18656 34468
rect 19432 34561 19441 34595
rect 19441 34561 19475 34595
rect 19475 34561 19484 34595
rect 19432 34552 19484 34561
rect 23940 34552 23992 34604
rect 25044 34552 25096 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 22284 34484 22336 34536
rect 22836 34527 22888 34536
rect 22836 34493 22845 34527
rect 22845 34493 22879 34527
rect 22879 34493 22888 34527
rect 22836 34484 22888 34493
rect 24492 34484 24544 34536
rect 26424 34595 26476 34604
rect 26424 34561 26433 34595
rect 26433 34561 26467 34595
rect 26467 34561 26476 34595
rect 26424 34552 26476 34561
rect 27344 34552 27396 34604
rect 26148 34527 26200 34536
rect 26148 34493 26157 34527
rect 26157 34493 26191 34527
rect 26191 34493 26200 34527
rect 26148 34484 26200 34493
rect 27988 34527 28040 34536
rect 27988 34493 27997 34527
rect 27997 34493 28031 34527
rect 28031 34493 28040 34527
rect 27988 34484 28040 34493
rect 31668 34484 31720 34536
rect 19524 34416 19576 34468
rect 7196 34348 7248 34400
rect 13084 34391 13136 34400
rect 13084 34357 13093 34391
rect 13093 34357 13127 34391
rect 13127 34357 13136 34391
rect 13084 34348 13136 34357
rect 13636 34348 13688 34400
rect 14648 34348 14700 34400
rect 16488 34348 16540 34400
rect 18972 34348 19024 34400
rect 19248 34348 19300 34400
rect 23848 34416 23900 34468
rect 27620 34416 27672 34468
rect 24860 34348 24912 34400
rect 28172 34391 28224 34400
rect 28172 34357 28181 34391
rect 28181 34357 28215 34391
rect 28215 34357 28224 34391
rect 28172 34348 28224 34357
rect 28264 34348 28316 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5540 34144 5592 34196
rect 6000 34144 6052 34196
rect 6368 34144 6420 34196
rect 7840 34187 7892 34196
rect 7840 34153 7849 34187
rect 7849 34153 7883 34187
rect 7883 34153 7892 34187
rect 7840 34144 7892 34153
rect 9496 34144 9548 34196
rect 6092 34076 6144 34128
rect 7012 34119 7064 34128
rect 7012 34085 7021 34119
rect 7021 34085 7055 34119
rect 7055 34085 7064 34119
rect 7012 34076 7064 34085
rect 7104 34076 7156 34128
rect 5356 34008 5408 34060
rect 7472 34051 7524 34060
rect 7472 34017 7481 34051
rect 7481 34017 7515 34051
rect 7515 34017 7524 34051
rect 7472 34008 7524 34017
rect 8208 34008 8260 34060
rect 8392 34119 8444 34128
rect 8392 34085 8401 34119
rect 8401 34085 8435 34119
rect 8435 34085 8444 34119
rect 8392 34076 8444 34085
rect 8944 34076 8996 34128
rect 9128 34076 9180 34128
rect 9864 34187 9916 34196
rect 9864 34153 9873 34187
rect 9873 34153 9907 34187
rect 9907 34153 9916 34187
rect 9864 34144 9916 34153
rect 11520 34144 11572 34196
rect 12440 34144 12492 34196
rect 8484 34008 8536 34060
rect 9404 34008 9456 34060
rect 9496 34051 9548 34060
rect 9496 34017 9505 34051
rect 9505 34017 9539 34051
rect 9539 34017 9548 34051
rect 9496 34008 9548 34017
rect 4712 33983 4764 33992
rect 4712 33949 4721 33983
rect 4721 33949 4755 33983
rect 4755 33949 4764 33983
rect 4712 33940 4764 33949
rect 6276 33940 6328 33992
rect 6828 33983 6880 33992
rect 6828 33949 6837 33983
rect 6837 33949 6871 33983
rect 6871 33949 6880 33983
rect 6828 33940 6880 33949
rect 6920 33983 6972 33992
rect 6920 33949 6929 33983
rect 6929 33949 6963 33983
rect 6963 33949 6972 33983
rect 6920 33940 6972 33949
rect 7196 33983 7248 33992
rect 7196 33949 7205 33983
rect 7205 33949 7239 33983
rect 7239 33949 7248 33983
rect 7196 33940 7248 33949
rect 7288 33940 7340 33992
rect 7748 33940 7800 33992
rect 5264 33872 5316 33924
rect 4620 33804 4672 33856
rect 6552 33804 6604 33856
rect 6644 33847 6696 33856
rect 6644 33813 6653 33847
rect 6653 33813 6687 33847
rect 6687 33813 6696 33847
rect 6644 33804 6696 33813
rect 7104 33804 7156 33856
rect 7380 33847 7432 33856
rect 7380 33813 7389 33847
rect 7389 33813 7423 33847
rect 7423 33813 7432 33847
rect 7380 33804 7432 33813
rect 8116 33983 8168 33992
rect 8116 33949 8125 33983
rect 8125 33949 8159 33983
rect 8159 33949 8168 33983
rect 8116 33940 8168 33949
rect 9956 34008 10008 34060
rect 10232 33983 10284 33992
rect 10232 33949 10241 33983
rect 10241 33949 10275 33983
rect 10275 33949 10284 33983
rect 10232 33940 10284 33949
rect 10692 34008 10744 34060
rect 12164 34076 12216 34128
rect 13820 34187 13872 34196
rect 13820 34153 13829 34187
rect 13829 34153 13863 34187
rect 13863 34153 13872 34187
rect 13820 34144 13872 34153
rect 14096 34187 14148 34196
rect 14096 34153 14105 34187
rect 14105 34153 14139 34187
rect 14139 34153 14148 34187
rect 14096 34144 14148 34153
rect 11428 34051 11480 34060
rect 11428 34017 11437 34051
rect 11437 34017 11471 34051
rect 11471 34017 11480 34051
rect 11428 34008 11480 34017
rect 12348 34008 12400 34060
rect 9496 33804 9548 33856
rect 10416 33804 10468 33856
rect 12256 33983 12308 33992
rect 12256 33949 12265 33983
rect 12265 33949 12299 33983
rect 12299 33949 12308 33983
rect 12256 33940 12308 33949
rect 13084 34051 13136 34060
rect 13084 34017 13093 34051
rect 13093 34017 13127 34051
rect 13127 34017 13136 34051
rect 13084 34008 13136 34017
rect 12716 33983 12768 33992
rect 12716 33949 12725 33983
rect 12725 33949 12759 33983
rect 12759 33949 12768 33983
rect 12716 33940 12768 33949
rect 12992 33940 13044 33992
rect 14004 34008 14056 34060
rect 13728 33983 13780 33992
rect 13728 33949 13737 33983
rect 13737 33949 13771 33983
rect 13771 33949 13780 33983
rect 13728 33940 13780 33949
rect 11060 33915 11112 33924
rect 11060 33881 11069 33915
rect 11069 33881 11103 33915
rect 11103 33881 11112 33915
rect 11060 33872 11112 33881
rect 15660 34144 15712 34196
rect 16120 34144 16172 34196
rect 14280 34076 14332 34128
rect 14556 34076 14608 34128
rect 14648 34119 14700 34128
rect 14648 34085 14657 34119
rect 14657 34085 14691 34119
rect 14691 34085 14700 34119
rect 14648 34076 14700 34085
rect 14740 34076 14792 34128
rect 14372 33983 14424 33992
rect 14372 33949 14381 33983
rect 14381 33949 14415 33983
rect 14415 33949 14424 33983
rect 14372 33940 14424 33949
rect 14924 34008 14976 34060
rect 17316 34144 17368 34196
rect 15200 33983 15252 33992
rect 15200 33949 15209 33983
rect 15209 33949 15243 33983
rect 15243 33949 15252 33983
rect 15200 33940 15252 33949
rect 15292 33983 15344 33992
rect 15292 33949 15301 33983
rect 15301 33949 15335 33983
rect 15335 33949 15344 33983
rect 15292 33940 15344 33949
rect 16672 34008 16724 34060
rect 13820 33804 13872 33856
rect 13912 33804 13964 33856
rect 14924 33915 14976 33924
rect 14924 33881 14933 33915
rect 14933 33881 14967 33915
rect 14967 33881 14976 33915
rect 14924 33872 14976 33881
rect 14648 33804 14700 33856
rect 15844 33872 15896 33924
rect 15752 33847 15804 33856
rect 15752 33813 15761 33847
rect 15761 33813 15795 33847
rect 15795 33813 15804 33847
rect 15752 33804 15804 33813
rect 16028 33804 16080 33856
rect 17132 33983 17184 33992
rect 17132 33949 17141 33983
rect 17141 33949 17175 33983
rect 17175 33949 17184 33983
rect 17132 33940 17184 33949
rect 16304 33872 16356 33924
rect 18328 34008 18380 34060
rect 19524 34008 19576 34060
rect 22836 34144 22888 34196
rect 24768 34144 24820 34196
rect 22652 34076 22704 34128
rect 29368 34144 29420 34196
rect 18144 33983 18196 33992
rect 18144 33949 18153 33983
rect 18153 33949 18187 33983
rect 18187 33949 18196 33983
rect 18144 33940 18196 33949
rect 18236 33983 18288 33992
rect 18236 33949 18245 33983
rect 18245 33949 18279 33983
rect 18279 33949 18288 33983
rect 18236 33940 18288 33949
rect 18512 33940 18564 33992
rect 18972 33983 19024 33992
rect 18972 33949 18981 33983
rect 18981 33949 19015 33983
rect 19015 33949 19024 33983
rect 18972 33940 19024 33949
rect 21640 33983 21692 33992
rect 21640 33949 21649 33983
rect 21649 33949 21683 33983
rect 21683 33949 21692 33983
rect 21640 33940 21692 33949
rect 22008 33983 22060 33992
rect 22008 33949 22017 33983
rect 22017 33949 22051 33983
rect 22051 33949 22060 33983
rect 22008 33940 22060 33949
rect 22284 33940 22336 33992
rect 23204 33940 23256 33992
rect 23664 34051 23716 34060
rect 23664 34017 23673 34051
rect 23673 34017 23707 34051
rect 23707 34017 23716 34051
rect 23664 34008 23716 34017
rect 24124 33940 24176 33992
rect 20260 33872 20312 33924
rect 23940 33872 23992 33924
rect 22008 33804 22060 33856
rect 22376 33804 22428 33856
rect 23480 33804 23532 33856
rect 24032 33847 24084 33856
rect 24032 33813 24041 33847
rect 24041 33813 24075 33847
rect 24075 33813 24084 33847
rect 24032 33804 24084 33813
rect 27620 34076 27672 34128
rect 29460 34076 29512 34128
rect 25320 34008 25372 34060
rect 25504 34008 25556 34060
rect 27344 34008 27396 34060
rect 28172 34008 28224 34060
rect 24860 33940 24912 33992
rect 25780 33872 25832 33924
rect 26148 33872 26200 33924
rect 26608 33915 26660 33924
rect 26608 33881 26617 33915
rect 26617 33881 26651 33915
rect 26651 33881 26660 33915
rect 26608 33872 26660 33881
rect 26884 33872 26936 33924
rect 30196 33940 30248 33992
rect 32496 33940 32548 33992
rect 28908 33872 28960 33924
rect 27988 33804 28040 33856
rect 28540 33804 28592 33856
rect 29184 33872 29236 33924
rect 29920 33872 29972 33924
rect 31576 33804 31628 33856
rect 32864 33804 32916 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 5264 33600 5316 33652
rect 6184 33600 6236 33652
rect 5356 33464 5408 33516
rect 5540 33532 5592 33584
rect 7196 33600 7248 33652
rect 8116 33600 8168 33652
rect 8300 33600 8352 33652
rect 9404 33600 9456 33652
rect 10692 33600 10744 33652
rect 11428 33600 11480 33652
rect 12256 33600 12308 33652
rect 14924 33600 14976 33652
rect 15384 33600 15436 33652
rect 6644 33575 6696 33584
rect 6644 33541 6653 33575
rect 6653 33541 6687 33575
rect 6687 33541 6696 33575
rect 6644 33532 6696 33541
rect 5540 33439 5592 33448
rect 5540 33405 5549 33439
rect 5549 33405 5583 33439
rect 5583 33405 5592 33439
rect 5540 33396 5592 33405
rect 5264 33328 5316 33380
rect 6184 33507 6236 33516
rect 6184 33473 6193 33507
rect 6193 33473 6227 33507
rect 6227 33473 6236 33507
rect 6184 33464 6236 33473
rect 6460 33396 6512 33448
rect 6736 33507 6788 33516
rect 6736 33473 6745 33507
rect 6745 33473 6779 33507
rect 6779 33473 6788 33507
rect 6736 33464 6788 33473
rect 7196 33464 7248 33516
rect 7380 33464 7432 33516
rect 6184 33303 6236 33312
rect 6184 33269 6193 33303
rect 6193 33269 6227 33303
rect 6227 33269 6236 33303
rect 6184 33260 6236 33269
rect 7288 33328 7340 33380
rect 6920 33260 6972 33312
rect 7196 33260 7248 33312
rect 9588 33532 9640 33584
rect 9680 33532 9732 33584
rect 12716 33532 12768 33584
rect 8116 33439 8168 33448
rect 8116 33405 8125 33439
rect 8125 33405 8159 33439
rect 8159 33405 8168 33439
rect 8116 33396 8168 33405
rect 8576 33260 8628 33312
rect 10416 33464 10468 33516
rect 9404 33396 9456 33448
rect 11060 33396 11112 33448
rect 11520 33396 11572 33448
rect 9496 33328 9548 33380
rect 10416 33328 10468 33380
rect 12164 33507 12216 33516
rect 12164 33473 12173 33507
rect 12173 33473 12207 33507
rect 12207 33473 12216 33507
rect 12164 33464 12216 33473
rect 12440 33507 12492 33516
rect 12440 33473 12449 33507
rect 12449 33473 12483 33507
rect 12483 33473 12492 33507
rect 12440 33464 12492 33473
rect 12992 33396 13044 33448
rect 13360 33507 13412 33516
rect 13360 33473 13369 33507
rect 13369 33473 13403 33507
rect 13403 33473 13412 33507
rect 13360 33464 13412 33473
rect 13820 33507 13872 33516
rect 13820 33473 13829 33507
rect 13829 33473 13863 33507
rect 13863 33473 13872 33507
rect 13820 33464 13872 33473
rect 14004 33507 14056 33516
rect 14004 33473 14013 33507
rect 14013 33473 14047 33507
rect 14047 33473 14056 33507
rect 14004 33464 14056 33473
rect 14188 33507 14240 33516
rect 14188 33473 14197 33507
rect 14197 33473 14231 33507
rect 14231 33473 14240 33507
rect 14188 33464 14240 33473
rect 14372 33507 14424 33516
rect 14372 33473 14381 33507
rect 14381 33473 14415 33507
rect 14415 33473 14424 33507
rect 14372 33464 14424 33473
rect 14464 33507 14516 33516
rect 14464 33473 14473 33507
rect 14473 33473 14507 33507
rect 14507 33473 14516 33507
rect 14464 33464 14516 33473
rect 11980 33328 12032 33380
rect 13728 33396 13780 33448
rect 13912 33439 13964 33448
rect 13912 33405 13921 33439
rect 13921 33405 13955 33439
rect 13955 33405 13964 33439
rect 13912 33396 13964 33405
rect 14280 33396 14332 33448
rect 14740 33507 14792 33516
rect 14740 33473 14749 33507
rect 14749 33473 14783 33507
rect 14783 33473 14792 33507
rect 14740 33464 14792 33473
rect 15568 33532 15620 33584
rect 15200 33464 15252 33516
rect 16396 33600 16448 33652
rect 18328 33600 18380 33652
rect 18512 33600 18564 33652
rect 19248 33600 19300 33652
rect 20260 33600 20312 33652
rect 15844 33532 15896 33584
rect 16120 33507 16172 33516
rect 16120 33473 16129 33507
rect 16129 33473 16163 33507
rect 16163 33473 16172 33507
rect 16120 33464 16172 33473
rect 16304 33575 16356 33584
rect 16304 33541 16313 33575
rect 16313 33541 16347 33575
rect 16347 33541 16356 33575
rect 16304 33532 16356 33541
rect 16672 33575 16724 33584
rect 16672 33541 16681 33575
rect 16681 33541 16715 33575
rect 16715 33541 16724 33575
rect 16672 33532 16724 33541
rect 18972 33532 19024 33584
rect 19156 33532 19208 33584
rect 21824 33643 21876 33652
rect 21824 33609 21833 33643
rect 21833 33609 21867 33643
rect 21867 33609 21876 33643
rect 21824 33600 21876 33609
rect 23020 33600 23072 33652
rect 22560 33532 22612 33584
rect 24676 33600 24728 33652
rect 25044 33600 25096 33652
rect 25780 33600 25832 33652
rect 16856 33507 16908 33516
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 18052 33464 18104 33516
rect 18512 33464 18564 33516
rect 18604 33507 18656 33516
rect 18604 33473 18613 33507
rect 18613 33473 18647 33507
rect 18647 33473 18656 33507
rect 18604 33464 18656 33473
rect 18696 33507 18748 33516
rect 18696 33473 18705 33507
rect 18705 33473 18739 33507
rect 18739 33473 18748 33507
rect 18696 33464 18748 33473
rect 18880 33507 18932 33516
rect 18880 33473 18889 33507
rect 18889 33473 18923 33507
rect 18923 33473 18932 33507
rect 18880 33464 18932 33473
rect 24400 33532 24452 33584
rect 26700 33600 26752 33652
rect 32312 33600 32364 33652
rect 27988 33532 28040 33584
rect 29920 33532 29972 33584
rect 32864 33532 32916 33584
rect 15292 33439 15344 33448
rect 15292 33405 15301 33439
rect 15301 33405 15335 33439
rect 15335 33405 15344 33439
rect 15292 33396 15344 33405
rect 18420 33396 18472 33448
rect 18788 33396 18840 33448
rect 19156 33396 19208 33448
rect 19432 33396 19484 33448
rect 9404 33260 9456 33312
rect 13268 33328 13320 33380
rect 14096 33328 14148 33380
rect 15568 33371 15620 33380
rect 15568 33337 15577 33371
rect 15577 33337 15611 33371
rect 15611 33337 15620 33371
rect 15568 33328 15620 33337
rect 18696 33328 18748 33380
rect 19524 33328 19576 33380
rect 22744 33396 22796 33448
rect 26056 33464 26108 33516
rect 27436 33507 27488 33516
rect 27436 33473 27445 33507
rect 27445 33473 27479 33507
rect 27479 33473 27488 33507
rect 27436 33464 27488 33473
rect 13912 33260 13964 33312
rect 14648 33260 14700 33312
rect 19432 33260 19484 33312
rect 22284 33260 22336 33312
rect 23204 33260 23256 33312
rect 25504 33396 25556 33448
rect 25964 33396 26016 33448
rect 26424 33396 26476 33448
rect 27160 33396 27212 33448
rect 27712 33439 27764 33448
rect 27712 33405 27721 33439
rect 27721 33405 27755 33439
rect 27755 33405 27764 33439
rect 27712 33396 27764 33405
rect 26884 33328 26936 33380
rect 23664 33303 23716 33312
rect 23664 33269 23673 33303
rect 23673 33269 23707 33303
rect 23707 33269 23716 33303
rect 23664 33260 23716 33269
rect 26240 33303 26292 33312
rect 26240 33269 26249 33303
rect 26249 33269 26283 33303
rect 26283 33269 26292 33303
rect 26240 33260 26292 33269
rect 26608 33260 26660 33312
rect 29000 33464 29052 33516
rect 29460 33507 29512 33516
rect 29460 33473 29469 33507
rect 29469 33473 29503 33507
rect 29503 33473 29512 33507
rect 29460 33464 29512 33473
rect 31668 33507 31720 33516
rect 31668 33473 31677 33507
rect 31677 33473 31711 33507
rect 31711 33473 31720 33507
rect 31668 33464 31720 33473
rect 29184 33439 29236 33448
rect 29184 33405 29193 33439
rect 29193 33405 29227 33439
rect 29227 33405 29236 33439
rect 29184 33396 29236 33405
rect 29644 33439 29696 33448
rect 29644 33405 29653 33439
rect 29653 33405 29687 33439
rect 29687 33405 29696 33439
rect 29644 33396 29696 33405
rect 31392 33439 31444 33448
rect 31392 33405 31401 33439
rect 31401 33405 31435 33439
rect 31435 33405 31444 33439
rect 31392 33396 31444 33405
rect 32404 33439 32456 33448
rect 32404 33405 32413 33439
rect 32413 33405 32447 33439
rect 32447 33405 32456 33439
rect 32404 33396 32456 33405
rect 29368 33260 29420 33312
rect 32220 33260 32272 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4436 32988 4488 33040
rect 5080 33056 5132 33108
rect 5264 33099 5316 33108
rect 5264 33065 5273 33099
rect 5273 33065 5307 33099
rect 5307 33065 5316 33099
rect 5264 33056 5316 33065
rect 5540 33056 5592 33108
rect 6184 33056 6236 33108
rect 5172 32988 5224 33040
rect 6460 33099 6512 33108
rect 6460 33065 6469 33099
rect 6469 33065 6503 33099
rect 6503 33065 6512 33099
rect 6460 33056 6512 33065
rect 6552 33099 6604 33108
rect 6552 33065 6561 33099
rect 6561 33065 6595 33099
rect 6595 33065 6604 33099
rect 6552 33056 6604 33065
rect 6644 33056 6696 33108
rect 7196 33056 7248 33108
rect 7288 33099 7340 33108
rect 7288 33065 7297 33099
rect 7297 33065 7331 33099
rect 7331 33065 7340 33099
rect 7288 33056 7340 33065
rect 8116 33056 8168 33108
rect 10232 33056 10284 33108
rect 10968 33056 11020 33108
rect 3332 32852 3384 32904
rect 4804 32963 4856 32972
rect 4804 32929 4813 32963
rect 4813 32929 4847 32963
rect 4847 32929 4856 32963
rect 4804 32920 4856 32929
rect 2964 32784 3016 32836
rect 4344 32827 4396 32836
rect 4344 32793 4353 32827
rect 4353 32793 4387 32827
rect 4387 32793 4396 32827
rect 4344 32784 4396 32793
rect 5080 32895 5132 32904
rect 5080 32861 5089 32895
rect 5089 32861 5123 32895
rect 5123 32861 5132 32895
rect 5080 32852 5132 32861
rect 5264 32852 5316 32904
rect 5448 32852 5500 32904
rect 5632 32852 5684 32904
rect 5816 32895 5868 32904
rect 5816 32861 5825 32895
rect 5825 32861 5859 32895
rect 5859 32861 5868 32895
rect 5816 32852 5868 32861
rect 5908 32852 5960 32904
rect 6552 32920 6604 32972
rect 6644 32963 6696 32972
rect 6644 32929 6653 32963
rect 6653 32929 6687 32963
rect 6687 32929 6696 32963
rect 6644 32920 6696 32929
rect 6736 32920 6788 32972
rect 6092 32895 6144 32904
rect 6092 32861 6101 32895
rect 6101 32861 6135 32895
rect 6135 32861 6144 32895
rect 6092 32852 6144 32861
rect 6184 32852 6236 32904
rect 4804 32716 4856 32768
rect 5080 32716 5132 32768
rect 5816 32716 5868 32768
rect 6092 32716 6144 32768
rect 6644 32784 6696 32836
rect 7104 32895 7156 32904
rect 7104 32861 7113 32895
rect 7113 32861 7147 32895
rect 7147 32861 7156 32895
rect 7104 32852 7156 32861
rect 7380 32988 7432 33040
rect 7932 32852 7984 32904
rect 8024 32895 8076 32904
rect 8024 32861 8033 32895
rect 8033 32861 8067 32895
rect 8067 32861 8076 32895
rect 8024 32852 8076 32861
rect 8760 32920 8812 32972
rect 10048 32988 10100 33040
rect 10140 32988 10192 33040
rect 12256 33056 12308 33108
rect 18236 33056 18288 33108
rect 18328 33056 18380 33108
rect 22100 33056 22152 33108
rect 7748 32784 7800 32836
rect 8392 32895 8444 32904
rect 8392 32861 8401 32895
rect 8401 32861 8435 32895
rect 8435 32861 8444 32895
rect 8392 32852 8444 32861
rect 9680 32920 9732 32972
rect 9496 32895 9548 32904
rect 9496 32861 9505 32895
rect 9505 32861 9539 32895
rect 9539 32861 9548 32895
rect 9496 32852 9548 32861
rect 10232 32920 10284 32972
rect 11336 32920 11388 32972
rect 8760 32784 8812 32836
rect 9772 32827 9824 32836
rect 9772 32793 9781 32827
rect 9781 32793 9815 32827
rect 9815 32793 9824 32827
rect 9772 32784 9824 32793
rect 10324 32895 10376 32904
rect 10324 32861 10333 32895
rect 10333 32861 10367 32895
rect 10367 32861 10376 32895
rect 10324 32852 10376 32861
rect 10508 32852 10560 32904
rect 10968 32852 11020 32904
rect 15844 32988 15896 33040
rect 12164 32852 12216 32904
rect 6736 32716 6788 32768
rect 6828 32716 6880 32768
rect 9956 32716 10008 32768
rect 10416 32784 10468 32836
rect 10232 32759 10284 32768
rect 10232 32725 10241 32759
rect 10241 32725 10275 32759
rect 10275 32725 10284 32759
rect 10232 32716 10284 32725
rect 10968 32716 11020 32768
rect 14096 32895 14148 32904
rect 14096 32861 14105 32895
rect 14105 32861 14139 32895
rect 14139 32861 14148 32895
rect 14096 32852 14148 32861
rect 16120 32920 16172 32972
rect 19892 32920 19944 32972
rect 22468 33056 22520 33108
rect 24492 33099 24544 33108
rect 24492 33065 24501 33099
rect 24501 33065 24535 33099
rect 24535 33065 24544 33099
rect 24492 33056 24544 33065
rect 24860 33056 24912 33108
rect 24124 32988 24176 33040
rect 24584 32988 24636 33040
rect 29644 33056 29696 33108
rect 22376 32963 22428 32972
rect 22376 32929 22385 32963
rect 22385 32929 22419 32963
rect 22419 32929 22428 32963
rect 22376 32920 22428 32929
rect 23388 32920 23440 32972
rect 23664 32920 23716 32972
rect 16580 32852 16632 32904
rect 20076 32852 20128 32904
rect 20260 32895 20312 32904
rect 20260 32861 20268 32895
rect 20268 32861 20302 32895
rect 20302 32861 20312 32895
rect 20260 32852 20312 32861
rect 14372 32827 14424 32836
rect 14372 32793 14381 32827
rect 14381 32793 14415 32827
rect 14415 32793 14424 32827
rect 14372 32784 14424 32793
rect 14924 32784 14976 32836
rect 14188 32716 14240 32768
rect 19248 32784 19300 32836
rect 21824 32895 21876 32904
rect 21824 32861 21833 32895
rect 21833 32861 21867 32895
rect 21867 32861 21876 32895
rect 21824 32852 21876 32861
rect 24032 32852 24084 32904
rect 24400 32895 24452 32904
rect 24400 32861 24409 32895
rect 24409 32861 24443 32895
rect 24443 32861 24452 32895
rect 24400 32852 24452 32861
rect 24676 32852 24728 32904
rect 24860 32852 24912 32904
rect 25044 32852 25096 32904
rect 19340 32759 19392 32768
rect 19340 32725 19349 32759
rect 19349 32725 19383 32759
rect 19383 32725 19392 32759
rect 19340 32716 19392 32725
rect 20720 32784 20772 32836
rect 21916 32784 21968 32836
rect 25320 32963 25372 32972
rect 25320 32929 25329 32963
rect 25329 32929 25363 32963
rect 25363 32929 25372 32963
rect 28264 33031 28316 33040
rect 28264 32997 28273 33031
rect 28273 32997 28307 33031
rect 28307 32997 28316 33031
rect 28264 32988 28316 32997
rect 28356 32988 28408 33040
rect 30012 32988 30064 33040
rect 31392 33099 31444 33108
rect 31392 33065 31401 33099
rect 31401 33065 31435 33099
rect 31435 33065 31444 33099
rect 31392 33056 31444 33065
rect 32404 33056 32456 33108
rect 25320 32920 25372 32929
rect 27712 32920 27764 32972
rect 25412 32895 25464 32904
rect 25412 32861 25421 32895
rect 25421 32861 25455 32895
rect 25455 32861 25464 32895
rect 25412 32852 25464 32861
rect 25504 32895 25556 32904
rect 25504 32861 25513 32895
rect 25513 32861 25547 32895
rect 25547 32861 25556 32895
rect 25504 32852 25556 32861
rect 25780 32852 25832 32904
rect 27528 32852 27580 32904
rect 19984 32759 20036 32768
rect 19984 32725 19993 32759
rect 19993 32725 20027 32759
rect 20027 32725 20036 32759
rect 19984 32716 20036 32725
rect 21732 32716 21784 32768
rect 23664 32716 23716 32768
rect 24032 32716 24084 32768
rect 24952 32716 25004 32768
rect 26700 32784 26752 32836
rect 27896 32895 27948 32904
rect 27896 32861 27905 32895
rect 27905 32861 27939 32895
rect 27939 32861 27948 32895
rect 27896 32852 27948 32861
rect 29184 32920 29236 32972
rect 29276 32963 29328 32972
rect 29276 32929 29285 32963
rect 29285 32929 29319 32963
rect 29319 32929 29328 32963
rect 29276 32920 29328 32929
rect 31668 32920 31720 32972
rect 28080 32852 28132 32904
rect 28540 32895 28592 32904
rect 28540 32861 28549 32895
rect 28549 32861 28583 32895
rect 28583 32861 28592 32895
rect 28540 32852 28592 32861
rect 28816 32895 28868 32904
rect 28816 32861 28825 32895
rect 28825 32861 28859 32895
rect 28859 32861 28868 32895
rect 28816 32852 28868 32861
rect 29000 32852 29052 32904
rect 29920 32852 29972 32904
rect 31576 32895 31628 32904
rect 31576 32861 31585 32895
rect 31585 32861 31619 32895
rect 31619 32861 31628 32895
rect 31576 32852 31628 32861
rect 32128 32920 32180 32972
rect 28632 32827 28684 32836
rect 28632 32793 28641 32827
rect 28641 32793 28675 32827
rect 28675 32793 28684 32827
rect 28632 32784 28684 32793
rect 31944 32895 31996 32904
rect 31944 32861 31953 32895
rect 31953 32861 31987 32895
rect 31987 32861 31996 32895
rect 31944 32852 31996 32861
rect 32220 32895 32272 32904
rect 32220 32861 32229 32895
rect 32229 32861 32263 32895
rect 32263 32861 32272 32895
rect 32220 32852 32272 32861
rect 32404 32895 32456 32904
rect 32404 32861 32413 32895
rect 32413 32861 32447 32895
rect 32447 32861 32456 32895
rect 32404 32852 32456 32861
rect 33416 32852 33468 32904
rect 25228 32716 25280 32768
rect 26148 32716 26200 32768
rect 27160 32716 27212 32768
rect 30380 32716 30432 32768
rect 31116 32716 31168 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 1308 32444 1360 32496
rect 4620 32512 4672 32564
rect 5264 32512 5316 32564
rect 6092 32512 6144 32564
rect 6736 32555 6788 32564
rect 6736 32521 6745 32555
rect 6745 32521 6779 32555
rect 6779 32521 6788 32555
rect 6736 32512 6788 32521
rect 6920 32512 6972 32564
rect 4436 32444 4488 32496
rect 4712 32376 4764 32428
rect 4804 32419 4856 32428
rect 4804 32385 4813 32419
rect 4813 32385 4847 32419
rect 4847 32385 4856 32419
rect 4804 32376 4856 32385
rect 5264 32419 5316 32428
rect 2504 32308 2556 32360
rect 4620 32308 4672 32360
rect 5264 32385 5273 32419
rect 5273 32385 5307 32419
rect 5307 32385 5316 32419
rect 5264 32376 5316 32385
rect 5448 32376 5500 32428
rect 6460 32444 6512 32496
rect 4528 32240 4580 32292
rect 4896 32240 4948 32292
rect 5724 32351 5776 32360
rect 5724 32317 5733 32351
rect 5733 32317 5767 32351
rect 5767 32317 5776 32351
rect 5724 32308 5776 32317
rect 6184 32308 6236 32360
rect 7104 32376 7156 32428
rect 6552 32308 6604 32360
rect 7472 32419 7524 32428
rect 7472 32385 7481 32419
rect 7481 32385 7515 32419
rect 7515 32385 7524 32419
rect 7472 32376 7524 32385
rect 7564 32419 7616 32428
rect 7564 32385 7573 32419
rect 7573 32385 7607 32419
rect 7607 32385 7616 32419
rect 7564 32376 7616 32385
rect 9864 32512 9916 32564
rect 9036 32487 9088 32496
rect 9036 32453 9045 32487
rect 9045 32453 9079 32487
rect 9079 32453 9088 32487
rect 9036 32444 9088 32453
rect 10600 32487 10652 32496
rect 10600 32453 10609 32487
rect 10609 32453 10643 32487
rect 10643 32453 10652 32487
rect 10600 32444 10652 32453
rect 12900 32512 12952 32564
rect 16764 32512 16816 32564
rect 13912 32444 13964 32496
rect 8300 32376 8352 32428
rect 11796 32419 11848 32428
rect 11796 32385 11805 32419
rect 11805 32385 11839 32419
rect 11839 32385 11848 32419
rect 11796 32376 11848 32385
rect 14648 32376 14700 32428
rect 16580 32444 16632 32496
rect 17500 32444 17552 32496
rect 15844 32419 15896 32428
rect 15844 32385 15853 32419
rect 15853 32385 15887 32419
rect 15887 32385 15896 32419
rect 15844 32376 15896 32385
rect 2596 32172 2648 32224
rect 4988 32172 5040 32224
rect 5080 32215 5132 32224
rect 5080 32181 5089 32215
rect 5089 32181 5123 32215
rect 5123 32181 5132 32215
rect 5080 32172 5132 32181
rect 5448 32215 5500 32224
rect 5448 32181 5457 32215
rect 5457 32181 5491 32215
rect 5491 32181 5500 32215
rect 5448 32172 5500 32181
rect 6092 32240 6144 32292
rect 7472 32240 7524 32292
rect 8484 32308 8536 32360
rect 9496 32308 9548 32360
rect 9588 32308 9640 32360
rect 10324 32308 10376 32360
rect 12348 32308 12400 32360
rect 13912 32308 13964 32360
rect 14924 32308 14976 32360
rect 16212 32419 16264 32428
rect 16212 32385 16221 32419
rect 16221 32385 16255 32419
rect 16255 32385 16264 32419
rect 16212 32376 16264 32385
rect 16396 32376 16448 32428
rect 18880 32512 18932 32564
rect 18328 32444 18380 32496
rect 18052 32376 18104 32428
rect 17684 32351 17736 32360
rect 17684 32317 17693 32351
rect 17693 32317 17727 32351
rect 17727 32317 17736 32351
rect 17684 32308 17736 32317
rect 7932 32240 7984 32292
rect 8392 32240 8444 32292
rect 11244 32240 11296 32292
rect 16120 32240 16172 32292
rect 17960 32351 18012 32360
rect 17960 32317 17969 32351
rect 17969 32317 18003 32351
rect 18003 32317 18012 32351
rect 17960 32308 18012 32317
rect 18420 32419 18472 32428
rect 18420 32385 18429 32419
rect 18429 32385 18463 32419
rect 18463 32385 18472 32419
rect 18420 32376 18472 32385
rect 19800 32512 19852 32564
rect 19892 32555 19944 32564
rect 19892 32521 19901 32555
rect 19901 32521 19935 32555
rect 19935 32521 19944 32555
rect 19892 32512 19944 32521
rect 21640 32512 21692 32564
rect 21732 32512 21784 32564
rect 19248 32419 19300 32428
rect 19248 32385 19257 32419
rect 19257 32385 19291 32419
rect 19291 32385 19300 32419
rect 19248 32376 19300 32385
rect 19340 32419 19392 32428
rect 19340 32385 19349 32419
rect 19349 32385 19383 32419
rect 19383 32385 19392 32419
rect 19340 32376 19392 32385
rect 19432 32419 19484 32428
rect 19432 32385 19441 32419
rect 19441 32385 19475 32419
rect 19475 32385 19484 32419
rect 19432 32376 19484 32385
rect 21272 32444 21324 32496
rect 22008 32512 22060 32564
rect 19984 32376 20036 32428
rect 21640 32419 21692 32428
rect 21640 32385 21649 32419
rect 21649 32385 21683 32419
rect 21683 32385 21692 32419
rect 21640 32376 21692 32385
rect 22560 32444 22612 32496
rect 22744 32555 22796 32564
rect 22744 32521 22753 32555
rect 22753 32521 22787 32555
rect 22787 32521 22796 32555
rect 22744 32512 22796 32521
rect 22928 32512 22980 32564
rect 21824 32419 21876 32428
rect 21824 32385 21833 32419
rect 21833 32385 21867 32419
rect 21867 32385 21876 32419
rect 21824 32376 21876 32385
rect 21916 32419 21968 32428
rect 21916 32385 21926 32419
rect 21926 32385 21960 32419
rect 21960 32385 21968 32419
rect 21916 32376 21968 32385
rect 22836 32376 22888 32428
rect 23480 32555 23532 32564
rect 23480 32521 23489 32555
rect 23489 32521 23523 32555
rect 23523 32521 23532 32555
rect 23480 32512 23532 32521
rect 24124 32512 24176 32564
rect 25320 32512 25372 32564
rect 26056 32512 26108 32564
rect 26240 32512 26292 32564
rect 26516 32512 26568 32564
rect 28080 32512 28132 32564
rect 29184 32512 29236 32564
rect 30288 32512 30340 32564
rect 30380 32555 30432 32564
rect 30380 32521 30389 32555
rect 30389 32521 30423 32555
rect 30423 32521 30432 32555
rect 30380 32512 30432 32521
rect 30748 32555 30800 32564
rect 30748 32521 30757 32555
rect 30757 32521 30791 32555
rect 30791 32521 30800 32555
rect 30748 32512 30800 32521
rect 31300 32512 31352 32564
rect 23204 32444 23256 32496
rect 24860 32444 24912 32496
rect 23388 32419 23440 32428
rect 23388 32385 23397 32419
rect 23397 32385 23431 32419
rect 23431 32385 23440 32419
rect 23388 32376 23440 32385
rect 23756 32376 23808 32428
rect 24308 32376 24360 32428
rect 26424 32444 26476 32496
rect 27528 32444 27580 32496
rect 27712 32444 27764 32496
rect 26608 32419 26660 32428
rect 19340 32240 19392 32292
rect 19892 32240 19944 32292
rect 23480 32308 23532 32360
rect 24032 32351 24084 32360
rect 24032 32317 24041 32351
rect 24041 32317 24075 32351
rect 24075 32317 24084 32351
rect 24032 32308 24084 32317
rect 26608 32385 26617 32419
rect 26617 32385 26651 32419
rect 26651 32385 26660 32419
rect 26608 32376 26660 32385
rect 27988 32376 28040 32428
rect 28172 32487 28224 32496
rect 28172 32453 28181 32487
rect 28181 32453 28215 32487
rect 28215 32453 28224 32487
rect 28172 32444 28224 32453
rect 29920 32487 29972 32496
rect 29920 32453 29929 32487
rect 29929 32453 29963 32487
rect 29963 32453 29972 32487
rect 29920 32444 29972 32453
rect 30012 32487 30064 32496
rect 30012 32453 30021 32487
rect 30021 32453 30055 32487
rect 30055 32453 30064 32487
rect 30012 32444 30064 32453
rect 29092 32376 29144 32428
rect 26240 32308 26292 32360
rect 7380 32172 7432 32224
rect 7656 32172 7708 32224
rect 8852 32172 8904 32224
rect 11428 32172 11480 32224
rect 11888 32172 11940 32224
rect 15476 32172 15528 32224
rect 15936 32215 15988 32224
rect 15936 32181 15945 32215
rect 15945 32181 15979 32215
rect 15979 32181 15988 32215
rect 15936 32172 15988 32181
rect 17500 32215 17552 32224
rect 17500 32181 17509 32215
rect 17509 32181 17543 32215
rect 17543 32181 17552 32215
rect 17500 32172 17552 32181
rect 20444 32172 20496 32224
rect 23112 32172 23164 32224
rect 24308 32172 24360 32224
rect 25136 32172 25188 32224
rect 25688 32172 25740 32224
rect 26148 32172 26200 32224
rect 26424 32351 26476 32360
rect 26424 32317 26433 32351
rect 26433 32317 26467 32351
rect 26467 32317 26476 32351
rect 26424 32308 26476 32317
rect 26516 32351 26568 32360
rect 26516 32317 26525 32351
rect 26525 32317 26559 32351
rect 26559 32317 26568 32351
rect 26516 32308 26568 32317
rect 26976 32351 27028 32360
rect 26976 32317 26985 32351
rect 26985 32317 27019 32351
rect 27019 32317 27028 32351
rect 26976 32308 27028 32317
rect 27712 32308 27764 32360
rect 28356 32308 28408 32360
rect 29276 32419 29328 32428
rect 29276 32385 29285 32419
rect 29285 32385 29319 32419
rect 29319 32385 29328 32419
rect 29276 32376 29328 32385
rect 29644 32419 29696 32428
rect 29644 32385 29653 32419
rect 29653 32385 29687 32419
rect 29687 32385 29696 32419
rect 29644 32376 29696 32385
rect 29828 32419 29880 32428
rect 29828 32385 29835 32419
rect 29835 32385 29880 32419
rect 29828 32376 29880 32385
rect 30196 32376 30248 32428
rect 29460 32308 29512 32360
rect 31024 32444 31076 32496
rect 30472 32376 30524 32428
rect 29736 32240 29788 32292
rect 30656 32351 30708 32360
rect 30656 32317 30665 32351
rect 30665 32317 30699 32351
rect 30699 32317 30708 32351
rect 30656 32308 30708 32317
rect 30932 32351 30984 32360
rect 30932 32317 30941 32351
rect 30941 32317 30975 32351
rect 30975 32317 30984 32351
rect 30932 32308 30984 32317
rect 31300 32419 31352 32428
rect 31300 32385 31309 32419
rect 31309 32385 31343 32419
rect 31343 32385 31352 32419
rect 31300 32376 31352 32385
rect 32220 32512 32272 32564
rect 33416 32555 33468 32564
rect 33416 32521 33425 32555
rect 33425 32521 33459 32555
rect 33459 32521 33468 32555
rect 33416 32512 33468 32521
rect 31852 32444 31904 32496
rect 32680 32487 32732 32496
rect 32680 32453 32689 32487
rect 32689 32453 32723 32487
rect 32723 32453 32732 32487
rect 32680 32444 32732 32453
rect 31576 32376 31628 32428
rect 31484 32308 31536 32360
rect 31576 32240 31628 32292
rect 32588 32419 32640 32428
rect 32588 32385 32597 32419
rect 32597 32385 32631 32419
rect 32631 32385 32640 32419
rect 32588 32376 32640 32385
rect 32772 32419 32824 32428
rect 32772 32385 32781 32419
rect 32781 32385 32815 32419
rect 32815 32385 32824 32419
rect 32772 32376 32824 32385
rect 32312 32351 32364 32360
rect 32312 32317 32321 32351
rect 32321 32317 32355 32351
rect 32355 32317 32364 32351
rect 32312 32308 32364 32317
rect 26424 32172 26476 32224
rect 26792 32215 26844 32224
rect 26792 32181 26801 32215
rect 26801 32181 26835 32215
rect 26835 32181 26844 32215
rect 26792 32172 26844 32181
rect 27804 32215 27856 32224
rect 27804 32181 27813 32215
rect 27813 32181 27847 32215
rect 27847 32181 27856 32215
rect 27804 32172 27856 32181
rect 28172 32172 28224 32224
rect 28632 32215 28684 32224
rect 28632 32181 28641 32215
rect 28641 32181 28675 32215
rect 28675 32181 28684 32215
rect 28632 32172 28684 32181
rect 29460 32172 29512 32224
rect 29644 32172 29696 32224
rect 29920 32172 29972 32224
rect 32128 32240 32180 32292
rect 32864 32172 32916 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2504 31968 2556 32020
rect 4160 31968 4212 32020
rect 4436 31968 4488 32020
rect 7012 31968 7064 32020
rect 7564 31968 7616 32020
rect 8024 32011 8076 32020
rect 8024 31977 8033 32011
rect 8033 31977 8067 32011
rect 8067 31977 8076 32011
rect 8024 31968 8076 31977
rect 10232 31968 10284 32020
rect 10600 31968 10652 32020
rect 2412 31900 2464 31952
rect 1308 31832 1360 31884
rect 2596 31764 2648 31816
rect 2780 31807 2832 31816
rect 2780 31773 2789 31807
rect 2789 31773 2823 31807
rect 2823 31773 2832 31807
rect 2780 31764 2832 31773
rect 3332 31807 3384 31816
rect 3332 31773 3341 31807
rect 3341 31773 3375 31807
rect 3375 31773 3384 31807
rect 3332 31764 3384 31773
rect 6552 31900 6604 31952
rect 6920 31900 6972 31952
rect 3700 31628 3752 31680
rect 4712 31832 4764 31884
rect 5080 31832 5132 31884
rect 5632 31832 5684 31884
rect 5448 31764 5500 31816
rect 5816 31807 5868 31816
rect 5816 31773 5825 31807
rect 5825 31773 5859 31807
rect 5859 31773 5868 31807
rect 5816 31764 5868 31773
rect 6092 31764 6144 31816
rect 7472 31875 7524 31884
rect 7472 31841 7481 31875
rect 7481 31841 7515 31875
rect 7515 31841 7524 31875
rect 7472 31832 7524 31841
rect 8116 31900 8168 31952
rect 8392 31832 8444 31884
rect 4344 31696 4396 31748
rect 5080 31696 5132 31748
rect 6828 31807 6880 31816
rect 6828 31773 6837 31807
rect 6837 31773 6871 31807
rect 6871 31773 6880 31807
rect 6828 31764 6880 31773
rect 7564 31807 7616 31816
rect 7564 31773 7573 31807
rect 7573 31773 7607 31807
rect 7607 31773 7616 31807
rect 7564 31764 7616 31773
rect 7840 31807 7892 31816
rect 7840 31773 7849 31807
rect 7849 31773 7883 31807
rect 7883 31773 7892 31807
rect 7840 31764 7892 31773
rect 4252 31628 4304 31680
rect 4896 31628 4948 31680
rect 5540 31628 5592 31680
rect 5724 31628 5776 31680
rect 7656 31696 7708 31748
rect 6092 31628 6144 31680
rect 6460 31628 6512 31680
rect 8944 31832 8996 31884
rect 9588 31943 9640 31952
rect 9588 31909 9597 31943
rect 9597 31909 9631 31943
rect 9631 31909 9640 31943
rect 9588 31900 9640 31909
rect 10140 31900 10192 31952
rect 13728 32011 13780 32020
rect 13728 31977 13737 32011
rect 13737 31977 13771 32011
rect 13771 31977 13780 32011
rect 13728 31968 13780 31977
rect 9680 31832 9732 31884
rect 10048 31875 10100 31884
rect 10048 31841 10057 31875
rect 10057 31841 10091 31875
rect 10091 31841 10100 31875
rect 10048 31832 10100 31841
rect 14004 31900 14056 31952
rect 15936 31968 15988 32020
rect 17684 31968 17736 32020
rect 15476 31943 15528 31952
rect 15476 31909 15485 31943
rect 15485 31909 15519 31943
rect 15519 31909 15528 31943
rect 15476 31900 15528 31909
rect 17408 31900 17460 31952
rect 19984 31968 20036 32020
rect 20904 31968 20956 32020
rect 21272 31968 21324 32020
rect 22100 31968 22152 32020
rect 23848 31968 23900 32020
rect 17868 31900 17920 31952
rect 19432 31900 19484 31952
rect 8668 31628 8720 31680
rect 9036 31739 9088 31748
rect 9036 31705 9045 31739
rect 9045 31705 9079 31739
rect 9079 31705 9088 31739
rect 9036 31696 9088 31705
rect 9220 31807 9272 31816
rect 9220 31773 9229 31807
rect 9229 31773 9263 31807
rect 9263 31773 9272 31807
rect 9220 31764 9272 31773
rect 9588 31764 9640 31816
rect 9772 31807 9824 31816
rect 9772 31773 9781 31807
rect 9781 31773 9815 31807
rect 9815 31773 9824 31807
rect 9772 31764 9824 31773
rect 10600 31807 10652 31816
rect 10600 31773 10609 31807
rect 10609 31773 10643 31807
rect 10643 31773 10652 31807
rect 10600 31764 10652 31773
rect 10968 31807 11020 31816
rect 10968 31773 10972 31807
rect 10972 31773 11006 31807
rect 11006 31773 11020 31807
rect 10968 31764 11020 31773
rect 11244 31807 11296 31816
rect 11244 31773 11289 31807
rect 11289 31773 11296 31807
rect 11244 31764 11296 31773
rect 11428 31807 11480 31816
rect 11428 31773 11437 31807
rect 11437 31773 11471 31807
rect 11471 31773 11480 31807
rect 11428 31764 11480 31773
rect 9128 31628 9180 31680
rect 9956 31628 10008 31680
rect 10140 31628 10192 31680
rect 11152 31739 11204 31748
rect 11152 31705 11161 31739
rect 11161 31705 11195 31739
rect 11195 31705 11204 31739
rect 11152 31696 11204 31705
rect 14096 31832 14148 31884
rect 14924 31832 14976 31884
rect 18696 31832 18748 31884
rect 19248 31832 19300 31884
rect 12072 31764 12124 31816
rect 13452 31764 13504 31816
rect 15108 31807 15160 31816
rect 15108 31773 15117 31807
rect 15117 31773 15151 31807
rect 15151 31773 15160 31807
rect 15108 31764 15160 31773
rect 12992 31696 13044 31748
rect 14372 31696 14424 31748
rect 11704 31628 11756 31680
rect 15476 31764 15528 31816
rect 17500 31764 17552 31816
rect 17868 31807 17920 31816
rect 17868 31773 17877 31807
rect 17877 31773 17911 31807
rect 17911 31773 17920 31807
rect 17868 31764 17920 31773
rect 21364 31900 21416 31952
rect 22560 31943 22612 31952
rect 22560 31909 22569 31943
rect 22569 31909 22603 31943
rect 22603 31909 22612 31943
rect 22560 31900 22612 31909
rect 17316 31696 17368 31748
rect 15936 31628 15988 31680
rect 18420 31696 18472 31748
rect 19708 31764 19760 31816
rect 19800 31807 19852 31816
rect 19800 31773 19809 31807
rect 19809 31773 19843 31807
rect 19843 31773 19852 31807
rect 19800 31764 19852 31773
rect 20536 31832 20588 31884
rect 21916 31832 21968 31884
rect 24124 31900 24176 31952
rect 25504 31968 25556 32020
rect 25596 31968 25648 32020
rect 27344 31968 27396 32020
rect 28632 31968 28684 32020
rect 29276 31968 29328 32020
rect 24584 31900 24636 31952
rect 25136 31900 25188 31952
rect 19984 31807 20036 31816
rect 19984 31773 19993 31807
rect 19993 31773 20027 31807
rect 20027 31773 20036 31807
rect 19984 31764 20036 31773
rect 21640 31764 21692 31816
rect 22468 31764 22520 31816
rect 24032 31832 24084 31884
rect 24768 31875 24820 31884
rect 21272 31696 21324 31748
rect 22376 31739 22428 31748
rect 22376 31705 22385 31739
rect 22385 31705 22419 31739
rect 22419 31705 22428 31739
rect 22376 31696 22428 31705
rect 23020 31807 23072 31816
rect 23020 31773 23029 31807
rect 23029 31773 23063 31807
rect 23063 31773 23072 31807
rect 23020 31764 23072 31773
rect 17776 31671 17828 31680
rect 17776 31637 17785 31671
rect 17785 31637 17819 31671
rect 17819 31637 17828 31671
rect 17776 31628 17828 31637
rect 20168 31628 20220 31680
rect 23664 31739 23716 31748
rect 23664 31705 23673 31739
rect 23673 31705 23707 31739
rect 23707 31705 23716 31739
rect 23664 31696 23716 31705
rect 24308 31764 24360 31816
rect 24768 31841 24777 31875
rect 24777 31841 24811 31875
rect 24811 31841 24820 31875
rect 24768 31832 24820 31841
rect 26148 31832 26200 31884
rect 27620 31900 27672 31952
rect 27712 31900 27764 31952
rect 27344 31875 27396 31884
rect 27344 31841 27353 31875
rect 27353 31841 27387 31875
rect 27387 31841 27396 31875
rect 27344 31832 27396 31841
rect 28356 31900 28408 31952
rect 29828 31968 29880 32020
rect 30380 32011 30432 32020
rect 30380 31977 30389 32011
rect 30389 31977 30423 32011
rect 30423 31977 30432 32011
rect 30380 31968 30432 31977
rect 31300 31968 31352 32020
rect 32312 31968 32364 32020
rect 32588 32011 32640 32020
rect 32588 31977 32597 32011
rect 32597 31977 32631 32011
rect 32631 31977 32640 32011
rect 32588 31968 32640 31977
rect 30840 31900 30892 31952
rect 32772 31943 32824 31952
rect 32772 31909 32781 31943
rect 32781 31909 32815 31943
rect 32815 31909 32824 31943
rect 32772 31900 32824 31909
rect 24768 31696 24820 31748
rect 24952 31696 25004 31748
rect 25320 31764 25372 31816
rect 25688 31807 25740 31816
rect 25688 31773 25697 31807
rect 25697 31773 25731 31807
rect 25731 31773 25740 31807
rect 25688 31764 25740 31773
rect 25872 31807 25924 31816
rect 25872 31773 25881 31807
rect 25881 31773 25915 31807
rect 25915 31773 25924 31807
rect 25872 31764 25924 31773
rect 26148 31696 26200 31748
rect 26424 31807 26476 31816
rect 26424 31773 26433 31807
rect 26433 31773 26467 31807
rect 26467 31773 26476 31807
rect 26424 31764 26476 31773
rect 27068 31764 27120 31816
rect 27160 31807 27212 31816
rect 27160 31773 27169 31807
rect 27169 31773 27203 31807
rect 27203 31773 27212 31807
rect 27160 31764 27212 31773
rect 27252 31807 27304 31816
rect 27252 31773 27261 31807
rect 27261 31773 27295 31807
rect 27295 31773 27304 31807
rect 27252 31764 27304 31773
rect 27436 31807 27488 31816
rect 27436 31773 27445 31807
rect 27445 31773 27479 31807
rect 27479 31773 27488 31807
rect 27436 31764 27488 31773
rect 27620 31807 27672 31816
rect 27620 31773 27629 31807
rect 27629 31773 27663 31807
rect 27663 31773 27672 31807
rect 27620 31764 27672 31773
rect 28080 31807 28132 31816
rect 28080 31773 28090 31807
rect 28090 31773 28124 31807
rect 28124 31773 28132 31807
rect 28080 31764 28132 31773
rect 28264 31807 28316 31816
rect 28264 31773 28273 31807
rect 28273 31773 28307 31807
rect 28307 31773 28316 31807
rect 28264 31764 28316 31773
rect 28540 31875 28592 31884
rect 28540 31841 28549 31875
rect 28549 31841 28583 31875
rect 28583 31841 28592 31875
rect 28540 31832 28592 31841
rect 28908 31832 28960 31884
rect 31116 31875 31168 31884
rect 31116 31841 31125 31875
rect 31125 31841 31159 31875
rect 31159 31841 31168 31875
rect 31116 31832 31168 31841
rect 31392 31832 31444 31884
rect 31576 31832 31628 31884
rect 28724 31764 28776 31816
rect 28816 31764 28868 31816
rect 28448 31696 28500 31748
rect 23756 31628 23808 31680
rect 24584 31628 24636 31680
rect 25228 31671 25280 31680
rect 25228 31637 25237 31671
rect 25237 31637 25271 31671
rect 25271 31637 25280 31671
rect 25228 31628 25280 31637
rect 25688 31628 25740 31680
rect 25780 31628 25832 31680
rect 26516 31628 26568 31680
rect 27528 31628 27580 31680
rect 28816 31671 28868 31680
rect 28816 31637 28825 31671
rect 28825 31637 28859 31671
rect 28859 31637 28868 31671
rect 28816 31628 28868 31637
rect 29368 31696 29420 31748
rect 30012 31807 30064 31816
rect 30012 31773 30021 31807
rect 30021 31773 30055 31807
rect 30055 31773 30064 31807
rect 30012 31764 30064 31773
rect 30104 31764 30156 31816
rect 30380 31764 30432 31816
rect 30472 31807 30524 31816
rect 30472 31773 30481 31807
rect 30481 31773 30515 31807
rect 30515 31773 30524 31807
rect 30472 31764 30524 31773
rect 30932 31807 30984 31816
rect 30932 31773 30938 31807
rect 30938 31773 30972 31807
rect 30972 31773 30984 31807
rect 30932 31764 30984 31773
rect 31024 31764 31076 31816
rect 31300 31764 31352 31816
rect 29828 31696 29880 31748
rect 31484 31739 31536 31748
rect 31484 31705 31493 31739
rect 31493 31705 31527 31739
rect 31527 31705 31536 31739
rect 31484 31696 31536 31705
rect 31852 31764 31904 31816
rect 30472 31628 30524 31680
rect 31392 31628 31444 31680
rect 32312 31764 32364 31816
rect 32680 31764 32732 31816
rect 32404 31739 32456 31748
rect 32404 31705 32413 31739
rect 32413 31705 32447 31739
rect 32447 31705 32456 31739
rect 32404 31696 32456 31705
rect 32588 31671 32640 31680
rect 32588 31637 32613 31671
rect 32613 31637 32640 31671
rect 32588 31628 32640 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 1308 31356 1360 31408
rect 2412 31399 2464 31408
rect 2412 31365 2421 31399
rect 2421 31365 2455 31399
rect 2455 31365 2464 31399
rect 2412 31356 2464 31365
rect 4252 31424 4304 31476
rect 5724 31424 5776 31476
rect 6828 31424 6880 31476
rect 6920 31467 6972 31476
rect 6920 31433 6929 31467
rect 6929 31433 6963 31467
rect 6963 31433 6972 31467
rect 6920 31424 6972 31433
rect 4160 31399 4212 31408
rect 4160 31365 4169 31399
rect 4169 31365 4203 31399
rect 4203 31365 4212 31399
rect 4160 31356 4212 31365
rect 4620 31356 4672 31408
rect 4712 31288 4764 31340
rect 5540 31356 5592 31408
rect 2780 31220 2832 31272
rect 4068 31220 4120 31272
rect 4620 31220 4672 31272
rect 5172 31331 5224 31340
rect 5172 31297 5181 31331
rect 5181 31297 5215 31331
rect 5215 31297 5224 31331
rect 5172 31288 5224 31297
rect 2964 31152 3016 31204
rect 5540 31263 5592 31272
rect 5540 31229 5549 31263
rect 5549 31229 5583 31263
rect 5583 31229 5592 31263
rect 5540 31220 5592 31229
rect 6276 31288 6328 31340
rect 6552 31331 6604 31340
rect 6552 31297 6561 31331
rect 6561 31297 6595 31331
rect 6595 31297 6604 31331
rect 6552 31288 6604 31297
rect 6828 31288 6880 31340
rect 7656 31424 7708 31476
rect 7932 31424 7984 31476
rect 7472 31356 7524 31408
rect 9220 31424 9272 31476
rect 9680 31424 9732 31476
rect 10048 31424 10100 31476
rect 11796 31424 11848 31476
rect 13912 31424 13964 31476
rect 10876 31356 10928 31408
rect 14372 31424 14424 31476
rect 19340 31424 19392 31476
rect 21088 31424 21140 31476
rect 21180 31424 21232 31476
rect 24308 31424 24360 31476
rect 7380 31331 7432 31340
rect 7380 31297 7389 31331
rect 7389 31297 7423 31331
rect 7423 31297 7432 31331
rect 7380 31288 7432 31297
rect 7840 31288 7892 31340
rect 8484 31331 8536 31340
rect 8484 31297 8493 31331
rect 8493 31297 8527 31331
rect 8527 31297 8536 31331
rect 8484 31288 8536 31297
rect 6920 31220 6972 31272
rect 7564 31220 7616 31272
rect 5724 31152 5776 31204
rect 7472 31152 7524 31204
rect 8576 31152 8628 31204
rect 8944 31331 8996 31340
rect 8944 31297 8953 31331
rect 8953 31297 8987 31331
rect 8987 31297 8996 31331
rect 8944 31288 8996 31297
rect 9128 31331 9180 31340
rect 9128 31297 9137 31331
rect 9137 31297 9171 31331
rect 9171 31297 9180 31331
rect 9128 31288 9180 31297
rect 9220 31331 9272 31340
rect 9220 31297 9229 31331
rect 9229 31297 9263 31331
rect 9263 31297 9272 31331
rect 9220 31288 9272 31297
rect 9496 31288 9548 31340
rect 9956 31288 10008 31340
rect 10692 31288 10744 31340
rect 10140 31220 10192 31272
rect 10508 31220 10560 31272
rect 9128 31152 9180 31204
rect 9772 31152 9824 31204
rect 11336 31331 11388 31340
rect 11336 31297 11345 31331
rect 11345 31297 11379 31331
rect 11379 31297 11388 31331
rect 11336 31288 11388 31297
rect 11704 31331 11756 31340
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 11980 31288 12032 31340
rect 11888 31220 11940 31272
rect 14924 31331 14976 31340
rect 14924 31297 14933 31331
rect 14933 31297 14967 31331
rect 14967 31297 14976 31331
rect 14924 31288 14976 31297
rect 15384 31331 15436 31340
rect 15384 31297 15393 31331
rect 15393 31297 15427 31331
rect 15427 31297 15436 31331
rect 15384 31288 15436 31297
rect 1768 31084 1820 31136
rect 4896 31084 4948 31136
rect 5632 31084 5684 31136
rect 5816 31084 5868 31136
rect 6092 31084 6144 31136
rect 8484 31127 8536 31136
rect 8484 31093 8493 31127
rect 8493 31093 8527 31127
rect 8527 31093 8536 31127
rect 8484 31084 8536 31093
rect 9036 31084 9088 31136
rect 11336 31084 11388 31136
rect 12348 31152 12400 31204
rect 13912 31220 13964 31272
rect 15660 31220 15712 31272
rect 16212 31220 16264 31272
rect 17592 31356 17644 31408
rect 17776 31356 17828 31408
rect 17868 31288 17920 31340
rect 18788 31331 18840 31340
rect 18788 31297 18797 31331
rect 18797 31297 18831 31331
rect 18831 31297 18840 31331
rect 18788 31288 18840 31297
rect 18880 31331 18932 31340
rect 18880 31297 18889 31331
rect 18889 31297 18923 31331
rect 18923 31297 18932 31331
rect 18880 31288 18932 31297
rect 22100 31356 22152 31408
rect 25872 31424 25924 31476
rect 27896 31424 27948 31476
rect 25320 31399 25372 31408
rect 25320 31365 25329 31399
rect 25329 31365 25363 31399
rect 25363 31365 25372 31399
rect 25320 31356 25372 31365
rect 26608 31356 26660 31408
rect 26700 31356 26752 31408
rect 18052 31220 18104 31272
rect 20168 31331 20220 31340
rect 20168 31297 20177 31331
rect 20177 31297 20211 31331
rect 20211 31297 20220 31331
rect 20168 31288 20220 31297
rect 20260 31288 20312 31340
rect 20444 31331 20496 31340
rect 20444 31297 20453 31331
rect 20453 31297 20487 31331
rect 20487 31297 20496 31331
rect 20444 31288 20496 31297
rect 15752 31152 15804 31204
rect 19156 31152 19208 31204
rect 20720 31331 20772 31340
rect 20720 31297 20729 31331
rect 20729 31297 20763 31331
rect 20763 31297 20772 31331
rect 20720 31288 20772 31297
rect 20628 31220 20680 31272
rect 20904 31331 20956 31340
rect 20904 31297 20913 31331
rect 20913 31297 20947 31331
rect 20947 31297 20956 31331
rect 20904 31288 20956 31297
rect 20812 31152 20864 31204
rect 21272 31288 21324 31340
rect 13268 31084 13320 31136
rect 14280 31084 14332 31136
rect 16856 31084 16908 31136
rect 17316 31127 17368 31136
rect 17316 31093 17325 31127
rect 17325 31093 17359 31127
rect 17359 31093 17368 31127
rect 17316 31084 17368 31093
rect 17592 31084 17644 31136
rect 18788 31084 18840 31136
rect 20536 31127 20588 31136
rect 20536 31093 20545 31127
rect 20545 31093 20579 31127
rect 20579 31093 20588 31127
rect 20536 31084 20588 31093
rect 20720 31084 20772 31136
rect 23204 31288 23256 31340
rect 23572 31288 23624 31340
rect 23020 31263 23072 31272
rect 23020 31229 23029 31263
rect 23029 31229 23063 31263
rect 23063 31229 23072 31263
rect 23020 31220 23072 31229
rect 25872 31288 25924 31340
rect 24308 31220 24360 31272
rect 24952 31263 25004 31272
rect 24952 31229 24961 31263
rect 24961 31229 24995 31263
rect 24995 31229 25004 31263
rect 24952 31220 25004 31229
rect 22560 31084 22612 31136
rect 23020 31084 23072 31136
rect 23204 31127 23256 31136
rect 23204 31093 23213 31127
rect 23213 31093 23247 31127
rect 23247 31093 23256 31127
rect 25412 31220 25464 31272
rect 25596 31220 25648 31272
rect 26240 31331 26292 31340
rect 26240 31297 26249 31331
rect 26249 31297 26283 31331
rect 26283 31297 26292 31331
rect 26240 31288 26292 31297
rect 26884 31288 26936 31340
rect 27528 31288 27580 31340
rect 27712 31288 27764 31340
rect 28724 31356 28776 31408
rect 26424 31220 26476 31272
rect 26516 31263 26568 31272
rect 26516 31229 26525 31263
rect 26525 31229 26559 31263
rect 26559 31229 26568 31263
rect 26516 31220 26568 31229
rect 28632 31288 28684 31340
rect 30748 31424 30800 31476
rect 31024 31467 31076 31476
rect 31024 31433 31033 31467
rect 31033 31433 31067 31467
rect 31067 31433 31076 31467
rect 31024 31424 31076 31433
rect 29184 31356 29236 31408
rect 31852 31356 31904 31408
rect 32680 31424 32732 31476
rect 32404 31356 32456 31408
rect 32772 31356 32824 31408
rect 28908 31288 28960 31340
rect 29828 31331 29880 31340
rect 29828 31297 29837 31331
rect 29837 31297 29871 31331
rect 29871 31297 29880 31331
rect 29828 31288 29880 31297
rect 30196 31331 30248 31340
rect 30196 31297 30205 31331
rect 30205 31297 30239 31331
rect 30239 31297 30248 31331
rect 30196 31288 30248 31297
rect 30380 31331 30432 31340
rect 30380 31297 30389 31331
rect 30389 31297 30423 31331
rect 30423 31297 30432 31331
rect 30380 31288 30432 31297
rect 30472 31331 30524 31340
rect 30472 31297 30481 31331
rect 30481 31297 30515 31331
rect 30515 31297 30524 31331
rect 30472 31288 30524 31297
rect 32588 31331 32640 31340
rect 25228 31152 25280 31204
rect 23204 31084 23256 31093
rect 25596 31084 25648 31136
rect 26332 31127 26384 31136
rect 26332 31093 26341 31127
rect 26341 31093 26375 31127
rect 26375 31093 26384 31127
rect 26332 31084 26384 31093
rect 26516 31084 26568 31136
rect 27620 31152 27672 31204
rect 30564 31220 30616 31272
rect 32588 31297 32597 31331
rect 32597 31297 32631 31331
rect 32631 31297 32640 31331
rect 32588 31288 32640 31297
rect 32680 31331 32732 31340
rect 32680 31297 32689 31331
rect 32689 31297 32723 31331
rect 32723 31297 32732 31331
rect 32680 31288 32732 31297
rect 30748 31220 30800 31272
rect 31300 31220 31352 31272
rect 27896 31152 27948 31204
rect 28080 31195 28132 31204
rect 28080 31161 28089 31195
rect 28089 31161 28123 31195
rect 28123 31161 28132 31195
rect 28080 31152 28132 31161
rect 28264 31152 28316 31204
rect 27344 31084 27396 31136
rect 27436 31084 27488 31136
rect 30104 31152 30156 31204
rect 30288 31195 30340 31204
rect 30288 31161 30297 31195
rect 30297 31161 30331 31195
rect 30331 31161 30340 31195
rect 30288 31152 30340 31161
rect 32220 31152 32272 31204
rect 33324 31288 33376 31340
rect 29000 31084 29052 31136
rect 30012 31084 30064 31136
rect 30196 31084 30248 31136
rect 33048 31084 33100 31136
rect 33140 31084 33192 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4068 30880 4120 30932
rect 3148 30812 3200 30864
rect 3700 30744 3752 30796
rect 3240 30676 3292 30728
rect 4620 30880 4672 30932
rect 4896 30880 4948 30932
rect 4988 30880 5040 30932
rect 5724 30880 5776 30932
rect 5908 30880 5960 30932
rect 7564 30880 7616 30932
rect 7840 30880 7892 30932
rect 8484 30880 8536 30932
rect 8668 30880 8720 30932
rect 9220 30880 9272 30932
rect 4436 30744 4488 30796
rect 7288 30812 7340 30864
rect 5172 30744 5224 30796
rect 7748 30812 7800 30864
rect 11244 30880 11296 30932
rect 9680 30812 9732 30864
rect 1768 30651 1820 30660
rect 1768 30617 1777 30651
rect 1777 30617 1811 30651
rect 1811 30617 1820 30651
rect 1768 30608 1820 30617
rect 3056 30608 3108 30660
rect 1308 30540 1360 30592
rect 4804 30676 4856 30728
rect 4528 30540 4580 30592
rect 4988 30651 5040 30660
rect 4988 30617 4997 30651
rect 4997 30617 5031 30651
rect 5031 30617 5040 30651
rect 4988 30608 5040 30617
rect 5540 30676 5592 30728
rect 6736 30719 6788 30728
rect 6736 30685 6745 30719
rect 6745 30685 6779 30719
rect 6779 30685 6788 30719
rect 6736 30676 6788 30685
rect 6920 30719 6972 30728
rect 6920 30685 6929 30719
rect 6929 30685 6963 30719
rect 6963 30685 6972 30719
rect 6920 30676 6972 30685
rect 7104 30719 7156 30728
rect 7104 30685 7113 30719
rect 7113 30685 7147 30719
rect 7147 30685 7156 30719
rect 7104 30676 7156 30685
rect 7196 30676 7248 30728
rect 5724 30608 5776 30660
rect 6092 30608 6144 30660
rect 6460 30608 6512 30660
rect 5356 30540 5408 30592
rect 5540 30583 5592 30592
rect 5540 30549 5549 30583
rect 5549 30549 5583 30583
rect 5583 30549 5592 30583
rect 5540 30540 5592 30549
rect 6000 30583 6052 30592
rect 6000 30549 6009 30583
rect 6009 30549 6043 30583
rect 6043 30549 6052 30583
rect 6000 30540 6052 30549
rect 6552 30583 6604 30592
rect 6552 30549 6561 30583
rect 6561 30549 6595 30583
rect 6595 30549 6604 30583
rect 6552 30540 6604 30549
rect 7564 30719 7616 30728
rect 7564 30685 7573 30719
rect 7573 30685 7607 30719
rect 7607 30685 7616 30719
rect 7564 30676 7616 30685
rect 7932 30719 7984 30728
rect 7932 30685 7941 30719
rect 7941 30685 7975 30719
rect 7975 30685 7984 30719
rect 7932 30676 7984 30685
rect 8116 30719 8168 30728
rect 8116 30685 8125 30719
rect 8125 30685 8159 30719
rect 8159 30685 8168 30719
rect 8116 30676 8168 30685
rect 8668 30744 8720 30796
rect 9312 30744 9364 30796
rect 11152 30812 11204 30864
rect 10232 30744 10284 30796
rect 11428 30787 11480 30796
rect 11428 30753 11437 30787
rect 11437 30753 11471 30787
rect 11471 30753 11480 30787
rect 11428 30744 11480 30753
rect 9588 30676 9640 30728
rect 10416 30676 10468 30728
rect 14280 30880 14332 30932
rect 11980 30676 12032 30728
rect 12348 30676 12400 30728
rect 9496 30608 9548 30660
rect 15016 30812 15068 30864
rect 15292 30812 15344 30864
rect 15936 30812 15988 30864
rect 16212 30744 16264 30796
rect 17868 30880 17920 30932
rect 21364 30923 21416 30932
rect 21364 30889 21373 30923
rect 21373 30889 21407 30923
rect 21407 30889 21416 30923
rect 21364 30880 21416 30889
rect 21732 30880 21784 30932
rect 14832 30676 14884 30728
rect 15752 30676 15804 30728
rect 14096 30651 14148 30660
rect 14096 30617 14105 30651
rect 14105 30617 14139 30651
rect 14139 30617 14148 30651
rect 14096 30608 14148 30617
rect 14648 30651 14700 30660
rect 14648 30617 14657 30651
rect 14657 30617 14691 30651
rect 14691 30617 14700 30651
rect 14648 30608 14700 30617
rect 15660 30608 15712 30660
rect 16120 30719 16172 30728
rect 16120 30685 16129 30719
rect 16129 30685 16163 30719
rect 16163 30685 16172 30719
rect 16120 30676 16172 30685
rect 20996 30812 21048 30864
rect 21916 30812 21968 30864
rect 16212 30651 16264 30660
rect 16212 30617 16221 30651
rect 16221 30617 16255 30651
rect 16255 30617 16264 30651
rect 16212 30608 16264 30617
rect 17960 30676 18012 30728
rect 18880 30676 18932 30728
rect 17684 30651 17736 30660
rect 17684 30617 17693 30651
rect 17693 30617 17727 30651
rect 17727 30617 17736 30651
rect 17684 30608 17736 30617
rect 17868 30651 17920 30660
rect 17868 30617 17877 30651
rect 17877 30617 17911 30651
rect 17911 30617 17920 30651
rect 17868 30608 17920 30617
rect 19340 30676 19392 30728
rect 20168 30744 20220 30796
rect 20904 30744 20956 30796
rect 19800 30719 19852 30728
rect 19800 30685 19809 30719
rect 19809 30685 19843 30719
rect 19843 30685 19852 30719
rect 19800 30676 19852 30685
rect 8116 30540 8168 30592
rect 10508 30583 10560 30592
rect 10508 30549 10517 30583
rect 10517 30549 10551 30583
rect 10551 30549 10560 30583
rect 10508 30540 10560 30549
rect 10876 30540 10928 30592
rect 13176 30583 13228 30592
rect 13176 30549 13185 30583
rect 13185 30549 13219 30583
rect 13219 30549 13228 30583
rect 13176 30540 13228 30549
rect 13268 30540 13320 30592
rect 15200 30540 15252 30592
rect 17132 30583 17184 30592
rect 17132 30549 17141 30583
rect 17141 30549 17175 30583
rect 17175 30549 17184 30583
rect 17132 30540 17184 30549
rect 17224 30540 17276 30592
rect 19248 30608 19300 30660
rect 20260 30676 20312 30728
rect 20720 30676 20772 30728
rect 21732 30719 21784 30728
rect 21732 30685 21741 30719
rect 21741 30685 21775 30719
rect 21775 30685 21784 30719
rect 21732 30676 21784 30685
rect 22008 30719 22060 30728
rect 22008 30685 22017 30719
rect 22017 30685 22051 30719
rect 22051 30685 22060 30719
rect 22008 30676 22060 30685
rect 22836 30880 22888 30932
rect 25872 30880 25924 30932
rect 23020 30812 23072 30864
rect 23388 30812 23440 30864
rect 20628 30608 20680 30660
rect 18880 30583 18932 30592
rect 18880 30549 18889 30583
rect 18889 30549 18923 30583
rect 18923 30549 18932 30583
rect 18880 30540 18932 30549
rect 19156 30540 19208 30592
rect 21364 30583 21416 30592
rect 21364 30549 21373 30583
rect 21373 30549 21407 30583
rect 21407 30549 21416 30583
rect 21364 30540 21416 30549
rect 23204 30676 23256 30728
rect 23480 30676 23532 30728
rect 27620 30880 27672 30932
rect 28080 30880 28132 30932
rect 23940 30676 23992 30728
rect 27528 30744 27580 30796
rect 24860 30676 24912 30728
rect 25044 30676 25096 30728
rect 26608 30719 26660 30728
rect 26608 30685 26617 30719
rect 26617 30685 26651 30719
rect 26651 30685 26660 30719
rect 26608 30676 26660 30685
rect 27068 30719 27120 30728
rect 27068 30685 27077 30719
rect 27077 30685 27111 30719
rect 27111 30685 27120 30719
rect 27068 30676 27120 30685
rect 27436 30676 27488 30728
rect 27620 30719 27672 30728
rect 27620 30685 27629 30719
rect 27629 30685 27663 30719
rect 27663 30685 27672 30719
rect 27620 30676 27672 30685
rect 28540 30744 28592 30796
rect 27896 30719 27948 30728
rect 27896 30685 27905 30719
rect 27905 30685 27939 30719
rect 27939 30685 27948 30719
rect 27896 30676 27948 30685
rect 28080 30719 28132 30728
rect 28080 30685 28089 30719
rect 28089 30685 28123 30719
rect 28123 30685 28132 30719
rect 28080 30676 28132 30685
rect 23204 30540 23256 30592
rect 23572 30540 23624 30592
rect 24216 30651 24268 30660
rect 24216 30617 24225 30651
rect 24225 30617 24259 30651
rect 24259 30617 24268 30651
rect 24216 30608 24268 30617
rect 24308 30608 24360 30660
rect 26332 30651 26384 30660
rect 26332 30617 26341 30651
rect 26341 30617 26375 30651
rect 26375 30617 26384 30651
rect 26332 30608 26384 30617
rect 26424 30608 26476 30660
rect 27712 30608 27764 30660
rect 28724 30676 28776 30728
rect 28632 30651 28684 30660
rect 28632 30617 28641 30651
rect 28641 30617 28675 30651
rect 28675 30617 28684 30651
rect 28632 30608 28684 30617
rect 28908 30812 28960 30864
rect 29000 30744 29052 30796
rect 30472 30812 30524 30864
rect 31484 30880 31536 30932
rect 31668 30812 31720 30864
rect 30288 30744 30340 30796
rect 29368 30676 29420 30728
rect 30012 30676 30064 30728
rect 30196 30676 30248 30728
rect 36268 30676 36320 30728
rect 30748 30651 30800 30660
rect 30748 30617 30757 30651
rect 30757 30617 30791 30651
rect 30791 30617 30800 30651
rect 30748 30608 30800 30617
rect 24768 30540 24820 30592
rect 24860 30583 24912 30592
rect 24860 30549 24869 30583
rect 24869 30549 24903 30583
rect 24903 30549 24912 30583
rect 24860 30540 24912 30549
rect 25412 30540 25464 30592
rect 26148 30540 26200 30592
rect 27620 30540 27672 30592
rect 28172 30540 28224 30592
rect 28816 30540 28868 30592
rect 29552 30583 29604 30592
rect 29552 30549 29561 30583
rect 29561 30549 29595 30583
rect 29595 30549 29604 30583
rect 29552 30540 29604 30549
rect 31300 30540 31352 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 3056 30336 3108 30388
rect 5264 30268 5316 30320
rect 3700 30243 3752 30252
rect 3700 30209 3709 30243
rect 3709 30209 3743 30243
rect 3743 30209 3752 30243
rect 3700 30200 3752 30209
rect 1308 30132 1360 30184
rect 3976 30175 4028 30184
rect 3976 30141 3985 30175
rect 3985 30141 4019 30175
rect 4019 30141 4028 30175
rect 3976 30132 4028 30141
rect 5264 30132 5316 30184
rect 5724 30336 5776 30388
rect 6000 30336 6052 30388
rect 6276 30336 6328 30388
rect 10140 30336 10192 30388
rect 10692 30379 10744 30388
rect 10692 30345 10717 30379
rect 10717 30345 10744 30379
rect 10692 30336 10744 30345
rect 10876 30379 10928 30388
rect 10876 30345 10885 30379
rect 10885 30345 10919 30379
rect 10919 30345 10928 30379
rect 10876 30336 10928 30345
rect 11428 30336 11480 30388
rect 14096 30379 14148 30388
rect 14096 30345 14105 30379
rect 14105 30345 14139 30379
rect 14139 30345 14148 30379
rect 14096 30336 14148 30345
rect 14648 30336 14700 30388
rect 19064 30336 19116 30388
rect 5724 30243 5776 30252
rect 5724 30209 5733 30243
rect 5733 30209 5767 30243
rect 5767 30209 5776 30243
rect 5724 30200 5776 30209
rect 6736 30200 6788 30252
rect 7288 30200 7340 30252
rect 5816 30175 5868 30184
rect 5816 30141 5825 30175
rect 5825 30141 5859 30175
rect 5859 30141 5868 30175
rect 5816 30132 5868 30141
rect 7012 30132 7064 30184
rect 7656 30175 7708 30184
rect 7656 30141 7665 30175
rect 7665 30141 7699 30175
rect 7699 30141 7708 30175
rect 7656 30132 7708 30141
rect 8576 30132 8628 30184
rect 9128 30311 9180 30320
rect 9128 30277 9137 30311
rect 9137 30277 9171 30311
rect 9171 30277 9180 30311
rect 9128 30268 9180 30277
rect 10232 30268 10284 30320
rect 8852 30243 8904 30252
rect 8852 30209 8861 30243
rect 8861 30209 8895 30243
rect 8895 30209 8904 30243
rect 8852 30200 8904 30209
rect 8944 30200 8996 30252
rect 10600 30268 10652 30320
rect 9588 30132 9640 30184
rect 10968 30200 11020 30252
rect 3608 30064 3660 30116
rect 6920 30064 6972 30116
rect 11060 30132 11112 30184
rect 11244 30243 11296 30252
rect 11244 30209 11253 30243
rect 11253 30209 11287 30243
rect 11287 30209 11296 30243
rect 11244 30200 11296 30209
rect 11796 30243 11848 30252
rect 11796 30209 11805 30243
rect 11805 30209 11839 30243
rect 11839 30209 11848 30243
rect 11796 30200 11848 30209
rect 14280 30268 14332 30320
rect 13176 30175 13228 30184
rect 13176 30141 13185 30175
rect 13185 30141 13219 30175
rect 13219 30141 13228 30175
rect 13176 30132 13228 30141
rect 14280 30132 14332 30184
rect 5172 29996 5224 30048
rect 7104 29996 7156 30048
rect 7932 29996 7984 30048
rect 8116 30039 8168 30048
rect 8116 30005 8125 30039
rect 8125 30005 8159 30039
rect 8159 30005 8168 30039
rect 8116 29996 8168 30005
rect 8392 29996 8444 30048
rect 8852 29996 8904 30048
rect 9588 29996 9640 30048
rect 13912 30064 13964 30116
rect 14004 30064 14056 30116
rect 14832 30243 14884 30252
rect 14832 30209 14841 30243
rect 14841 30209 14875 30243
rect 14875 30209 14884 30243
rect 14832 30200 14884 30209
rect 18604 30268 18656 30320
rect 15108 30200 15160 30252
rect 17592 30200 17644 30252
rect 17684 30175 17736 30184
rect 17684 30141 17693 30175
rect 17693 30141 17727 30175
rect 17727 30141 17736 30175
rect 17684 30132 17736 30141
rect 18328 30175 18380 30184
rect 18328 30141 18337 30175
rect 18337 30141 18371 30175
rect 18371 30141 18380 30175
rect 18328 30132 18380 30141
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 18972 30268 19024 30320
rect 18880 30243 18932 30252
rect 18880 30209 18889 30243
rect 18889 30209 18923 30243
rect 18923 30209 18932 30243
rect 18880 30200 18932 30209
rect 19616 30336 19668 30388
rect 20720 30336 20772 30388
rect 21824 30336 21876 30388
rect 24860 30336 24912 30388
rect 10784 29996 10836 30048
rect 11612 29996 11664 30048
rect 13268 29996 13320 30048
rect 16856 30064 16908 30116
rect 18972 30132 19024 30184
rect 19248 30243 19300 30252
rect 19248 30209 19257 30243
rect 19257 30209 19291 30243
rect 19291 30209 19300 30243
rect 19248 30200 19300 30209
rect 19340 30175 19392 30184
rect 19340 30141 19349 30175
rect 19349 30141 19383 30175
rect 19383 30141 19392 30175
rect 19340 30132 19392 30141
rect 21640 30268 21692 30320
rect 20628 30200 20680 30252
rect 20720 30200 20772 30252
rect 22008 30243 22060 30252
rect 22008 30209 22017 30243
rect 22017 30209 22051 30243
rect 22051 30209 22060 30243
rect 22008 30200 22060 30209
rect 22468 30200 22520 30252
rect 23204 30268 23256 30320
rect 22744 30243 22796 30252
rect 22744 30209 22753 30243
rect 22753 30209 22787 30243
rect 22787 30209 22796 30243
rect 22744 30200 22796 30209
rect 22836 30243 22888 30252
rect 23848 30268 23900 30320
rect 24308 30268 24360 30320
rect 24492 30268 24544 30320
rect 26884 30336 26936 30388
rect 27068 30336 27120 30388
rect 27436 30336 27488 30388
rect 27712 30336 27764 30388
rect 27988 30336 28040 30388
rect 22836 30209 22871 30243
rect 22871 30209 22888 30243
rect 22836 30200 22888 30209
rect 22376 30132 22428 30184
rect 22284 30064 22336 30116
rect 23756 30243 23808 30252
rect 23756 30209 23765 30243
rect 23765 30209 23799 30243
rect 23799 30209 23808 30243
rect 23756 30200 23808 30209
rect 26148 30200 26200 30252
rect 19340 29996 19392 30048
rect 19616 30039 19668 30048
rect 19616 30005 19625 30039
rect 19625 30005 19659 30039
rect 19659 30005 19668 30039
rect 19616 29996 19668 30005
rect 20076 29996 20128 30048
rect 22100 29996 22152 30048
rect 22468 29996 22520 30048
rect 22652 30064 22704 30116
rect 23940 30175 23992 30184
rect 23940 30141 23949 30175
rect 23949 30141 23983 30175
rect 23983 30141 23992 30175
rect 23940 30132 23992 30141
rect 22928 29996 22980 30048
rect 23204 29996 23256 30048
rect 26240 30132 26292 30184
rect 26608 30200 26660 30252
rect 27344 30200 27396 30252
rect 28080 30268 28132 30320
rect 28264 30268 28316 30320
rect 28448 30200 28500 30252
rect 28172 30132 28224 30184
rect 28264 30132 28316 30184
rect 27896 30064 27948 30116
rect 28080 30064 28132 30116
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 28908 30243 28960 30252
rect 28908 30209 28917 30243
rect 28917 30209 28951 30243
rect 28951 30209 28960 30243
rect 28908 30200 28960 30209
rect 29000 30243 29052 30252
rect 29000 30209 29009 30243
rect 29009 30209 29043 30243
rect 29043 30209 29052 30243
rect 29000 30200 29052 30209
rect 29368 30200 29420 30252
rect 29552 30243 29604 30252
rect 29552 30209 29561 30243
rect 29561 30209 29595 30243
rect 29595 30209 29604 30243
rect 29552 30200 29604 30209
rect 30012 30268 30064 30320
rect 30196 30200 30248 30252
rect 29184 30132 29236 30184
rect 30656 30243 30708 30252
rect 30656 30209 30665 30243
rect 30665 30209 30699 30243
rect 30699 30209 30708 30243
rect 30656 30200 30708 30209
rect 31116 30200 31168 30252
rect 31484 30200 31536 30252
rect 33048 30243 33100 30252
rect 33048 30209 33057 30243
rect 33057 30209 33091 30243
rect 33091 30209 33100 30243
rect 33048 30200 33100 30209
rect 33324 30243 33376 30252
rect 33324 30209 33333 30243
rect 33333 30209 33367 30243
rect 33367 30209 33376 30243
rect 33324 30200 33376 30209
rect 33416 30243 33468 30252
rect 33416 30209 33425 30243
rect 33425 30209 33459 30243
rect 33459 30209 33468 30243
rect 33416 30200 33468 30209
rect 32404 30132 32456 30184
rect 34428 30243 34480 30252
rect 34428 30209 34437 30243
rect 34437 30209 34471 30243
rect 34471 30209 34480 30243
rect 34428 30200 34480 30209
rect 30472 30107 30524 30116
rect 26884 29996 26936 30048
rect 27436 29996 27488 30048
rect 28540 29996 28592 30048
rect 30472 30073 30481 30107
rect 30481 30073 30515 30107
rect 30515 30073 30524 30107
rect 30472 30064 30524 30073
rect 28908 29996 28960 30048
rect 29644 29996 29696 30048
rect 30564 29996 30616 30048
rect 31576 29996 31628 30048
rect 34336 30132 34388 30184
rect 33232 30064 33284 30116
rect 33600 29996 33652 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1308 29792 1360 29844
rect 3608 29792 3660 29844
rect 3976 29792 4028 29844
rect 8944 29792 8996 29844
rect 9220 29792 9272 29844
rect 10416 29792 10468 29844
rect 10508 29792 10560 29844
rect 10968 29792 11020 29844
rect 15476 29792 15528 29844
rect 3148 29656 3200 29708
rect 3240 29699 3292 29708
rect 3240 29665 3249 29699
rect 3249 29665 3283 29699
rect 3283 29665 3292 29699
rect 3240 29656 3292 29665
rect 3700 29656 3752 29708
rect 4068 29588 4120 29640
rect 6276 29656 6328 29708
rect 7104 29656 7156 29708
rect 5540 29588 5592 29640
rect 5632 29631 5684 29640
rect 5632 29597 5641 29631
rect 5641 29597 5675 29631
rect 5675 29597 5684 29631
rect 5632 29588 5684 29597
rect 5816 29588 5868 29640
rect 6552 29588 6604 29640
rect 7564 29588 7616 29640
rect 8392 29656 8444 29708
rect 8116 29631 8168 29640
rect 8116 29597 8125 29631
rect 8125 29597 8159 29631
rect 8159 29597 8168 29631
rect 8116 29588 8168 29597
rect 8668 29588 8720 29640
rect 5356 29520 5408 29572
rect 3056 29452 3108 29504
rect 4712 29452 4764 29504
rect 5172 29495 5224 29504
rect 5172 29461 5181 29495
rect 5181 29461 5215 29495
rect 5215 29461 5224 29495
rect 5172 29452 5224 29461
rect 5724 29495 5776 29504
rect 5724 29461 5733 29495
rect 5733 29461 5767 29495
rect 5767 29461 5776 29495
rect 5724 29452 5776 29461
rect 9128 29724 9180 29776
rect 9772 29656 9824 29708
rect 9312 29588 9364 29640
rect 11612 29656 11664 29708
rect 13084 29724 13136 29776
rect 13360 29724 13412 29776
rect 10416 29588 10468 29640
rect 10600 29588 10652 29640
rect 10784 29588 10836 29640
rect 11796 29631 11848 29640
rect 11796 29597 11805 29631
rect 11805 29597 11839 29631
rect 11839 29597 11848 29631
rect 11796 29588 11848 29597
rect 12256 29631 12308 29640
rect 12256 29597 12265 29631
rect 12265 29597 12299 29631
rect 12299 29597 12308 29631
rect 12256 29588 12308 29597
rect 12624 29631 12676 29640
rect 12624 29597 12633 29631
rect 12633 29597 12667 29631
rect 12667 29597 12676 29631
rect 12624 29588 12676 29597
rect 9220 29452 9272 29504
rect 13636 29588 13688 29640
rect 16028 29724 16080 29776
rect 17316 29792 17368 29844
rect 18604 29835 18656 29844
rect 18604 29801 18613 29835
rect 18613 29801 18647 29835
rect 18647 29801 18656 29835
rect 18604 29792 18656 29801
rect 18972 29792 19024 29844
rect 14096 29699 14148 29708
rect 14096 29665 14105 29699
rect 14105 29665 14139 29699
rect 14139 29665 14148 29699
rect 14096 29656 14148 29665
rect 13820 29631 13872 29640
rect 13820 29597 13829 29631
rect 13829 29597 13863 29631
rect 13863 29597 13872 29631
rect 13820 29588 13872 29597
rect 14372 29631 14424 29640
rect 14372 29597 14381 29631
rect 14381 29597 14415 29631
rect 14415 29597 14424 29631
rect 14372 29588 14424 29597
rect 15292 29699 15344 29708
rect 15292 29665 15301 29699
rect 15301 29665 15335 29699
rect 15335 29665 15344 29699
rect 15292 29656 15344 29665
rect 16580 29699 16632 29708
rect 16580 29665 16589 29699
rect 16589 29665 16623 29699
rect 16623 29665 16632 29699
rect 16580 29656 16632 29665
rect 15752 29588 15804 29640
rect 17408 29656 17460 29708
rect 18328 29724 18380 29776
rect 18788 29724 18840 29776
rect 23940 29792 23992 29844
rect 19708 29724 19760 29776
rect 20168 29724 20220 29776
rect 21272 29724 21324 29776
rect 21548 29724 21600 29776
rect 22100 29767 22152 29776
rect 22100 29733 22109 29767
rect 22109 29733 22143 29767
rect 22143 29733 22152 29767
rect 22100 29724 22152 29733
rect 22192 29767 22244 29776
rect 22192 29733 22201 29767
rect 22201 29733 22235 29767
rect 22235 29733 22244 29767
rect 22192 29724 22244 29733
rect 22284 29724 22336 29776
rect 14004 29520 14056 29572
rect 9496 29452 9548 29504
rect 10232 29452 10284 29504
rect 13176 29452 13228 29504
rect 13268 29452 13320 29504
rect 13360 29452 13412 29504
rect 13636 29452 13688 29504
rect 15568 29520 15620 29572
rect 16212 29563 16264 29572
rect 16212 29529 16221 29563
rect 16221 29529 16255 29563
rect 16255 29529 16264 29563
rect 16212 29520 16264 29529
rect 17040 29588 17092 29640
rect 17684 29588 17736 29640
rect 17960 29588 18012 29640
rect 18512 29631 18564 29640
rect 18512 29597 18521 29631
rect 18521 29597 18555 29631
rect 18555 29597 18564 29631
rect 18512 29588 18564 29597
rect 19708 29631 19760 29640
rect 19708 29597 19717 29631
rect 19717 29597 19751 29631
rect 19751 29597 19760 29631
rect 19708 29588 19760 29597
rect 15844 29452 15896 29504
rect 16120 29452 16172 29504
rect 16672 29452 16724 29504
rect 16764 29495 16816 29504
rect 16764 29461 16773 29495
rect 16773 29461 16807 29495
rect 16807 29461 16816 29495
rect 16764 29452 16816 29461
rect 17776 29520 17828 29572
rect 17868 29520 17920 29572
rect 17040 29452 17092 29504
rect 17960 29452 18012 29504
rect 18236 29495 18288 29504
rect 18236 29461 18245 29495
rect 18245 29461 18279 29495
rect 18279 29461 18288 29495
rect 18236 29452 18288 29461
rect 18420 29520 18472 29572
rect 19616 29520 19668 29572
rect 20812 29631 20864 29640
rect 20812 29597 20821 29631
rect 20821 29597 20855 29631
rect 20855 29597 20864 29631
rect 20812 29588 20864 29597
rect 20904 29631 20956 29640
rect 20904 29597 20913 29631
rect 20913 29597 20947 29631
rect 20947 29597 20956 29631
rect 20904 29588 20956 29597
rect 20996 29631 21048 29640
rect 20996 29597 21005 29631
rect 21005 29597 21039 29631
rect 21039 29597 21048 29631
rect 20996 29588 21048 29597
rect 21272 29588 21324 29640
rect 21456 29520 21508 29572
rect 22008 29656 22060 29708
rect 21732 29588 21784 29640
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 22836 29631 22888 29640
rect 22836 29597 22845 29631
rect 22845 29597 22879 29631
rect 22879 29597 22888 29631
rect 22836 29588 22888 29597
rect 23296 29631 23348 29640
rect 23296 29597 23305 29631
rect 23305 29597 23339 29631
rect 23339 29597 23348 29631
rect 23296 29588 23348 29597
rect 24492 29724 24544 29776
rect 26148 29724 26200 29776
rect 26332 29792 26384 29844
rect 27160 29792 27212 29844
rect 28448 29792 28500 29844
rect 28908 29792 28960 29844
rect 29184 29792 29236 29844
rect 29828 29792 29880 29844
rect 32036 29792 32088 29844
rect 26976 29656 27028 29708
rect 27528 29699 27580 29708
rect 27528 29665 27537 29699
rect 27537 29665 27571 29699
rect 27571 29665 27580 29699
rect 27528 29656 27580 29665
rect 28540 29724 28592 29776
rect 29000 29724 29052 29776
rect 29092 29724 29144 29776
rect 28908 29656 28960 29708
rect 25780 29631 25832 29640
rect 25780 29597 25789 29631
rect 25789 29597 25823 29631
rect 25823 29597 25832 29631
rect 25780 29588 25832 29597
rect 26792 29588 26844 29640
rect 26884 29631 26936 29640
rect 26884 29597 26893 29631
rect 26893 29597 26927 29631
rect 26927 29597 26936 29631
rect 26884 29588 26936 29597
rect 27068 29631 27120 29640
rect 27068 29597 27077 29631
rect 27077 29597 27111 29631
rect 27111 29597 27120 29631
rect 27068 29588 27120 29597
rect 27344 29588 27396 29640
rect 27712 29588 27764 29640
rect 28264 29631 28316 29640
rect 28264 29597 28273 29631
rect 28273 29597 28307 29631
rect 28307 29597 28316 29631
rect 28264 29588 28316 29597
rect 28448 29588 28500 29640
rect 30472 29588 30524 29640
rect 23664 29520 23716 29572
rect 25228 29563 25280 29572
rect 25228 29529 25237 29563
rect 25237 29529 25271 29563
rect 25271 29529 25280 29563
rect 25228 29520 25280 29529
rect 20996 29452 21048 29504
rect 21640 29452 21692 29504
rect 23020 29452 23072 29504
rect 25688 29452 25740 29504
rect 26148 29520 26200 29572
rect 26608 29563 26660 29572
rect 26608 29529 26617 29563
rect 26617 29529 26651 29563
rect 26651 29529 26660 29563
rect 26608 29520 26660 29529
rect 27528 29520 27580 29572
rect 30288 29520 30340 29572
rect 30748 29520 30800 29572
rect 30840 29520 30892 29572
rect 32956 29588 33008 29640
rect 31944 29520 31996 29572
rect 27988 29495 28040 29504
rect 27988 29461 27997 29495
rect 27997 29461 28031 29495
rect 28031 29461 28040 29495
rect 27988 29452 28040 29461
rect 28172 29452 28224 29504
rect 28816 29452 28868 29504
rect 30932 29452 30984 29504
rect 31116 29452 31168 29504
rect 31484 29452 31536 29504
rect 31576 29495 31628 29504
rect 31576 29461 31585 29495
rect 31585 29461 31619 29495
rect 31619 29461 31628 29495
rect 31576 29452 31628 29461
rect 31852 29495 31904 29504
rect 31852 29461 31861 29495
rect 31861 29461 31895 29495
rect 31895 29461 31904 29495
rect 31852 29452 31904 29461
rect 32312 29495 32364 29504
rect 32312 29461 32321 29495
rect 32321 29461 32355 29495
rect 32355 29461 32364 29495
rect 32312 29452 32364 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 1308 29180 1360 29232
rect 7748 29248 7800 29300
rect 16028 29248 16080 29300
rect 3056 29180 3108 29232
rect 3608 29180 3660 29232
rect 4804 29180 4856 29232
rect 6460 29180 6512 29232
rect 7104 29223 7156 29232
rect 7104 29189 7113 29223
rect 7113 29189 7147 29223
rect 7147 29189 7156 29223
rect 7104 29180 7156 29189
rect 4068 29044 4120 29096
rect 7196 29155 7248 29164
rect 7196 29121 7205 29155
rect 7205 29121 7239 29155
rect 7239 29121 7248 29155
rect 7196 29112 7248 29121
rect 9404 29180 9456 29232
rect 10324 29180 10376 29232
rect 10692 29180 10744 29232
rect 14372 29180 14424 29232
rect 15292 29180 15344 29232
rect 16396 29180 16448 29232
rect 16764 29180 16816 29232
rect 7748 29155 7800 29164
rect 7748 29121 7757 29155
rect 7757 29121 7791 29155
rect 7791 29121 7800 29155
rect 7748 29112 7800 29121
rect 8668 29112 8720 29164
rect 9220 29112 9272 29164
rect 9588 29155 9640 29164
rect 9588 29121 9597 29155
rect 9597 29121 9631 29155
rect 9631 29121 9640 29155
rect 9588 29112 9640 29121
rect 9956 29155 10008 29164
rect 9956 29121 9965 29155
rect 9965 29121 9999 29155
rect 9999 29121 10008 29155
rect 9956 29112 10008 29121
rect 11796 29112 11848 29164
rect 12256 29112 12308 29164
rect 12716 29112 12768 29164
rect 12900 29155 12952 29164
rect 12900 29121 12909 29155
rect 12909 29121 12943 29155
rect 12943 29121 12952 29155
rect 12900 29112 12952 29121
rect 13268 29112 13320 29164
rect 7472 29087 7524 29096
rect 7472 29053 7481 29087
rect 7481 29053 7515 29087
rect 7515 29053 7524 29087
rect 7472 29044 7524 29053
rect 2412 28908 2464 28960
rect 5264 28908 5316 28960
rect 5356 28908 5408 28960
rect 7012 28976 7064 29028
rect 9404 29044 9456 29096
rect 11152 29044 11204 29096
rect 8116 28976 8168 29028
rect 10048 28976 10100 29028
rect 9588 28908 9640 28960
rect 11704 28908 11756 28960
rect 12440 28976 12492 29028
rect 12808 29044 12860 29096
rect 13176 29087 13228 29096
rect 13176 29053 13185 29087
rect 13185 29053 13219 29087
rect 13219 29053 13228 29087
rect 13176 29044 13228 29053
rect 13452 29087 13504 29096
rect 13452 29053 13461 29087
rect 13461 29053 13495 29087
rect 13495 29053 13504 29087
rect 13452 29044 13504 29053
rect 13636 29155 13688 29164
rect 13636 29121 13645 29155
rect 13645 29121 13679 29155
rect 13679 29121 13688 29155
rect 13636 29112 13688 29121
rect 13820 29044 13872 29096
rect 14188 29112 14240 29164
rect 14464 29155 14516 29164
rect 14464 29121 14473 29155
rect 14473 29121 14507 29155
rect 14507 29121 14516 29155
rect 14464 29112 14516 29121
rect 15752 29112 15804 29164
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 14372 29044 14424 29096
rect 15292 29087 15344 29096
rect 15292 29053 15301 29087
rect 15301 29053 15335 29087
rect 15335 29053 15344 29087
rect 15292 29044 15344 29053
rect 15476 29044 15528 29096
rect 15568 29087 15620 29096
rect 15568 29053 15577 29087
rect 15577 29053 15611 29087
rect 15611 29053 15620 29087
rect 15568 29044 15620 29053
rect 15660 29087 15712 29096
rect 15660 29053 15669 29087
rect 15669 29053 15703 29087
rect 15703 29053 15712 29087
rect 15660 29044 15712 29053
rect 15844 29044 15896 29096
rect 16212 29044 16264 29096
rect 17224 29112 17276 29164
rect 17776 29112 17828 29164
rect 18512 29248 18564 29300
rect 19064 29248 19116 29300
rect 18052 29112 18104 29164
rect 20260 29180 20312 29232
rect 18972 29112 19024 29164
rect 21640 29248 21692 29300
rect 21824 29248 21876 29300
rect 20628 29155 20680 29164
rect 20628 29121 20637 29155
rect 20637 29121 20671 29155
rect 20671 29121 20680 29155
rect 20628 29112 20680 29121
rect 20812 29155 20864 29164
rect 20812 29121 20821 29155
rect 20821 29121 20855 29155
rect 20855 29121 20864 29155
rect 20812 29112 20864 29121
rect 20996 29112 21048 29164
rect 21180 29155 21232 29164
rect 21180 29121 21189 29155
rect 21189 29121 21223 29155
rect 21223 29121 21232 29155
rect 21180 29112 21232 29121
rect 21456 29155 21508 29164
rect 21456 29121 21465 29155
rect 21465 29121 21499 29155
rect 21499 29121 21508 29155
rect 21456 29112 21508 29121
rect 21640 29112 21692 29164
rect 22652 29291 22704 29300
rect 22652 29257 22661 29291
rect 22661 29257 22695 29291
rect 22695 29257 22704 29291
rect 22652 29248 22704 29257
rect 22744 29248 22796 29300
rect 23388 29248 23440 29300
rect 22836 29155 22888 29164
rect 22836 29121 22845 29155
rect 22845 29121 22879 29155
rect 22879 29121 22888 29155
rect 22836 29112 22888 29121
rect 23296 29112 23348 29164
rect 24952 29248 25004 29300
rect 26608 29248 26660 29300
rect 26792 29248 26844 29300
rect 29184 29248 29236 29300
rect 32680 29248 32732 29300
rect 24492 29180 24544 29232
rect 28172 29180 28224 29232
rect 14280 29019 14332 29028
rect 14280 28985 14289 29019
rect 14289 28985 14323 29019
rect 14323 28985 14332 29019
rect 14280 28976 14332 28985
rect 14924 29019 14976 29028
rect 14924 28985 14933 29019
rect 14933 28985 14967 29019
rect 14967 28985 14976 29019
rect 14924 28976 14976 28985
rect 15384 29019 15436 29028
rect 15384 28985 15393 29019
rect 15393 28985 15427 29019
rect 15427 28985 15436 29019
rect 15384 28976 15436 28985
rect 17040 29087 17092 29096
rect 17040 29053 17049 29087
rect 17049 29053 17083 29087
rect 17083 29053 17092 29087
rect 17040 29044 17092 29053
rect 17224 28976 17276 29028
rect 17684 29044 17736 29096
rect 14832 28908 14884 28960
rect 16580 28908 16632 28960
rect 18052 28976 18104 29028
rect 20168 28976 20220 29028
rect 21364 29019 21416 29028
rect 21364 28985 21373 29019
rect 21373 28985 21407 29019
rect 21407 28985 21416 29019
rect 21364 28976 21416 28985
rect 22284 29044 22336 29096
rect 22928 29044 22980 29096
rect 23204 28976 23256 29028
rect 23296 28976 23348 29028
rect 21824 28951 21876 28960
rect 21824 28917 21833 28951
rect 21833 28917 21867 28951
rect 21867 28917 21876 28951
rect 21824 28908 21876 28917
rect 21916 28908 21968 28960
rect 23388 28908 23440 28960
rect 26148 29112 26200 29164
rect 26700 29112 26752 29164
rect 27528 29155 27580 29164
rect 27528 29121 27537 29155
rect 27537 29121 27571 29155
rect 27571 29121 27580 29155
rect 27528 29112 27580 29121
rect 27804 29112 27856 29164
rect 28264 29155 28316 29164
rect 28264 29121 28273 29155
rect 28273 29121 28307 29155
rect 28307 29121 28316 29155
rect 28264 29112 28316 29121
rect 25596 29044 25648 29096
rect 26608 29044 26660 29096
rect 26884 29044 26936 29096
rect 29000 29112 29052 29164
rect 29552 29155 29604 29164
rect 29552 29121 29561 29155
rect 29561 29121 29595 29155
rect 29595 29121 29604 29155
rect 29552 29112 29604 29121
rect 30380 29223 30432 29232
rect 30380 29189 30389 29223
rect 30389 29189 30423 29223
rect 30423 29189 30432 29223
rect 30380 29180 30432 29189
rect 30748 29223 30800 29232
rect 30748 29189 30757 29223
rect 30757 29189 30791 29223
rect 30791 29189 30800 29223
rect 30748 29180 30800 29189
rect 30932 29180 30984 29232
rect 30656 29155 30708 29164
rect 30656 29121 30665 29155
rect 30665 29121 30699 29155
rect 30699 29121 30708 29155
rect 30656 29112 30708 29121
rect 27712 28976 27764 29028
rect 28448 29019 28500 29028
rect 28448 28985 28457 29019
rect 28457 28985 28491 29019
rect 28491 28985 28500 29019
rect 28448 28976 28500 28985
rect 26516 28908 26568 28960
rect 26884 28908 26936 28960
rect 28080 28951 28132 28960
rect 28080 28917 28089 28951
rect 28089 28917 28123 28951
rect 28123 28917 28132 28951
rect 28080 28908 28132 28917
rect 28540 28908 28592 28960
rect 30012 29019 30064 29028
rect 30012 28985 30021 29019
rect 30021 28985 30055 29019
rect 30055 28985 30064 29019
rect 30012 28976 30064 28985
rect 30472 29044 30524 29096
rect 31484 29112 31536 29164
rect 36176 29180 36228 29232
rect 31668 29112 31720 29164
rect 33784 29112 33836 29164
rect 35808 29155 35860 29164
rect 35808 29121 35817 29155
rect 35817 29121 35851 29155
rect 35851 29121 35860 29155
rect 35808 29112 35860 29121
rect 31944 28976 31996 29028
rect 30656 28908 30708 28960
rect 30840 28908 30892 28960
rect 34520 29044 34572 29096
rect 34796 29044 34848 29096
rect 35624 29019 35676 29028
rect 35624 28985 35633 29019
rect 35633 28985 35667 29019
rect 35667 28985 35676 29019
rect 35624 28976 35676 28985
rect 35808 28908 35860 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1308 28568 1360 28620
rect 3608 28611 3660 28620
rect 3608 28577 3617 28611
rect 3617 28577 3651 28611
rect 3651 28577 3660 28611
rect 3608 28568 3660 28577
rect 5816 28704 5868 28756
rect 6920 28704 6972 28756
rect 8576 28704 8628 28756
rect 9956 28704 10008 28756
rect 10140 28704 10192 28756
rect 11152 28704 11204 28756
rect 15016 28704 15068 28756
rect 15292 28704 15344 28756
rect 15752 28747 15804 28756
rect 15752 28713 15761 28747
rect 15761 28713 15795 28747
rect 15795 28713 15804 28747
rect 15752 28704 15804 28713
rect 16488 28704 16540 28756
rect 19248 28704 19300 28756
rect 21180 28704 21232 28756
rect 22284 28747 22336 28756
rect 22284 28713 22293 28747
rect 22293 28713 22327 28747
rect 22327 28713 22336 28747
rect 22284 28704 22336 28713
rect 5356 28568 5408 28620
rect 6276 28679 6328 28688
rect 6276 28645 6285 28679
rect 6285 28645 6319 28679
rect 6319 28645 6328 28679
rect 6276 28636 6328 28645
rect 7104 28636 7156 28688
rect 7472 28636 7524 28688
rect 2780 28432 2832 28484
rect 4068 28432 4120 28484
rect 5264 28432 5316 28484
rect 5724 28543 5776 28552
rect 5724 28509 5733 28543
rect 5733 28509 5767 28543
rect 5767 28509 5776 28543
rect 5724 28500 5776 28509
rect 7564 28611 7616 28620
rect 7564 28577 7573 28611
rect 7573 28577 7607 28611
rect 7607 28577 7616 28611
rect 7564 28568 7616 28577
rect 7748 28636 7800 28688
rect 9220 28636 9272 28688
rect 7932 28611 7984 28620
rect 7932 28577 7941 28611
rect 7941 28577 7975 28611
rect 7975 28577 7984 28611
rect 7932 28568 7984 28577
rect 6460 28543 6512 28552
rect 6460 28509 6469 28543
rect 6469 28509 6503 28543
rect 6503 28509 6512 28543
rect 6460 28500 6512 28509
rect 7012 28500 7064 28552
rect 7288 28543 7340 28552
rect 7288 28509 7297 28543
rect 7297 28509 7331 28543
rect 7331 28509 7340 28543
rect 7288 28500 7340 28509
rect 7380 28543 7432 28552
rect 7380 28509 7389 28543
rect 7389 28509 7423 28543
rect 7423 28509 7432 28543
rect 7380 28500 7432 28509
rect 7932 28432 7984 28484
rect 8668 28500 8720 28552
rect 9220 28543 9272 28552
rect 9220 28509 9229 28543
rect 9229 28509 9263 28543
rect 9263 28509 9272 28543
rect 9220 28500 9272 28509
rect 9404 28543 9456 28552
rect 9404 28509 9413 28543
rect 9413 28509 9447 28543
rect 9447 28509 9456 28543
rect 9404 28500 9456 28509
rect 9772 28636 9824 28688
rect 10232 28636 10284 28688
rect 10324 28636 10376 28688
rect 15200 28636 15252 28688
rect 16856 28636 16908 28688
rect 9680 28543 9732 28552
rect 9680 28509 9689 28543
rect 9689 28509 9723 28543
rect 9723 28509 9732 28543
rect 9680 28500 9732 28509
rect 9772 28543 9824 28552
rect 9772 28509 9781 28543
rect 9781 28509 9815 28543
rect 9815 28509 9824 28543
rect 9772 28500 9824 28509
rect 10324 28543 10376 28552
rect 10324 28509 10333 28543
rect 10333 28509 10367 28543
rect 10367 28509 10376 28543
rect 10324 28500 10376 28509
rect 10600 28500 10652 28552
rect 12716 28568 12768 28620
rect 12900 28611 12952 28620
rect 12900 28577 12909 28611
rect 12909 28577 12943 28611
rect 12943 28577 12952 28611
rect 12900 28568 12952 28577
rect 10968 28500 11020 28552
rect 11796 28500 11848 28552
rect 4804 28364 4856 28416
rect 6736 28407 6788 28416
rect 6736 28373 6745 28407
rect 6745 28373 6779 28407
rect 6779 28373 6788 28407
rect 6736 28364 6788 28373
rect 7288 28364 7340 28416
rect 9128 28364 9180 28416
rect 9312 28407 9364 28416
rect 9312 28373 9321 28407
rect 9321 28373 9355 28407
rect 9355 28373 9364 28407
rect 9312 28364 9364 28373
rect 10232 28432 10284 28484
rect 12348 28543 12400 28552
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 13084 28500 13136 28552
rect 13268 28500 13320 28552
rect 13544 28500 13596 28552
rect 13728 28543 13780 28552
rect 13728 28509 13737 28543
rect 13737 28509 13771 28543
rect 13771 28509 13780 28543
rect 13728 28500 13780 28509
rect 12164 28432 12216 28484
rect 13176 28432 13228 28484
rect 10876 28364 10928 28416
rect 10968 28407 11020 28416
rect 10968 28373 10977 28407
rect 10977 28373 11011 28407
rect 11011 28373 11020 28407
rect 10968 28364 11020 28373
rect 11704 28407 11756 28416
rect 11704 28373 11713 28407
rect 11713 28373 11747 28407
rect 11747 28373 11756 28407
rect 11704 28364 11756 28373
rect 11796 28364 11848 28416
rect 14188 28432 14240 28484
rect 15016 28500 15068 28552
rect 15384 28543 15436 28552
rect 15384 28509 15393 28543
rect 15393 28509 15427 28543
rect 15427 28509 15436 28543
rect 15384 28500 15436 28509
rect 15568 28543 15620 28552
rect 15568 28509 15577 28543
rect 15577 28509 15611 28543
rect 15611 28509 15620 28543
rect 15568 28500 15620 28509
rect 15660 28500 15712 28552
rect 16028 28543 16080 28552
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 16764 28568 16816 28620
rect 16396 28543 16448 28552
rect 16396 28509 16405 28543
rect 16405 28509 16439 28543
rect 16439 28509 16448 28543
rect 16396 28500 16448 28509
rect 16580 28543 16632 28552
rect 16580 28509 16589 28543
rect 16589 28509 16623 28543
rect 16623 28509 16632 28543
rect 16580 28500 16632 28509
rect 16672 28500 16724 28552
rect 18604 28568 18656 28620
rect 20720 28568 20772 28620
rect 22560 28636 22612 28688
rect 22836 28636 22888 28688
rect 22468 28611 22520 28620
rect 18788 28543 18840 28552
rect 18788 28509 18797 28543
rect 18797 28509 18831 28543
rect 18831 28509 18840 28543
rect 18788 28500 18840 28509
rect 18972 28543 19024 28552
rect 18972 28509 18981 28543
rect 18981 28509 19015 28543
rect 19015 28509 19024 28543
rect 18972 28500 19024 28509
rect 20260 28500 20312 28552
rect 20536 28543 20588 28552
rect 20536 28509 20545 28543
rect 20545 28509 20579 28543
rect 20579 28509 20588 28543
rect 20536 28500 20588 28509
rect 20996 28500 21048 28552
rect 21088 28543 21140 28552
rect 21088 28509 21097 28543
rect 21097 28509 21131 28543
rect 21131 28509 21140 28543
rect 21088 28500 21140 28509
rect 21364 28543 21416 28552
rect 21364 28509 21373 28543
rect 21373 28509 21407 28543
rect 21407 28509 21416 28543
rect 21364 28500 21416 28509
rect 13912 28364 13964 28416
rect 17132 28432 17184 28484
rect 17408 28432 17460 28484
rect 20168 28432 20220 28484
rect 22468 28577 22477 28611
rect 22477 28577 22511 28611
rect 22511 28577 22520 28611
rect 22468 28568 22520 28577
rect 22652 28568 22704 28620
rect 24400 28704 24452 28756
rect 25596 28704 25648 28756
rect 26700 28704 26752 28756
rect 27068 28704 27120 28756
rect 27712 28704 27764 28756
rect 28264 28747 28316 28756
rect 28264 28713 28273 28747
rect 28273 28713 28307 28747
rect 28307 28713 28316 28747
rect 28264 28704 28316 28713
rect 29552 28704 29604 28756
rect 29920 28704 29972 28756
rect 34888 28704 34940 28756
rect 24584 28636 24636 28688
rect 24768 28636 24820 28688
rect 25136 28636 25188 28688
rect 25780 28636 25832 28688
rect 24492 28568 24544 28620
rect 23020 28500 23072 28552
rect 15568 28364 15620 28416
rect 16396 28364 16448 28416
rect 16580 28364 16632 28416
rect 18880 28407 18932 28416
rect 18880 28373 18889 28407
rect 18889 28373 18923 28407
rect 18923 28373 18932 28407
rect 18880 28364 18932 28373
rect 20812 28364 20864 28416
rect 21364 28407 21416 28416
rect 21364 28373 21373 28407
rect 21373 28373 21407 28407
rect 21407 28373 21416 28407
rect 21364 28364 21416 28373
rect 21732 28364 21784 28416
rect 22376 28432 22428 28484
rect 23572 28432 23624 28484
rect 24860 28500 24912 28552
rect 24952 28543 25004 28552
rect 24952 28509 24961 28543
rect 24961 28509 24995 28543
rect 24995 28509 25004 28543
rect 24952 28500 25004 28509
rect 25044 28500 25096 28552
rect 25688 28568 25740 28620
rect 26700 28568 26752 28620
rect 26516 28543 26568 28552
rect 26516 28509 26525 28543
rect 26525 28509 26559 28543
rect 26559 28509 26568 28543
rect 26516 28500 26568 28509
rect 26608 28543 26660 28552
rect 26608 28509 26617 28543
rect 26617 28509 26651 28543
rect 26651 28509 26660 28543
rect 26608 28500 26660 28509
rect 24768 28432 24820 28484
rect 22192 28364 22244 28416
rect 23204 28364 23256 28416
rect 23756 28407 23808 28416
rect 23756 28373 23791 28407
rect 23791 28373 23808 28407
rect 23756 28364 23808 28373
rect 24124 28364 24176 28416
rect 24676 28364 24728 28416
rect 26332 28432 26384 28484
rect 27528 28568 27580 28620
rect 28080 28636 28132 28688
rect 28632 28636 28684 28688
rect 28908 28636 28960 28688
rect 27620 28500 27672 28552
rect 27252 28475 27304 28484
rect 27252 28441 27261 28475
rect 27261 28441 27295 28475
rect 27295 28441 27304 28475
rect 27252 28432 27304 28441
rect 27344 28475 27396 28484
rect 27344 28441 27353 28475
rect 27353 28441 27387 28475
rect 27387 28441 27396 28475
rect 27344 28432 27396 28441
rect 28816 28611 28868 28620
rect 28816 28577 28825 28611
rect 28825 28577 28859 28611
rect 28859 28577 28868 28611
rect 28816 28568 28868 28577
rect 30104 28568 30156 28620
rect 28264 28543 28316 28552
rect 28264 28509 28273 28543
rect 28273 28509 28307 28543
rect 28307 28509 28316 28543
rect 28264 28500 28316 28509
rect 28724 28500 28776 28552
rect 28632 28432 28684 28484
rect 29552 28432 29604 28484
rect 29920 28500 29972 28552
rect 30196 28500 30248 28552
rect 29828 28432 29880 28484
rect 28448 28364 28500 28416
rect 30840 28364 30892 28416
rect 31668 28364 31720 28416
rect 31852 28475 31904 28484
rect 31852 28441 31861 28475
rect 31861 28441 31895 28475
rect 31895 28441 31904 28475
rect 31852 28432 31904 28441
rect 32680 28568 32732 28620
rect 33324 28636 33376 28688
rect 34428 28636 34480 28688
rect 34796 28568 34848 28620
rect 32036 28543 32088 28552
rect 32036 28509 32071 28543
rect 32071 28509 32088 28543
rect 32036 28500 32088 28509
rect 33784 28543 33836 28552
rect 33784 28509 33793 28543
rect 33793 28509 33827 28543
rect 33827 28509 33836 28543
rect 33784 28500 33836 28509
rect 34704 28432 34756 28484
rect 34612 28364 34664 28416
rect 35624 28432 35676 28484
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 2780 28160 2832 28212
rect 3516 28160 3568 28212
rect 5724 28160 5776 28212
rect 7196 28160 7248 28212
rect 3424 28067 3476 28076
rect 3424 28033 3433 28067
rect 3433 28033 3467 28067
rect 3467 28033 3476 28067
rect 3424 28024 3476 28033
rect 3608 28024 3660 28076
rect 6000 28092 6052 28144
rect 6920 28135 6972 28144
rect 6920 28101 6929 28135
rect 6929 28101 6963 28135
rect 6963 28101 6972 28135
rect 6920 28092 6972 28101
rect 7012 28092 7064 28144
rect 5264 28024 5316 28076
rect 5908 28024 5960 28076
rect 6736 28024 6788 28076
rect 1400 27999 1452 28008
rect 1400 27965 1409 27999
rect 1409 27965 1443 27999
rect 1443 27965 1452 27999
rect 1400 27956 1452 27965
rect 3148 27999 3200 28008
rect 3148 27965 3157 27999
rect 3157 27965 3191 27999
rect 3191 27965 3200 27999
rect 3148 27956 3200 27965
rect 4988 27956 5040 28008
rect 7196 27999 7248 28008
rect 7196 27965 7205 27999
rect 7205 27965 7239 27999
rect 7239 27965 7248 27999
rect 7196 27956 7248 27965
rect 7748 28092 7800 28144
rect 9680 28160 9732 28212
rect 9772 28160 9824 28212
rect 10416 28160 10468 28212
rect 13176 28203 13228 28212
rect 13176 28169 13185 28203
rect 13185 28169 13219 28203
rect 13219 28169 13228 28203
rect 13176 28160 13228 28169
rect 15384 28160 15436 28212
rect 17868 28160 17920 28212
rect 8116 28024 8168 28076
rect 9312 28092 9364 28144
rect 8852 28067 8904 28076
rect 8852 28033 8861 28067
rect 8861 28033 8895 28067
rect 8895 28033 8904 28067
rect 8852 28024 8904 28033
rect 9036 28024 9088 28076
rect 9220 28067 9272 28076
rect 9220 28033 9229 28067
rect 9229 28033 9263 28067
rect 9263 28033 9272 28067
rect 9220 28024 9272 28033
rect 9588 28024 9640 28076
rect 9772 28024 9824 28076
rect 10968 28092 11020 28144
rect 11704 28092 11756 28144
rect 2504 27820 2556 27872
rect 4620 27820 4672 27872
rect 5264 27888 5316 27940
rect 8024 27956 8076 28008
rect 9680 27956 9732 28008
rect 10232 28067 10284 28076
rect 10232 28033 10241 28067
rect 10241 28033 10275 28067
rect 10275 28033 10284 28067
rect 10232 28024 10284 28033
rect 10324 28024 10376 28076
rect 10600 28067 10652 28076
rect 10600 28033 10609 28067
rect 10609 28033 10643 28067
rect 10643 28033 10652 28067
rect 10600 28024 10652 28033
rect 10784 28024 10836 28076
rect 11244 28067 11296 28076
rect 11244 28033 11253 28067
rect 11253 28033 11287 28067
rect 11287 28033 11296 28067
rect 11244 28024 11296 28033
rect 12256 28024 12308 28076
rect 12348 28067 12400 28076
rect 12348 28033 12357 28067
rect 12357 28033 12391 28067
rect 12391 28033 12400 28067
rect 12348 28024 12400 28033
rect 13084 28092 13136 28144
rect 18236 28092 18288 28144
rect 19156 28160 19208 28212
rect 19248 28160 19300 28212
rect 21824 28160 21876 28212
rect 24584 28160 24636 28212
rect 25136 28203 25188 28212
rect 25136 28169 25145 28203
rect 25145 28169 25179 28203
rect 25179 28169 25188 28203
rect 25136 28160 25188 28169
rect 26516 28160 26568 28212
rect 13544 28067 13596 28076
rect 13544 28033 13553 28067
rect 13553 28033 13587 28067
rect 13587 28033 13596 28067
rect 13544 28024 13596 28033
rect 14464 28024 14516 28076
rect 14832 28024 14884 28076
rect 15476 28067 15528 28076
rect 15476 28033 15485 28067
rect 15485 28033 15519 28067
rect 15519 28033 15528 28067
rect 15476 28024 15528 28033
rect 16304 28024 16356 28076
rect 16672 28024 16724 28076
rect 16948 28024 17000 28076
rect 17316 28067 17368 28076
rect 17316 28033 17325 28067
rect 17325 28033 17359 28067
rect 17359 28033 17368 28067
rect 17316 28024 17368 28033
rect 17500 28024 17552 28076
rect 17684 28024 17736 28076
rect 13452 27956 13504 28008
rect 13728 27956 13780 28008
rect 15660 27956 15712 28008
rect 16488 27956 16540 28008
rect 19156 28024 19208 28076
rect 20904 28092 20956 28144
rect 21180 28135 21232 28144
rect 21180 28101 21189 28135
rect 21189 28101 21223 28135
rect 21223 28101 21232 28135
rect 21180 28092 21232 28101
rect 22192 28135 22244 28144
rect 22192 28101 22201 28135
rect 22201 28101 22235 28135
rect 22235 28101 22244 28135
rect 22192 28092 22244 28101
rect 23756 28092 23808 28144
rect 25044 28092 25096 28144
rect 26424 28135 26476 28144
rect 26424 28101 26433 28135
rect 26433 28101 26467 28135
rect 26467 28101 26476 28135
rect 26424 28092 26476 28101
rect 27344 28160 27396 28212
rect 27528 28160 27580 28212
rect 27620 28203 27672 28212
rect 27620 28169 27629 28203
rect 27629 28169 27663 28203
rect 27663 28169 27672 28203
rect 27620 28160 27672 28169
rect 27712 28160 27764 28212
rect 19432 27956 19484 28008
rect 19524 27999 19576 28008
rect 19524 27965 19533 27999
rect 19533 27965 19567 27999
rect 19567 27965 19576 27999
rect 19524 27956 19576 27965
rect 21916 27956 21968 28008
rect 10048 27888 10100 27940
rect 11060 27888 11112 27940
rect 11520 27931 11572 27940
rect 11520 27897 11529 27931
rect 11529 27897 11563 27931
rect 11563 27897 11572 27931
rect 11520 27888 11572 27897
rect 18972 27888 19024 27940
rect 19616 27888 19668 27940
rect 19984 27888 20036 27940
rect 22376 28067 22428 28076
rect 22376 28033 22385 28067
rect 22385 28033 22419 28067
rect 22419 28033 22428 28067
rect 22376 28024 22428 28033
rect 22928 28067 22980 28076
rect 22928 28033 22937 28067
rect 22937 28033 22971 28067
rect 22971 28033 22980 28067
rect 22928 28024 22980 28033
rect 23112 28067 23164 28076
rect 23112 28033 23121 28067
rect 23121 28033 23155 28067
rect 23155 28033 23164 28067
rect 23112 28024 23164 28033
rect 23388 28067 23440 28076
rect 23388 28033 23397 28067
rect 23397 28033 23431 28067
rect 23431 28033 23440 28067
rect 23388 28024 23440 28033
rect 24768 28024 24820 28076
rect 26240 28024 26292 28076
rect 26884 28092 26936 28144
rect 28264 28092 28316 28144
rect 30012 28135 30064 28144
rect 30012 28101 30021 28135
rect 30021 28101 30055 28135
rect 30055 28101 30064 28135
rect 36360 28160 36412 28212
rect 30012 28092 30064 28101
rect 27068 28024 27120 28076
rect 22836 27999 22888 28008
rect 22836 27965 22845 27999
rect 22845 27965 22879 27999
rect 22879 27965 22888 27999
rect 22836 27956 22888 27965
rect 22928 27888 22980 27940
rect 7840 27820 7892 27872
rect 8116 27820 8168 27872
rect 9588 27820 9640 27872
rect 9680 27820 9732 27872
rect 10784 27863 10836 27872
rect 10784 27829 10793 27863
rect 10793 27829 10827 27863
rect 10827 27829 10836 27863
rect 10784 27820 10836 27829
rect 11612 27820 11664 27872
rect 12900 27820 12952 27872
rect 17960 27820 18012 27872
rect 20996 27863 21048 27872
rect 20996 27829 21005 27863
rect 21005 27829 21039 27863
rect 21039 27829 21048 27863
rect 20996 27820 21048 27829
rect 22560 27863 22612 27872
rect 22560 27829 22569 27863
rect 22569 27829 22603 27863
rect 22603 27829 22612 27863
rect 22560 27820 22612 27829
rect 22652 27863 22704 27872
rect 22652 27829 22661 27863
rect 22661 27829 22695 27863
rect 22695 27829 22704 27863
rect 22652 27820 22704 27829
rect 23296 27956 23348 28008
rect 24676 27956 24728 28008
rect 26332 27956 26384 28008
rect 25872 27888 25924 27940
rect 26976 27888 27028 27940
rect 28448 28067 28500 28076
rect 28448 28033 28457 28067
rect 28457 28033 28491 28067
rect 28491 28033 28500 28067
rect 28448 28024 28500 28033
rect 29644 28067 29696 28076
rect 29644 28033 29653 28067
rect 29653 28033 29687 28067
rect 29687 28033 29696 28067
rect 29644 28024 29696 28033
rect 29920 28067 29972 28076
rect 29920 28033 29929 28067
rect 29929 28033 29963 28067
rect 29963 28033 29972 28067
rect 29920 28024 29972 28033
rect 30196 28024 30248 28076
rect 28540 27956 28592 28008
rect 23112 27820 23164 27872
rect 26240 27820 26292 27872
rect 27068 27820 27120 27872
rect 30012 27956 30064 28008
rect 30380 27999 30432 28008
rect 30380 27965 30389 27999
rect 30389 27965 30423 27999
rect 30423 27965 30432 27999
rect 30380 27956 30432 27965
rect 30564 28067 30616 28076
rect 30564 28033 30573 28067
rect 30573 28033 30607 28067
rect 30607 28033 30616 28067
rect 30564 28024 30616 28033
rect 31392 28092 31444 28144
rect 31852 28092 31904 28144
rect 33324 28092 33376 28144
rect 32312 28024 32364 28076
rect 32404 28067 32456 28076
rect 32404 28033 32413 28067
rect 32413 28033 32447 28067
rect 32447 28033 32456 28067
rect 32404 28024 32456 28033
rect 32680 28067 32732 28076
rect 32680 28033 32689 28067
rect 32689 28033 32723 28067
rect 32723 28033 32732 28067
rect 32680 28024 32732 28033
rect 29000 27888 29052 27940
rect 29736 27888 29788 27940
rect 30472 27888 30524 27940
rect 27344 27863 27396 27872
rect 27344 27829 27353 27863
rect 27353 27829 27387 27863
rect 27387 27829 27396 27863
rect 27344 27820 27396 27829
rect 29092 27863 29144 27872
rect 29092 27829 29101 27863
rect 29101 27829 29135 27863
rect 29135 27829 29144 27863
rect 29092 27820 29144 27829
rect 29368 27820 29420 27872
rect 31852 27820 31904 27872
rect 32956 27863 33008 27872
rect 32956 27829 32965 27863
rect 32965 27829 32999 27863
rect 32999 27829 33008 27863
rect 32956 27820 33008 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2136 27616 2188 27668
rect 4988 27616 5040 27668
rect 5264 27616 5316 27668
rect 3148 27548 3200 27600
rect 7472 27616 7524 27668
rect 7748 27616 7800 27668
rect 10048 27616 10100 27668
rect 10232 27616 10284 27668
rect 11060 27616 11112 27668
rect 4528 27523 4580 27532
rect 4528 27489 4537 27523
rect 4537 27489 4571 27523
rect 4571 27489 4580 27523
rect 4528 27480 4580 27489
rect 5356 27480 5408 27532
rect 2412 27455 2464 27464
rect 2412 27421 2421 27455
rect 2421 27421 2455 27455
rect 2455 27421 2464 27455
rect 2412 27412 2464 27421
rect 4068 27412 4120 27464
rect 4620 27412 4672 27464
rect 6000 27412 6052 27464
rect 7380 27480 7432 27532
rect 6460 27412 6512 27464
rect 9036 27548 9088 27600
rect 15200 27616 15252 27668
rect 9220 27480 9272 27532
rect 12348 27480 12400 27532
rect 12716 27480 12768 27532
rect 14280 27548 14332 27600
rect 16948 27548 17000 27600
rect 17500 27548 17552 27600
rect 20720 27548 20772 27600
rect 22192 27616 22244 27668
rect 23296 27616 23348 27668
rect 25872 27616 25924 27668
rect 26700 27616 26752 27668
rect 27252 27616 27304 27668
rect 26332 27548 26384 27600
rect 29000 27616 29052 27668
rect 28816 27548 28868 27600
rect 30196 27616 30248 27668
rect 31024 27616 31076 27668
rect 31668 27659 31720 27668
rect 31668 27625 31677 27659
rect 31677 27625 31711 27659
rect 31711 27625 31720 27659
rect 31668 27616 31720 27625
rect 29184 27548 29236 27600
rect 15384 27480 15436 27532
rect 18972 27480 19024 27532
rect 21180 27480 21232 27532
rect 23388 27480 23440 27532
rect 25136 27523 25188 27532
rect 25136 27489 25145 27523
rect 25145 27489 25179 27523
rect 25179 27489 25188 27523
rect 25136 27480 25188 27489
rect 26240 27523 26292 27532
rect 26240 27489 26249 27523
rect 26249 27489 26283 27523
rect 26283 27489 26292 27523
rect 26240 27480 26292 27489
rect 26608 27480 26660 27532
rect 27344 27480 27396 27532
rect 29828 27523 29880 27532
rect 29828 27489 29837 27523
rect 29837 27489 29871 27523
rect 29871 27489 29880 27523
rect 29828 27480 29880 27489
rect 1400 27344 1452 27396
rect 4804 27387 4856 27396
rect 4804 27353 4813 27387
rect 4813 27353 4847 27387
rect 4847 27353 4856 27387
rect 4804 27344 4856 27353
rect 5356 27319 5408 27328
rect 5356 27285 5365 27319
rect 5365 27285 5399 27319
rect 5399 27285 5408 27319
rect 5356 27276 5408 27285
rect 5724 27319 5776 27328
rect 5724 27285 5733 27319
rect 5733 27285 5767 27319
rect 5767 27285 5776 27319
rect 5724 27276 5776 27285
rect 5908 27319 5960 27328
rect 5908 27285 5917 27319
rect 5917 27285 5951 27319
rect 5951 27285 5960 27319
rect 5908 27276 5960 27285
rect 6092 27344 6144 27396
rect 9128 27455 9180 27464
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 9496 27455 9548 27464
rect 9496 27421 9505 27455
rect 9505 27421 9539 27455
rect 9539 27421 9548 27455
rect 9496 27412 9548 27421
rect 9588 27412 9640 27464
rect 10416 27455 10468 27464
rect 10416 27421 10425 27455
rect 10425 27421 10459 27455
rect 10459 27421 10468 27455
rect 10416 27412 10468 27421
rect 10784 27412 10836 27464
rect 8024 27387 8076 27396
rect 8024 27353 8033 27387
rect 8033 27353 8067 27387
rect 8067 27353 8076 27387
rect 8024 27344 8076 27353
rect 8116 27344 8168 27396
rect 11336 27344 11388 27396
rect 11796 27455 11848 27464
rect 11796 27421 11806 27455
rect 11806 27421 11840 27455
rect 11840 27421 11848 27455
rect 11796 27412 11848 27421
rect 12164 27455 12216 27464
rect 12164 27421 12173 27455
rect 12173 27421 12207 27455
rect 12207 27421 12216 27455
rect 12164 27412 12216 27421
rect 12440 27455 12492 27464
rect 12440 27421 12449 27455
rect 12449 27421 12483 27455
rect 12483 27421 12492 27455
rect 12440 27412 12492 27421
rect 12900 27412 12952 27464
rect 13452 27455 13504 27464
rect 12256 27344 12308 27396
rect 12532 27344 12584 27396
rect 13452 27421 13461 27455
rect 13461 27421 13495 27455
rect 13495 27421 13504 27455
rect 13452 27412 13504 27421
rect 13544 27455 13596 27464
rect 13544 27421 13553 27455
rect 13553 27421 13587 27455
rect 13587 27421 13596 27455
rect 13544 27412 13596 27421
rect 14096 27412 14148 27464
rect 16304 27412 16356 27464
rect 17132 27412 17184 27464
rect 15476 27344 15528 27396
rect 15568 27387 15620 27396
rect 15568 27353 15577 27387
rect 15577 27353 15611 27387
rect 15611 27353 15620 27387
rect 15568 27344 15620 27353
rect 17040 27344 17092 27396
rect 18604 27387 18656 27396
rect 18604 27353 18613 27387
rect 18613 27353 18647 27387
rect 18647 27353 18656 27387
rect 18604 27344 18656 27353
rect 18696 27344 18748 27396
rect 19432 27412 19484 27464
rect 19616 27412 19668 27464
rect 19984 27412 20036 27464
rect 21272 27455 21324 27464
rect 21272 27421 21281 27455
rect 21281 27421 21315 27455
rect 21315 27421 21324 27455
rect 21272 27412 21324 27421
rect 23572 27455 23624 27464
rect 23572 27421 23581 27455
rect 23581 27421 23615 27455
rect 23615 27421 23624 27455
rect 23572 27412 23624 27421
rect 23756 27455 23808 27464
rect 23756 27421 23765 27455
rect 23765 27421 23799 27455
rect 23799 27421 23808 27455
rect 23756 27412 23808 27421
rect 23940 27455 23992 27464
rect 23940 27421 23949 27455
rect 23949 27421 23983 27455
rect 23983 27421 23992 27455
rect 23940 27412 23992 27421
rect 25872 27412 25924 27464
rect 21548 27387 21600 27396
rect 21548 27353 21557 27387
rect 21557 27353 21591 27387
rect 21591 27353 21600 27387
rect 21548 27344 21600 27353
rect 23112 27344 23164 27396
rect 27068 27412 27120 27464
rect 27528 27412 27580 27464
rect 31116 27548 31168 27600
rect 31208 27548 31260 27600
rect 31484 27548 31536 27600
rect 34612 27548 34664 27600
rect 30104 27480 30156 27532
rect 30656 27480 30708 27532
rect 30932 27480 30984 27532
rect 31024 27455 31076 27464
rect 31024 27421 31033 27455
rect 31033 27421 31067 27455
rect 31067 27421 31076 27455
rect 31024 27412 31076 27421
rect 10784 27276 10836 27328
rect 10968 27319 11020 27328
rect 10968 27285 10977 27319
rect 10977 27285 11011 27319
rect 11011 27285 11020 27319
rect 10968 27276 11020 27285
rect 11244 27276 11296 27328
rect 11704 27276 11756 27328
rect 16304 27276 16356 27328
rect 18328 27276 18380 27328
rect 18512 27276 18564 27328
rect 20904 27276 20956 27328
rect 21916 27276 21968 27328
rect 22836 27276 22888 27328
rect 26056 27276 26108 27328
rect 26608 27319 26660 27328
rect 26608 27285 26617 27319
rect 26617 27285 26651 27319
rect 26651 27285 26660 27319
rect 26608 27276 26660 27285
rect 27252 27344 27304 27396
rect 29092 27344 29144 27396
rect 31852 27455 31904 27464
rect 31852 27421 31861 27455
rect 31861 27421 31895 27455
rect 31895 27421 31904 27455
rect 31852 27412 31904 27421
rect 26884 27276 26936 27328
rect 27804 27276 27856 27328
rect 30104 27276 30156 27328
rect 30748 27319 30800 27328
rect 30748 27285 30757 27319
rect 30757 27285 30791 27319
rect 30791 27285 30800 27319
rect 30748 27276 30800 27285
rect 30932 27319 30984 27328
rect 30932 27285 30941 27319
rect 30941 27285 30975 27319
rect 30975 27285 30984 27319
rect 30932 27276 30984 27285
rect 33508 27276 33560 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 2872 27072 2924 27124
rect 3424 27072 3476 27124
rect 4620 27072 4672 27124
rect 7932 27072 7984 27124
rect 8116 27072 8168 27124
rect 9496 27072 9548 27124
rect 10876 27072 10928 27124
rect 2780 27004 2832 27056
rect 5356 27004 5408 27056
rect 6460 27004 6512 27056
rect 12992 27072 13044 27124
rect 13360 27072 13412 27124
rect 14740 27072 14792 27124
rect 12532 27004 12584 27056
rect 12716 27004 12768 27056
rect 5724 26936 5776 26988
rect 7196 26936 7248 26988
rect 7288 26979 7340 26988
rect 7288 26945 7297 26979
rect 7297 26945 7331 26979
rect 7331 26945 7340 26979
rect 7288 26936 7340 26945
rect 7656 26936 7708 26988
rect 9128 26936 9180 26988
rect 3700 26868 3752 26920
rect 4528 26868 4580 26920
rect 4988 26911 5040 26920
rect 4988 26877 4997 26911
rect 4997 26877 5031 26911
rect 5031 26877 5040 26911
rect 4988 26868 5040 26877
rect 4068 26800 4120 26852
rect 7472 26868 7524 26920
rect 5264 26800 5316 26852
rect 9588 26800 9640 26852
rect 11336 26979 11388 26988
rect 11336 26945 11345 26979
rect 11345 26945 11379 26979
rect 11379 26945 11388 26979
rect 11336 26936 11388 26945
rect 12164 26979 12216 26988
rect 12164 26945 12173 26979
rect 12173 26945 12207 26979
rect 12207 26945 12216 26979
rect 12164 26936 12216 26945
rect 12900 26936 12952 26988
rect 13452 26936 13504 26988
rect 14188 26936 14240 26988
rect 16488 27072 16540 27124
rect 18604 27072 18656 27124
rect 21548 27072 21600 27124
rect 10968 26800 11020 26852
rect 11152 26843 11204 26852
rect 11152 26809 11161 26843
rect 11161 26809 11195 26843
rect 11195 26809 11204 26843
rect 11152 26800 11204 26809
rect 14372 26911 14424 26920
rect 14372 26877 14381 26911
rect 14381 26877 14415 26911
rect 14415 26877 14424 26911
rect 14372 26868 14424 26877
rect 16396 26936 16448 26988
rect 16580 26936 16632 26988
rect 16028 26868 16080 26920
rect 17224 26979 17276 26988
rect 17224 26945 17233 26979
rect 17233 26945 17267 26979
rect 17267 26945 17276 26979
rect 17224 26936 17276 26945
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 17408 26936 17460 26945
rect 17500 26936 17552 26988
rect 17960 26936 18012 26988
rect 18512 27004 18564 27056
rect 18972 27004 19024 27056
rect 23112 27072 23164 27124
rect 22560 27004 22612 27056
rect 18144 26936 18196 26988
rect 17316 26868 17368 26920
rect 14740 26800 14792 26852
rect 5448 26732 5500 26784
rect 7288 26732 7340 26784
rect 9036 26732 9088 26784
rect 13360 26732 13412 26784
rect 13728 26732 13780 26784
rect 16948 26732 17000 26784
rect 18604 26936 18656 26988
rect 18696 26979 18748 26988
rect 18696 26945 18705 26979
rect 18705 26945 18739 26979
rect 18739 26945 18748 26979
rect 18696 26936 18748 26945
rect 20720 26936 20772 26988
rect 20904 26979 20956 26988
rect 20904 26945 20913 26979
rect 20913 26945 20947 26979
rect 20947 26945 20956 26979
rect 20904 26936 20956 26945
rect 21088 26936 21140 26988
rect 24952 27072 25004 27124
rect 25044 27072 25096 27124
rect 31484 27072 31536 27124
rect 25136 27004 25188 27056
rect 21456 26868 21508 26920
rect 21824 26868 21876 26920
rect 20352 26800 20404 26852
rect 22008 26800 22060 26852
rect 19524 26732 19576 26784
rect 19984 26732 20036 26784
rect 24768 26936 24820 26988
rect 26056 26979 26108 26988
rect 26056 26945 26065 26979
rect 26065 26945 26099 26979
rect 26099 26945 26108 26979
rect 26056 26936 26108 26945
rect 26240 26979 26292 26988
rect 26240 26945 26249 26979
rect 26249 26945 26283 26979
rect 26283 26945 26292 26979
rect 26240 26936 26292 26945
rect 26424 26936 26476 26988
rect 27160 27004 27212 27056
rect 32680 27004 32732 27056
rect 34428 27004 34480 27056
rect 27436 26979 27488 26988
rect 27436 26945 27445 26979
rect 27445 26945 27479 26979
rect 27479 26945 27488 26979
rect 27436 26936 27488 26945
rect 27528 26979 27580 26988
rect 27528 26945 27537 26979
rect 27537 26945 27571 26979
rect 27571 26945 27580 26979
rect 27528 26936 27580 26945
rect 31668 26936 31720 26988
rect 33140 26936 33192 26988
rect 33968 26936 34020 26988
rect 22192 26911 22244 26920
rect 22192 26877 22201 26911
rect 22201 26877 22235 26911
rect 22235 26877 22244 26911
rect 22192 26868 22244 26877
rect 22560 26868 22612 26920
rect 22928 26868 22980 26920
rect 23940 26868 23992 26920
rect 27620 26868 27672 26920
rect 24768 26800 24820 26852
rect 31208 26868 31260 26920
rect 31576 26868 31628 26920
rect 34704 26936 34756 26988
rect 23204 26732 23256 26784
rect 23480 26732 23532 26784
rect 24492 26775 24544 26784
rect 24492 26741 24501 26775
rect 24501 26741 24535 26775
rect 24535 26741 24544 26775
rect 24492 26732 24544 26741
rect 25964 26732 26016 26784
rect 26792 26732 26844 26784
rect 27160 26732 27212 26784
rect 28448 26732 28500 26784
rect 32036 26800 32088 26852
rect 34612 26800 34664 26852
rect 32496 26732 32548 26784
rect 35348 26732 35400 26784
rect 35440 26732 35492 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3700 26528 3752 26580
rect 5356 26528 5408 26580
rect 6000 26528 6052 26580
rect 6460 26528 6512 26580
rect 7288 26528 7340 26580
rect 7472 26528 7524 26580
rect 7656 26528 7708 26580
rect 11336 26528 11388 26580
rect 11520 26571 11572 26580
rect 11520 26537 11529 26571
rect 11529 26537 11563 26571
rect 11563 26537 11572 26571
rect 11520 26528 11572 26537
rect 12900 26528 12952 26580
rect 16948 26528 17000 26580
rect 18144 26571 18196 26580
rect 18144 26537 18153 26571
rect 18153 26537 18187 26571
rect 18187 26537 18196 26571
rect 18144 26528 18196 26537
rect 21088 26528 21140 26580
rect 22376 26528 22428 26580
rect 22928 26528 22980 26580
rect 24952 26528 25004 26580
rect 25872 26528 25924 26580
rect 4436 26460 4488 26512
rect 4804 26460 4856 26512
rect 8392 26460 8444 26512
rect 2872 26392 2924 26444
rect 2964 26392 3016 26444
rect 3884 26392 3936 26444
rect 4068 26392 4120 26444
rect 4344 26435 4396 26444
rect 4344 26401 4353 26435
rect 4353 26401 4387 26435
rect 4387 26401 4396 26435
rect 4344 26392 4396 26401
rect 5724 26392 5776 26444
rect 2780 26324 2832 26376
rect 4620 26324 4672 26376
rect 4988 26324 5040 26376
rect 7196 26392 7248 26444
rect 6092 26256 6144 26308
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 6552 26256 6604 26308
rect 9036 26392 9088 26444
rect 10324 26392 10376 26444
rect 9588 26324 9640 26376
rect 11336 26324 11388 26376
rect 11980 26392 12032 26444
rect 8116 26256 8168 26308
rect 2688 26188 2740 26240
rect 4712 26188 4764 26240
rect 5356 26188 5408 26240
rect 12164 26256 12216 26308
rect 13636 26460 13688 26512
rect 15200 26460 15252 26512
rect 17040 26460 17092 26512
rect 17224 26460 17276 26512
rect 20260 26503 20312 26512
rect 20260 26469 20269 26503
rect 20269 26469 20303 26503
rect 20303 26469 20312 26503
rect 20260 26460 20312 26469
rect 13360 26435 13412 26444
rect 13360 26401 13369 26435
rect 13369 26401 13403 26435
rect 13403 26401 13412 26435
rect 13360 26392 13412 26401
rect 12532 26324 12584 26376
rect 12808 26324 12860 26376
rect 12900 26299 12952 26308
rect 12900 26265 12909 26299
rect 12909 26265 12943 26299
rect 12943 26265 12952 26299
rect 12900 26256 12952 26265
rect 12992 26299 13044 26308
rect 12992 26265 13001 26299
rect 13001 26265 13035 26299
rect 13035 26265 13044 26299
rect 12992 26256 13044 26265
rect 13728 26367 13780 26376
rect 13728 26333 13737 26367
rect 13737 26333 13771 26367
rect 13771 26333 13780 26367
rect 13728 26324 13780 26333
rect 18144 26392 18196 26444
rect 18512 26392 18564 26444
rect 23296 26460 23348 26512
rect 23388 26460 23440 26512
rect 25596 26460 25648 26512
rect 26700 26528 26752 26580
rect 28816 26528 28868 26580
rect 22100 26392 22152 26444
rect 25044 26392 25096 26444
rect 13820 26256 13872 26308
rect 14096 26256 14148 26308
rect 9496 26188 9548 26240
rect 10600 26188 10652 26240
rect 10692 26188 10744 26240
rect 10968 26188 11020 26240
rect 11244 26188 11296 26240
rect 11336 26188 11388 26240
rect 11796 26188 11848 26240
rect 12716 26188 12768 26240
rect 13452 26188 13504 26240
rect 15844 26367 15896 26376
rect 15844 26333 15853 26367
rect 15853 26333 15887 26367
rect 15887 26333 15896 26367
rect 15844 26324 15896 26333
rect 16028 26367 16080 26376
rect 16028 26333 16037 26367
rect 16037 26333 16071 26367
rect 16071 26333 16080 26367
rect 16028 26324 16080 26333
rect 16948 26367 17000 26376
rect 16948 26333 16957 26367
rect 16957 26333 16991 26367
rect 16991 26333 17000 26367
rect 16948 26324 17000 26333
rect 18604 26324 18656 26376
rect 20352 26367 20404 26376
rect 20352 26333 20361 26367
rect 20361 26333 20395 26367
rect 20395 26333 20404 26367
rect 20352 26324 20404 26333
rect 15844 26188 15896 26240
rect 16028 26231 16080 26240
rect 16028 26197 16037 26231
rect 16037 26197 16071 26231
rect 16071 26197 16080 26231
rect 16028 26188 16080 26197
rect 16396 26188 16448 26240
rect 17316 26299 17368 26308
rect 17316 26265 17325 26299
rect 17325 26265 17359 26299
rect 17359 26265 17368 26299
rect 17316 26256 17368 26265
rect 17500 26299 17552 26308
rect 17500 26265 17509 26299
rect 17509 26265 17543 26299
rect 17543 26265 17552 26299
rect 17500 26256 17552 26265
rect 19248 26256 19300 26308
rect 19984 26299 20036 26308
rect 19984 26265 19993 26299
rect 19993 26265 20027 26299
rect 20027 26265 20036 26299
rect 19984 26256 20036 26265
rect 20260 26256 20312 26308
rect 22928 26324 22980 26376
rect 20720 26256 20772 26308
rect 21364 26256 21416 26308
rect 16764 26188 16816 26240
rect 19432 26188 19484 26240
rect 19616 26188 19668 26240
rect 21824 26256 21876 26308
rect 21916 26299 21968 26308
rect 21916 26265 21925 26299
rect 21925 26265 21959 26299
rect 21959 26265 21968 26299
rect 21916 26256 21968 26265
rect 22008 26256 22060 26308
rect 22744 26256 22796 26308
rect 23112 26324 23164 26376
rect 25412 26367 25464 26376
rect 25412 26333 25421 26367
rect 25421 26333 25455 26367
rect 25455 26333 25464 26367
rect 25412 26324 25464 26333
rect 25780 26392 25832 26444
rect 25872 26367 25924 26376
rect 25872 26333 25881 26367
rect 25881 26333 25915 26367
rect 25915 26333 25924 26367
rect 25872 26324 25924 26333
rect 26608 26392 26660 26444
rect 26976 26392 27028 26444
rect 26240 26367 26292 26376
rect 26240 26333 26249 26367
rect 26249 26333 26283 26367
rect 26283 26333 26292 26367
rect 26240 26324 26292 26333
rect 26700 26367 26752 26376
rect 26700 26333 26709 26367
rect 26709 26333 26743 26367
rect 26743 26333 26752 26367
rect 26700 26324 26752 26333
rect 21640 26188 21692 26240
rect 23664 26188 23716 26240
rect 25780 26299 25832 26308
rect 25780 26265 25789 26299
rect 25789 26265 25823 26299
rect 25823 26265 25832 26299
rect 25780 26256 25832 26265
rect 26976 26256 27028 26308
rect 27436 26367 27488 26376
rect 27436 26333 27445 26367
rect 27445 26333 27479 26367
rect 27479 26333 27488 26367
rect 27436 26324 27488 26333
rect 27712 26367 27764 26376
rect 27712 26333 27721 26367
rect 27721 26333 27755 26367
rect 27755 26333 27764 26367
rect 27712 26324 27764 26333
rect 27896 26367 27948 26376
rect 27896 26333 27903 26367
rect 27903 26333 27948 26367
rect 27896 26324 27948 26333
rect 27988 26367 28040 26376
rect 27988 26333 27997 26367
rect 27997 26333 28031 26367
rect 28031 26333 28040 26367
rect 27988 26324 28040 26333
rect 28448 26324 28500 26376
rect 29460 26324 29512 26376
rect 29644 26367 29696 26376
rect 29644 26333 29653 26367
rect 29653 26333 29687 26367
rect 29687 26333 29696 26367
rect 29644 26324 29696 26333
rect 31576 26528 31628 26580
rect 31760 26528 31812 26580
rect 32128 26528 32180 26580
rect 30380 26460 30432 26512
rect 30932 26460 30984 26512
rect 32128 26392 32180 26444
rect 32404 26392 32456 26444
rect 32680 26392 32732 26444
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 29920 26324 29972 26333
rect 27620 26256 27672 26308
rect 26424 26188 26476 26240
rect 26792 26188 26844 26240
rect 27252 26188 27304 26240
rect 31852 26324 31904 26376
rect 33968 26324 34020 26376
rect 32036 26299 32088 26308
rect 32036 26265 32045 26299
rect 32045 26265 32079 26299
rect 32079 26265 32088 26299
rect 32036 26256 32088 26265
rect 31944 26188 31996 26240
rect 33140 26256 33192 26308
rect 33324 26256 33376 26308
rect 34152 26367 34204 26376
rect 34152 26333 34161 26367
rect 34161 26333 34195 26367
rect 34195 26333 34204 26367
rect 34152 26324 34204 26333
rect 32404 26231 32456 26240
rect 32404 26197 32413 26231
rect 32413 26197 32447 26231
rect 32447 26197 32456 26231
rect 32404 26188 32456 26197
rect 33784 26188 33836 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 2136 26027 2188 26036
rect 2136 25993 2145 26027
rect 2145 25993 2179 26027
rect 2179 25993 2188 26027
rect 2136 25984 2188 25993
rect 3056 25984 3108 26036
rect 4344 25984 4396 26036
rect 4436 26027 4488 26036
rect 4436 25993 4445 26027
rect 4445 25993 4479 26027
rect 4479 25993 4488 26027
rect 4436 25984 4488 25993
rect 4712 25984 4764 26036
rect 5264 25984 5316 26036
rect 6092 26027 6144 26036
rect 6092 25993 6101 26027
rect 6101 25993 6135 26027
rect 6135 25993 6144 26027
rect 6092 25984 6144 25993
rect 2320 25780 2372 25832
rect 4620 25916 4672 25968
rect 7380 25916 7432 25968
rect 7840 25916 7892 25968
rect 3976 25848 4028 25900
rect 4344 25848 4396 25900
rect 1676 25644 1728 25696
rect 4712 25780 4764 25832
rect 3884 25712 3936 25764
rect 4988 25780 5040 25832
rect 5540 25780 5592 25832
rect 6552 25848 6604 25900
rect 7196 25848 7248 25900
rect 8484 25848 8536 25900
rect 6736 25780 6788 25832
rect 2872 25644 2924 25696
rect 3424 25644 3476 25696
rect 5264 25687 5316 25696
rect 5264 25653 5273 25687
rect 5273 25653 5307 25687
rect 5307 25653 5316 25687
rect 5264 25644 5316 25653
rect 5356 25644 5408 25696
rect 7840 25687 7892 25696
rect 7840 25653 7849 25687
rect 7849 25653 7883 25687
rect 7883 25653 7892 25687
rect 7840 25644 7892 25653
rect 9404 25916 9456 25968
rect 9496 25891 9548 25900
rect 9496 25857 9505 25891
rect 9505 25857 9539 25891
rect 9539 25857 9548 25891
rect 9496 25848 9548 25857
rect 9772 25959 9824 25968
rect 9772 25925 9781 25959
rect 9781 25925 9815 25959
rect 9815 25925 9824 25959
rect 9772 25916 9824 25925
rect 10140 25916 10192 25968
rect 10968 25959 11020 25968
rect 10968 25925 10977 25959
rect 10977 25925 11011 25959
rect 11011 25925 11020 25959
rect 10968 25916 11020 25925
rect 11244 25984 11296 26036
rect 11336 25916 11388 25968
rect 11520 25916 11572 25968
rect 10600 25891 10652 25900
rect 10600 25857 10609 25891
rect 10609 25857 10643 25891
rect 10643 25857 10652 25891
rect 10600 25848 10652 25857
rect 10784 25848 10836 25900
rect 11060 25891 11112 25900
rect 11060 25857 11069 25891
rect 11069 25857 11103 25891
rect 11103 25857 11112 25891
rect 11060 25848 11112 25857
rect 12624 25984 12676 26036
rect 13820 25984 13872 26036
rect 15108 25984 15160 26036
rect 19432 25984 19484 26036
rect 20444 25984 20496 26036
rect 16672 25916 16724 25968
rect 19984 25916 20036 25968
rect 20168 25916 20220 25968
rect 9588 25712 9640 25764
rect 11980 25823 12032 25832
rect 11980 25789 11989 25823
rect 11989 25789 12023 25823
rect 12023 25789 12032 25823
rect 11980 25780 12032 25789
rect 12624 25891 12676 25900
rect 12624 25857 12633 25891
rect 12633 25857 12667 25891
rect 12667 25857 12676 25891
rect 12624 25848 12676 25857
rect 12808 25891 12860 25900
rect 12808 25857 12822 25891
rect 12822 25857 12856 25891
rect 12856 25857 12860 25891
rect 12808 25848 12860 25857
rect 14464 25891 14516 25900
rect 14464 25857 14473 25891
rect 14473 25857 14507 25891
rect 14507 25857 14516 25891
rect 14464 25848 14516 25857
rect 14832 25891 14884 25900
rect 14832 25857 14840 25891
rect 14840 25857 14874 25891
rect 14874 25857 14884 25891
rect 14832 25848 14884 25857
rect 12532 25780 12584 25832
rect 15016 25891 15068 25900
rect 15016 25857 15025 25891
rect 15025 25857 15059 25891
rect 15059 25857 15068 25891
rect 15016 25848 15068 25857
rect 15200 25891 15252 25900
rect 15200 25857 15209 25891
rect 15209 25857 15243 25891
rect 15243 25857 15252 25891
rect 15200 25848 15252 25857
rect 15936 25891 15988 25900
rect 15936 25857 15945 25891
rect 15945 25857 15979 25891
rect 15979 25857 15988 25891
rect 15936 25848 15988 25857
rect 15108 25780 15160 25832
rect 15844 25823 15896 25832
rect 15844 25789 15853 25823
rect 15853 25789 15887 25823
rect 15887 25789 15896 25823
rect 15844 25780 15896 25789
rect 17868 25823 17920 25832
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 18144 25891 18196 25900
rect 18144 25857 18153 25891
rect 18153 25857 18187 25891
rect 18187 25857 18196 25891
rect 18144 25848 18196 25857
rect 18420 25891 18472 25900
rect 18420 25857 18429 25891
rect 18429 25857 18463 25891
rect 18463 25857 18472 25891
rect 18420 25848 18472 25857
rect 16488 25712 16540 25764
rect 18880 25848 18932 25900
rect 21364 25916 21416 25968
rect 18788 25780 18840 25832
rect 19524 25823 19576 25832
rect 19524 25789 19533 25823
rect 19533 25789 19567 25823
rect 19567 25789 19576 25823
rect 19524 25780 19576 25789
rect 19984 25780 20036 25832
rect 20352 25780 20404 25832
rect 21180 25823 21232 25832
rect 21180 25789 21189 25823
rect 21189 25789 21223 25823
rect 21223 25789 21232 25823
rect 21180 25780 21232 25789
rect 22008 25891 22060 25900
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 22836 25916 22888 25968
rect 29644 25984 29696 26036
rect 30564 25984 30616 26036
rect 32128 26027 32180 26036
rect 32128 25993 32137 26027
rect 32137 25993 32171 26027
rect 32171 25993 32180 26027
rect 32128 25984 32180 25993
rect 32312 25984 32364 26036
rect 21548 25780 21600 25832
rect 20812 25712 20864 25764
rect 9312 25644 9364 25696
rect 9404 25687 9456 25696
rect 9404 25653 9413 25687
rect 9413 25653 9447 25687
rect 9447 25653 9456 25687
rect 9404 25644 9456 25653
rect 9496 25644 9548 25696
rect 9772 25644 9824 25696
rect 10692 25644 10744 25696
rect 10968 25644 11020 25696
rect 12440 25644 12492 25696
rect 12992 25687 13044 25696
rect 12992 25653 13001 25687
rect 13001 25653 13035 25687
rect 13035 25653 13044 25687
rect 12992 25644 13044 25653
rect 14096 25687 14148 25696
rect 14096 25653 14105 25687
rect 14105 25653 14139 25687
rect 14139 25653 14148 25687
rect 14096 25644 14148 25653
rect 17868 25644 17920 25696
rect 18880 25644 18932 25696
rect 19616 25644 19668 25696
rect 19984 25644 20036 25696
rect 20352 25644 20404 25696
rect 21732 25644 21784 25696
rect 22560 25891 22612 25900
rect 22560 25857 22569 25891
rect 22569 25857 22603 25891
rect 22603 25857 22612 25891
rect 22560 25848 22612 25857
rect 23020 25780 23072 25832
rect 23572 25891 23624 25900
rect 23572 25857 23581 25891
rect 23581 25857 23615 25891
rect 23615 25857 23624 25891
rect 23572 25848 23624 25857
rect 23664 25891 23716 25900
rect 23664 25857 23674 25891
rect 23674 25857 23708 25891
rect 23708 25857 23716 25891
rect 23664 25848 23716 25857
rect 23848 25891 23900 25900
rect 23848 25857 23857 25891
rect 23857 25857 23891 25891
rect 23891 25857 23900 25891
rect 23848 25848 23900 25857
rect 23940 25891 23992 25900
rect 23940 25857 23949 25891
rect 23949 25857 23983 25891
rect 23983 25857 23992 25891
rect 23940 25848 23992 25857
rect 24952 25916 25004 25968
rect 25228 25916 25280 25968
rect 24216 25712 24268 25764
rect 24584 25891 24636 25900
rect 24584 25857 24593 25891
rect 24593 25857 24627 25891
rect 24627 25857 24636 25891
rect 24584 25848 24636 25857
rect 24860 25891 24912 25900
rect 24860 25857 24869 25891
rect 24869 25857 24903 25891
rect 24903 25857 24912 25891
rect 24860 25848 24912 25857
rect 25320 25891 25372 25900
rect 25320 25857 25329 25891
rect 25329 25857 25363 25891
rect 25363 25857 25372 25891
rect 25320 25848 25372 25857
rect 26056 25891 26108 25900
rect 26056 25857 26065 25891
rect 26065 25857 26099 25891
rect 26099 25857 26108 25891
rect 26056 25848 26108 25857
rect 26608 25848 26660 25900
rect 27620 25848 27672 25900
rect 28632 25780 28684 25832
rect 29184 25848 29236 25900
rect 30012 25916 30064 25968
rect 32588 25984 32640 26036
rect 29368 25780 29420 25832
rect 31024 25848 31076 25900
rect 32036 25848 32088 25900
rect 32588 25848 32640 25900
rect 32864 25916 32916 25968
rect 33508 25984 33560 26036
rect 34704 25984 34756 26036
rect 33324 25848 33376 25900
rect 34428 25916 34480 25968
rect 33968 25848 34020 25900
rect 34060 25891 34112 25900
rect 34060 25857 34069 25891
rect 34069 25857 34103 25891
rect 34103 25857 34112 25891
rect 34060 25848 34112 25857
rect 29736 25712 29788 25764
rect 33876 25780 33928 25832
rect 32128 25712 32180 25764
rect 32404 25712 32456 25764
rect 36084 25823 36136 25832
rect 36084 25789 36093 25823
rect 36093 25789 36127 25823
rect 36127 25789 36136 25823
rect 36084 25780 36136 25789
rect 23480 25644 23532 25696
rect 23940 25644 23992 25696
rect 29368 25644 29420 25696
rect 29920 25687 29972 25696
rect 29920 25653 29929 25687
rect 29929 25653 29963 25687
rect 29963 25653 29972 25687
rect 29920 25644 29972 25653
rect 30196 25644 30248 25696
rect 33508 25687 33560 25696
rect 33508 25653 33517 25687
rect 33517 25653 33551 25687
rect 33551 25653 33560 25687
rect 33508 25644 33560 25653
rect 35440 25644 35492 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3148 25483 3200 25492
rect 3148 25449 3157 25483
rect 3157 25449 3191 25483
rect 3191 25449 3200 25483
rect 3148 25440 3200 25449
rect 4620 25440 4672 25492
rect 4712 25440 4764 25492
rect 9404 25440 9456 25492
rect 9772 25483 9824 25492
rect 9772 25449 9781 25483
rect 9781 25449 9815 25483
rect 9815 25449 9824 25483
rect 9772 25440 9824 25449
rect 10140 25440 10192 25492
rect 10416 25440 10468 25492
rect 10968 25440 11020 25492
rect 18420 25440 18472 25492
rect 19800 25440 19852 25492
rect 7380 25372 7432 25424
rect 8208 25372 8260 25424
rect 8484 25415 8536 25424
rect 8484 25381 8493 25415
rect 8493 25381 8527 25415
rect 8527 25381 8536 25415
rect 8484 25372 8536 25381
rect 8852 25372 8904 25424
rect 9036 25372 9088 25424
rect 11152 25372 11204 25424
rect 11980 25372 12032 25424
rect 2872 25304 2924 25356
rect 5264 25347 5316 25356
rect 5264 25313 5273 25347
rect 5273 25313 5307 25347
rect 5307 25313 5316 25347
rect 5264 25304 5316 25313
rect 5540 25304 5592 25356
rect 6920 25304 6972 25356
rect 2780 25236 2832 25288
rect 3976 25236 4028 25288
rect 5908 25279 5960 25288
rect 5908 25245 5917 25279
rect 5917 25245 5951 25279
rect 5951 25245 5960 25279
rect 5908 25236 5960 25245
rect 1676 25211 1728 25220
rect 1676 25177 1685 25211
rect 1685 25177 1719 25211
rect 1719 25177 1728 25211
rect 1676 25168 1728 25177
rect 4068 25168 4120 25220
rect 6092 25168 6144 25220
rect 6828 25211 6880 25220
rect 6828 25177 6837 25211
rect 6837 25177 6871 25211
rect 6871 25177 6880 25211
rect 6828 25168 6880 25177
rect 6920 25211 6972 25220
rect 6920 25177 6929 25211
rect 6929 25177 6963 25211
rect 6963 25177 6972 25211
rect 6920 25168 6972 25177
rect 2320 25100 2372 25152
rect 3148 25100 3200 25152
rect 4620 25100 4672 25152
rect 5448 25100 5500 25152
rect 5724 25143 5776 25152
rect 5724 25109 5733 25143
rect 5733 25109 5767 25143
rect 5767 25109 5776 25143
rect 5724 25100 5776 25109
rect 7196 25279 7248 25288
rect 7196 25245 7205 25279
rect 7205 25245 7239 25279
rect 7239 25245 7248 25279
rect 7196 25236 7248 25245
rect 7380 25279 7432 25288
rect 7380 25245 7389 25279
rect 7389 25245 7423 25279
rect 7423 25245 7432 25279
rect 7380 25236 7432 25245
rect 7656 25236 7708 25288
rect 8024 25279 8076 25288
rect 8024 25245 8033 25279
rect 8033 25245 8067 25279
rect 8067 25245 8076 25279
rect 8024 25236 8076 25245
rect 8208 25279 8260 25288
rect 8208 25245 8217 25279
rect 8217 25245 8251 25279
rect 8251 25245 8260 25279
rect 8208 25236 8260 25245
rect 8484 25236 8536 25288
rect 9404 25279 9456 25288
rect 9404 25245 9413 25279
rect 9413 25245 9447 25279
rect 9447 25245 9456 25279
rect 9404 25236 9456 25245
rect 9588 25279 9640 25288
rect 9588 25245 9597 25279
rect 9597 25245 9631 25279
rect 9631 25245 9640 25279
rect 9588 25236 9640 25245
rect 9772 25236 9824 25288
rect 10048 25279 10100 25288
rect 10048 25245 10057 25279
rect 10057 25245 10091 25279
rect 10091 25245 10100 25279
rect 10048 25236 10100 25245
rect 10968 25236 11020 25288
rect 11612 25279 11664 25288
rect 11612 25245 11621 25279
rect 11621 25245 11655 25279
rect 11655 25245 11664 25279
rect 11612 25236 11664 25245
rect 11888 25304 11940 25356
rect 14464 25279 14516 25288
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 15844 25372 15896 25424
rect 15016 25304 15068 25356
rect 9036 25168 9088 25220
rect 10876 25168 10928 25220
rect 11336 25168 11388 25220
rect 12164 25168 12216 25220
rect 13084 25168 13136 25220
rect 13452 25168 13504 25220
rect 13820 25168 13872 25220
rect 14280 25168 14332 25220
rect 15108 25279 15160 25288
rect 15108 25245 15117 25279
rect 15117 25245 15151 25279
rect 15151 25245 15160 25279
rect 15108 25236 15160 25245
rect 15292 25236 15344 25288
rect 16304 25236 16356 25288
rect 16764 25279 16816 25288
rect 16764 25245 16773 25279
rect 16773 25245 16807 25279
rect 16807 25245 16816 25279
rect 16764 25236 16816 25245
rect 16948 25236 17000 25288
rect 18880 25372 18932 25424
rect 18972 25372 19024 25424
rect 21548 25440 21600 25492
rect 21824 25440 21876 25492
rect 22836 25440 22888 25492
rect 23296 25483 23348 25492
rect 23296 25449 23305 25483
rect 23305 25449 23339 25483
rect 23339 25449 23348 25483
rect 23296 25440 23348 25449
rect 24860 25483 24912 25492
rect 24860 25449 24869 25483
rect 24869 25449 24903 25483
rect 24903 25449 24912 25483
rect 24860 25440 24912 25449
rect 26424 25440 26476 25492
rect 33048 25440 33100 25492
rect 33324 25483 33376 25492
rect 33324 25449 33333 25483
rect 33333 25449 33367 25483
rect 33367 25449 33376 25483
rect 33324 25440 33376 25449
rect 33600 25440 33652 25492
rect 34428 25440 34480 25492
rect 20076 25372 20128 25424
rect 18880 25236 18932 25288
rect 21088 25304 21140 25356
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 20720 25236 20772 25245
rect 21640 25304 21692 25356
rect 23020 25372 23072 25424
rect 23664 25372 23716 25424
rect 25044 25415 25096 25424
rect 25044 25381 25053 25415
rect 25053 25381 25087 25415
rect 25087 25381 25096 25415
rect 25044 25372 25096 25381
rect 32128 25372 32180 25424
rect 23388 25304 23440 25356
rect 25320 25304 25372 25356
rect 32036 25304 32088 25356
rect 15936 25168 15988 25220
rect 16028 25211 16080 25220
rect 16028 25177 16037 25211
rect 16037 25177 16071 25211
rect 16071 25177 16080 25211
rect 16028 25168 16080 25177
rect 13728 25100 13780 25152
rect 14832 25100 14884 25152
rect 15844 25143 15896 25152
rect 15844 25109 15853 25143
rect 15853 25109 15887 25143
rect 15887 25109 15896 25143
rect 15844 25100 15896 25109
rect 16672 25168 16724 25220
rect 16764 25100 16816 25152
rect 18604 25211 18656 25220
rect 18604 25177 18613 25211
rect 18613 25177 18647 25211
rect 18647 25177 18656 25211
rect 18604 25168 18656 25177
rect 20168 25168 20220 25220
rect 21548 25279 21600 25288
rect 21548 25245 21557 25279
rect 21557 25245 21591 25279
rect 21591 25245 21600 25279
rect 21548 25236 21600 25245
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 22744 25236 22796 25288
rect 24216 25236 24268 25288
rect 25412 25236 25464 25288
rect 29000 25236 29052 25288
rect 20444 25100 20496 25152
rect 20536 25143 20588 25152
rect 20536 25109 20545 25143
rect 20545 25109 20579 25143
rect 20579 25109 20588 25143
rect 20536 25100 20588 25109
rect 22192 25168 22244 25220
rect 23020 25168 23072 25220
rect 26056 25168 26108 25220
rect 32128 25168 32180 25220
rect 32236 25245 32275 25266
rect 32275 25245 32288 25266
rect 32236 25214 32288 25245
rect 32496 25245 32548 25254
rect 32496 25211 32505 25245
rect 32505 25211 32539 25245
rect 32539 25211 32548 25245
rect 32496 25202 32548 25211
rect 32772 25236 32824 25288
rect 33692 25236 33744 25288
rect 33784 25236 33836 25288
rect 35440 25236 35492 25288
rect 22008 25100 22060 25152
rect 24860 25100 24912 25152
rect 28264 25100 28316 25152
rect 30012 25100 30064 25152
rect 36084 25168 36136 25220
rect 33968 25143 34020 25152
rect 33968 25109 33977 25143
rect 33977 25109 34011 25143
rect 34011 25109 34020 25143
rect 33968 25100 34020 25109
rect 34612 25100 34664 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 3976 24896 4028 24948
rect 2504 24828 2556 24880
rect 3148 24828 3200 24880
rect 5908 24896 5960 24948
rect 9220 24896 9272 24948
rect 11612 24896 11664 24948
rect 5724 24828 5776 24880
rect 6092 24828 6144 24880
rect 2872 24760 2924 24812
rect 6736 24760 6788 24812
rect 8024 24828 8076 24880
rect 7012 24803 7064 24812
rect 7012 24769 7021 24803
rect 7021 24769 7055 24803
rect 7055 24769 7064 24803
rect 7012 24760 7064 24769
rect 7288 24760 7340 24812
rect 3056 24692 3108 24744
rect 3976 24735 4028 24744
rect 3976 24701 3985 24735
rect 3985 24701 4019 24735
rect 4019 24701 4028 24735
rect 3976 24692 4028 24701
rect 8484 24692 8536 24744
rect 9036 24760 9088 24812
rect 9312 24828 9364 24880
rect 10600 24828 10652 24880
rect 12532 24896 12584 24948
rect 16304 24939 16356 24948
rect 16304 24905 16313 24939
rect 16313 24905 16347 24939
rect 16347 24905 16356 24939
rect 16304 24896 16356 24905
rect 21456 24896 21508 24948
rect 21824 24896 21876 24948
rect 22744 24939 22796 24948
rect 22744 24905 22753 24939
rect 22753 24905 22787 24939
rect 22787 24905 22796 24939
rect 22744 24896 22796 24905
rect 24032 24896 24084 24948
rect 25688 24896 25740 24948
rect 25872 24896 25924 24948
rect 27988 24896 28040 24948
rect 8852 24692 8904 24744
rect 9404 24803 9456 24812
rect 9404 24769 9413 24803
rect 9413 24769 9447 24803
rect 9447 24769 9456 24803
rect 9404 24760 9456 24769
rect 9588 24803 9640 24812
rect 9588 24769 9602 24803
rect 9602 24769 9636 24803
rect 9636 24769 9640 24803
rect 9588 24760 9640 24769
rect 11152 24803 11204 24812
rect 11152 24769 11161 24803
rect 11161 24769 11195 24803
rect 11195 24769 11204 24803
rect 11152 24760 11204 24769
rect 11336 24803 11388 24812
rect 11336 24769 11345 24803
rect 11345 24769 11379 24803
rect 11379 24769 11388 24803
rect 11336 24760 11388 24769
rect 9956 24692 10008 24744
rect 11796 24803 11848 24812
rect 11796 24769 11805 24803
rect 11805 24769 11839 24803
rect 11839 24769 11848 24803
rect 11796 24760 11848 24769
rect 12072 24760 12124 24812
rect 12256 24803 12308 24812
rect 12256 24769 12265 24803
rect 12265 24769 12299 24803
rect 12299 24769 12308 24803
rect 12256 24760 12308 24769
rect 13360 24828 13412 24880
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 12532 24760 12584 24769
rect 12808 24803 12860 24812
rect 12808 24769 12817 24803
rect 12817 24769 12851 24803
rect 12851 24769 12860 24803
rect 12808 24760 12860 24769
rect 12900 24760 12952 24812
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 14280 24760 14332 24812
rect 7012 24624 7064 24676
rect 8208 24624 8260 24676
rect 8576 24624 8628 24676
rect 10876 24624 10928 24676
rect 12440 24624 12492 24676
rect 13176 24692 13228 24744
rect 14832 24692 14884 24744
rect 16672 24760 16724 24812
rect 18512 24828 18564 24880
rect 18604 24828 18656 24880
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18788 24803 18840 24812
rect 18788 24769 18797 24803
rect 18797 24769 18831 24803
rect 18831 24769 18840 24803
rect 18788 24760 18840 24769
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 18972 24760 19024 24769
rect 20812 24828 20864 24880
rect 22008 24828 22060 24880
rect 19616 24803 19668 24812
rect 19616 24769 19625 24803
rect 19625 24769 19659 24803
rect 19659 24769 19668 24803
rect 19616 24760 19668 24769
rect 22928 24803 22980 24812
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 23388 24803 23440 24812
rect 23388 24769 23397 24803
rect 23397 24769 23431 24803
rect 23431 24769 23440 24803
rect 23388 24760 23440 24769
rect 23848 24760 23900 24812
rect 24952 24760 25004 24812
rect 17592 24692 17644 24744
rect 23756 24692 23808 24744
rect 24676 24692 24728 24744
rect 25872 24760 25924 24812
rect 25964 24803 26016 24812
rect 25964 24769 25973 24803
rect 25973 24769 26007 24803
rect 26007 24769 26016 24803
rect 25964 24760 26016 24769
rect 26056 24803 26108 24812
rect 26056 24769 26065 24803
rect 26065 24769 26099 24803
rect 26099 24769 26108 24803
rect 26056 24760 26108 24769
rect 26424 24760 26476 24812
rect 26608 24760 26660 24812
rect 27252 24803 27304 24812
rect 27252 24769 27261 24803
rect 27261 24769 27295 24803
rect 27295 24769 27304 24803
rect 27252 24760 27304 24769
rect 27528 24803 27580 24812
rect 27528 24769 27537 24803
rect 27537 24769 27571 24803
rect 27571 24769 27580 24803
rect 27528 24760 27580 24769
rect 27988 24760 28040 24812
rect 28264 24803 28316 24812
rect 28264 24769 28273 24803
rect 28273 24769 28307 24803
rect 28307 24769 28316 24803
rect 28264 24760 28316 24769
rect 29368 24896 29420 24948
rect 29552 24896 29604 24948
rect 32036 24896 32088 24948
rect 32588 24896 32640 24948
rect 35992 24896 36044 24948
rect 28908 24828 28960 24880
rect 29644 24828 29696 24880
rect 34152 24828 34204 24880
rect 13268 24624 13320 24676
rect 15200 24624 15252 24676
rect 17316 24624 17368 24676
rect 18420 24624 18472 24676
rect 18788 24624 18840 24676
rect 1676 24556 1728 24608
rect 5264 24556 5316 24608
rect 6460 24556 6512 24608
rect 9036 24556 9088 24608
rect 9680 24556 9732 24608
rect 9956 24556 10008 24608
rect 11152 24556 11204 24608
rect 11336 24599 11388 24608
rect 11336 24565 11345 24599
rect 11345 24565 11379 24599
rect 11379 24565 11388 24599
rect 11336 24556 11388 24565
rect 12348 24556 12400 24608
rect 16948 24599 17000 24608
rect 16948 24565 16957 24599
rect 16957 24565 16991 24599
rect 16991 24565 17000 24599
rect 16948 24556 17000 24565
rect 17040 24599 17092 24608
rect 17040 24565 17049 24599
rect 17049 24565 17083 24599
rect 17083 24565 17092 24599
rect 17040 24556 17092 24565
rect 17868 24599 17920 24608
rect 17868 24565 17877 24599
rect 17877 24565 17911 24599
rect 17911 24565 17920 24599
rect 17868 24556 17920 24565
rect 17960 24556 18012 24608
rect 20536 24624 20588 24676
rect 19432 24556 19484 24608
rect 20260 24556 20312 24608
rect 25044 24624 25096 24676
rect 26240 24624 26292 24676
rect 27160 24624 27212 24676
rect 23572 24556 23624 24608
rect 23756 24556 23808 24608
rect 24216 24556 24268 24608
rect 25136 24556 25188 24608
rect 27712 24667 27764 24676
rect 27712 24633 27721 24667
rect 27721 24633 27755 24667
rect 27755 24633 27764 24667
rect 27712 24624 27764 24633
rect 27896 24556 27948 24608
rect 28264 24556 28316 24608
rect 28816 24692 28868 24744
rect 29276 24735 29328 24744
rect 29276 24701 29285 24735
rect 29285 24701 29319 24735
rect 29319 24701 29328 24735
rect 29276 24692 29328 24701
rect 29644 24692 29696 24744
rect 29828 24692 29880 24744
rect 34336 24760 34388 24812
rect 35256 24760 35308 24812
rect 30656 24692 30708 24744
rect 31944 24692 31996 24744
rect 28724 24556 28776 24608
rect 29828 24556 29880 24608
rect 30288 24624 30340 24676
rect 35992 24803 36044 24812
rect 35992 24769 36001 24803
rect 36001 24769 36035 24803
rect 36035 24769 36044 24803
rect 35992 24760 36044 24769
rect 33692 24556 33744 24608
rect 34152 24556 34204 24608
rect 34336 24556 34388 24608
rect 35900 24556 35952 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3148 24395 3200 24404
rect 3148 24361 3157 24395
rect 3157 24361 3191 24395
rect 3191 24361 3200 24395
rect 3148 24352 3200 24361
rect 3608 24352 3660 24404
rect 3976 24352 4028 24404
rect 5816 24352 5868 24404
rect 6920 24352 6972 24404
rect 10968 24352 11020 24404
rect 6184 24284 6236 24336
rect 7288 24327 7340 24336
rect 7288 24293 7297 24327
rect 7297 24293 7331 24327
rect 7331 24293 7340 24327
rect 7288 24284 7340 24293
rect 1676 24259 1728 24268
rect 1676 24225 1685 24259
rect 1685 24225 1719 24259
rect 1719 24225 1728 24259
rect 1676 24216 1728 24225
rect 4804 24216 4856 24268
rect 5264 24259 5316 24268
rect 5264 24225 5273 24259
rect 5273 24225 5307 24259
rect 5307 24225 5316 24259
rect 5264 24216 5316 24225
rect 5448 24259 5500 24268
rect 5448 24225 5457 24259
rect 5457 24225 5491 24259
rect 5491 24225 5500 24259
rect 5448 24216 5500 24225
rect 10048 24284 10100 24336
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 2780 24148 2832 24200
rect 6368 24148 6420 24200
rect 7196 24148 7248 24200
rect 8300 24216 8352 24268
rect 7380 24191 7432 24200
rect 7380 24157 7389 24191
rect 7389 24157 7423 24191
rect 7423 24157 7432 24191
rect 7380 24148 7432 24157
rect 9772 24191 9824 24200
rect 9772 24157 9817 24191
rect 9817 24157 9824 24191
rect 9772 24148 9824 24157
rect 9956 24191 10008 24200
rect 9956 24157 9965 24191
rect 9965 24157 9999 24191
rect 9999 24157 10008 24191
rect 9956 24148 10008 24157
rect 10876 24216 10928 24268
rect 10508 24191 10560 24200
rect 10508 24157 10553 24191
rect 10553 24157 10560 24191
rect 10508 24148 10560 24157
rect 10692 24191 10744 24200
rect 10692 24157 10701 24191
rect 10701 24157 10735 24191
rect 10735 24157 10744 24191
rect 10692 24148 10744 24157
rect 11520 24216 11572 24268
rect 11980 24284 12032 24336
rect 12624 24352 12676 24404
rect 13268 24352 13320 24404
rect 13176 24284 13228 24336
rect 13728 24352 13780 24404
rect 14464 24352 14516 24404
rect 17868 24352 17920 24404
rect 19156 24352 19208 24404
rect 19800 24352 19852 24404
rect 20536 24352 20588 24404
rect 20996 24352 21048 24404
rect 21364 24395 21416 24404
rect 21364 24361 21373 24395
rect 21373 24361 21407 24395
rect 21407 24361 21416 24395
rect 21364 24352 21416 24361
rect 24032 24352 24084 24404
rect 26056 24352 26108 24404
rect 26240 24352 26292 24404
rect 26516 24352 26568 24404
rect 26608 24395 26660 24404
rect 26608 24361 26617 24395
rect 26617 24361 26651 24395
rect 26651 24361 26660 24395
rect 26608 24352 26660 24361
rect 5356 24080 5408 24132
rect 5540 24080 5592 24132
rect 5816 24123 5868 24132
rect 5816 24089 5825 24123
rect 5825 24089 5859 24123
rect 5859 24089 5868 24123
rect 5816 24080 5868 24089
rect 6000 24123 6052 24132
rect 6000 24089 6009 24123
rect 6009 24089 6043 24123
rect 6043 24089 6052 24123
rect 6000 24080 6052 24089
rect 6276 24080 6328 24132
rect 6552 24080 6604 24132
rect 6920 24012 6972 24064
rect 9588 24123 9640 24132
rect 9588 24089 9597 24123
rect 9597 24089 9631 24123
rect 9631 24089 9640 24123
rect 9588 24080 9640 24089
rect 9680 24123 9732 24132
rect 9680 24089 9689 24123
rect 9689 24089 9723 24123
rect 9723 24089 9732 24123
rect 9680 24080 9732 24089
rect 11980 24148 12032 24200
rect 11336 24123 11388 24132
rect 11336 24089 11345 24123
rect 11345 24089 11379 24123
rect 11379 24089 11388 24123
rect 11336 24080 11388 24089
rect 12992 24191 13044 24200
rect 12992 24157 13001 24191
rect 13001 24157 13035 24191
rect 13035 24157 13044 24191
rect 12992 24148 13044 24157
rect 13084 24191 13136 24200
rect 13084 24157 13094 24191
rect 13094 24157 13128 24191
rect 13128 24157 13136 24191
rect 13084 24148 13136 24157
rect 13268 24191 13320 24200
rect 13268 24157 13277 24191
rect 13277 24157 13311 24191
rect 13311 24157 13320 24191
rect 13268 24148 13320 24157
rect 16028 24284 16080 24336
rect 14740 24148 14792 24200
rect 14832 24191 14884 24200
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 16488 24216 16540 24268
rect 17592 24327 17644 24336
rect 17592 24293 17601 24327
rect 17601 24293 17635 24327
rect 17635 24293 17644 24327
rect 17592 24284 17644 24293
rect 17776 24284 17828 24336
rect 17960 24216 18012 24268
rect 18052 24216 18104 24268
rect 15844 24148 15896 24200
rect 12624 24123 12676 24132
rect 12624 24089 12633 24123
rect 12633 24089 12667 24123
rect 12667 24089 12676 24123
rect 12624 24080 12676 24089
rect 13728 24080 13780 24132
rect 14648 24123 14700 24132
rect 14648 24089 14657 24123
rect 14657 24089 14691 24123
rect 14691 24089 14700 24123
rect 14648 24080 14700 24089
rect 15016 24080 15068 24132
rect 17224 24080 17276 24132
rect 17776 24080 17828 24132
rect 18788 24191 18840 24200
rect 18788 24157 18797 24191
rect 18797 24157 18831 24191
rect 18831 24157 18840 24191
rect 18788 24148 18840 24157
rect 18972 24191 19024 24200
rect 18972 24157 18981 24191
rect 18981 24157 19015 24191
rect 19015 24157 19024 24191
rect 18972 24148 19024 24157
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20904 24284 20956 24336
rect 19892 24259 19944 24268
rect 19892 24225 19901 24259
rect 19901 24225 19935 24259
rect 19935 24225 19944 24259
rect 19892 24216 19944 24225
rect 21824 24284 21876 24336
rect 23388 24216 23440 24268
rect 20812 24191 20864 24200
rect 20812 24157 20821 24191
rect 20821 24157 20855 24191
rect 20855 24157 20864 24191
rect 20812 24148 20864 24157
rect 20904 24191 20956 24200
rect 20904 24157 20913 24191
rect 20913 24157 20947 24191
rect 20947 24157 20956 24191
rect 20904 24148 20956 24157
rect 21640 24148 21692 24200
rect 23204 24148 23256 24200
rect 24308 24148 24360 24200
rect 19800 24080 19852 24132
rect 20628 24123 20680 24132
rect 20628 24089 20637 24123
rect 20637 24089 20671 24123
rect 20671 24089 20680 24123
rect 20628 24080 20680 24089
rect 21088 24080 21140 24132
rect 23664 24080 23716 24132
rect 12256 24012 12308 24064
rect 14096 24012 14148 24064
rect 17592 24012 17644 24064
rect 19156 24012 19208 24064
rect 19248 24055 19300 24064
rect 19248 24021 19257 24055
rect 19257 24021 19291 24055
rect 19291 24021 19300 24055
rect 19248 24012 19300 24021
rect 19892 24012 19944 24064
rect 20352 24012 20404 24064
rect 20536 24055 20588 24064
rect 20536 24021 20545 24055
rect 20545 24021 20579 24055
rect 20579 24021 20588 24055
rect 20536 24012 20588 24021
rect 21916 24012 21968 24064
rect 24216 24012 24268 24064
rect 24860 24123 24912 24132
rect 24860 24089 24869 24123
rect 24869 24089 24903 24123
rect 24903 24089 24912 24123
rect 24860 24080 24912 24089
rect 25136 24191 25188 24200
rect 25136 24157 25145 24191
rect 25145 24157 25179 24191
rect 25179 24157 25188 24191
rect 25136 24148 25188 24157
rect 25780 24148 25832 24200
rect 25964 24148 26016 24200
rect 26608 24216 26660 24268
rect 26976 24352 27028 24404
rect 27804 24352 27856 24404
rect 27896 24395 27948 24404
rect 27896 24361 27905 24395
rect 27905 24361 27939 24395
rect 27939 24361 27948 24395
rect 27896 24352 27948 24361
rect 28816 24352 28868 24404
rect 27528 24284 27580 24336
rect 30288 24284 30340 24336
rect 26424 24191 26476 24200
rect 26424 24157 26433 24191
rect 26433 24157 26467 24191
rect 26467 24157 26476 24191
rect 26424 24148 26476 24157
rect 25228 24080 25280 24132
rect 26240 24123 26292 24132
rect 26240 24089 26249 24123
rect 26249 24089 26283 24123
rect 26283 24089 26292 24123
rect 26240 24080 26292 24089
rect 26884 24123 26936 24132
rect 26884 24089 26893 24123
rect 26893 24089 26927 24123
rect 26927 24089 26936 24123
rect 26884 24080 26936 24089
rect 26424 24012 26476 24064
rect 26516 24012 26568 24064
rect 27160 24148 27212 24200
rect 27528 24191 27580 24200
rect 27528 24157 27537 24191
rect 27537 24157 27571 24191
rect 27571 24157 27580 24191
rect 27528 24148 27580 24157
rect 27804 24216 27856 24268
rect 30012 24216 30064 24268
rect 28264 24148 28316 24200
rect 29276 24148 29328 24200
rect 30656 24191 30708 24200
rect 30656 24157 30665 24191
rect 30665 24157 30699 24191
rect 30699 24157 30708 24191
rect 30656 24148 30708 24157
rect 27620 24123 27672 24132
rect 27620 24089 27629 24123
rect 27629 24089 27663 24123
rect 27663 24089 27672 24123
rect 27620 24080 27672 24089
rect 28172 24080 28224 24132
rect 30932 24284 30984 24336
rect 31760 24395 31812 24404
rect 31760 24361 31769 24395
rect 31769 24361 31803 24395
rect 31803 24361 31812 24395
rect 31760 24352 31812 24361
rect 36176 24352 36228 24404
rect 31852 24284 31904 24336
rect 31024 24191 31076 24200
rect 31024 24157 31033 24191
rect 31033 24157 31067 24191
rect 31067 24157 31076 24191
rect 31024 24148 31076 24157
rect 30932 24123 30984 24132
rect 30932 24089 30941 24123
rect 30941 24089 30975 24123
rect 30975 24089 30984 24123
rect 30932 24080 30984 24089
rect 31300 24123 31352 24132
rect 31300 24089 31309 24123
rect 31309 24089 31343 24123
rect 31343 24089 31352 24123
rect 31300 24080 31352 24089
rect 31760 24216 31812 24268
rect 31576 24191 31628 24200
rect 31576 24157 31585 24191
rect 31585 24157 31619 24191
rect 31619 24157 31628 24191
rect 31576 24148 31628 24157
rect 36084 24191 36136 24200
rect 36084 24157 36093 24191
rect 36093 24157 36127 24191
rect 36127 24157 36136 24191
rect 36084 24148 36136 24157
rect 33416 24080 33468 24132
rect 29276 24012 29328 24064
rect 30840 24012 30892 24064
rect 31576 24012 31628 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 6092 23808 6144 23860
rect 8944 23808 8996 23860
rect 4068 23740 4120 23792
rect 5356 23783 5408 23792
rect 5356 23749 5365 23783
rect 5365 23749 5399 23783
rect 5399 23749 5408 23783
rect 5356 23740 5408 23749
rect 2964 23672 3016 23724
rect 4804 23672 4856 23724
rect 1400 23604 1452 23656
rect 1860 23647 1912 23656
rect 1860 23613 1869 23647
rect 1869 23613 1903 23647
rect 1903 23613 1912 23647
rect 1860 23604 1912 23613
rect 2412 23604 2464 23656
rect 5356 23536 5408 23588
rect 2044 23468 2096 23520
rect 2872 23468 2924 23520
rect 4712 23468 4764 23520
rect 5264 23468 5316 23520
rect 5816 23672 5868 23724
rect 12256 23808 12308 23860
rect 12808 23808 12860 23860
rect 14832 23808 14884 23860
rect 15016 23808 15068 23860
rect 15660 23851 15712 23860
rect 15660 23817 15669 23851
rect 15669 23817 15703 23851
rect 15703 23817 15712 23851
rect 15660 23808 15712 23817
rect 16396 23808 16448 23860
rect 17684 23808 17736 23860
rect 5632 23604 5684 23656
rect 5724 23604 5776 23656
rect 6460 23715 6512 23724
rect 6460 23681 6470 23715
rect 6470 23681 6504 23715
rect 6504 23681 6512 23715
rect 6460 23672 6512 23681
rect 6920 23672 6972 23724
rect 7380 23672 7432 23724
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 8300 23715 8352 23724
rect 8300 23681 8309 23715
rect 8309 23681 8343 23715
rect 8343 23681 8352 23715
rect 8300 23672 8352 23681
rect 9128 23740 9180 23792
rect 9312 23740 9364 23792
rect 7196 23604 7248 23656
rect 10508 23672 10560 23724
rect 11060 23604 11112 23656
rect 11888 23783 11940 23792
rect 11888 23749 11897 23783
rect 11897 23749 11931 23783
rect 11931 23749 11940 23783
rect 11888 23740 11940 23749
rect 11980 23740 12032 23792
rect 12808 23672 12860 23724
rect 13176 23715 13228 23724
rect 13176 23681 13180 23715
rect 13180 23681 13214 23715
rect 13214 23681 13228 23715
rect 13176 23672 13228 23681
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 13360 23715 13412 23724
rect 13360 23681 13369 23715
rect 13369 23681 13403 23715
rect 13403 23681 13412 23715
rect 13360 23672 13412 23681
rect 13544 23715 13596 23724
rect 13544 23681 13552 23715
rect 13552 23681 13586 23715
rect 13586 23681 13596 23715
rect 13544 23672 13596 23681
rect 13636 23715 13688 23724
rect 13636 23681 13645 23715
rect 13645 23681 13679 23715
rect 13679 23681 13688 23715
rect 13636 23672 13688 23681
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 15936 23740 15988 23792
rect 17868 23783 17920 23792
rect 17868 23749 17877 23783
rect 17877 23749 17911 23783
rect 17911 23749 17920 23783
rect 17868 23740 17920 23749
rect 18144 23808 18196 23860
rect 15844 23672 15896 23724
rect 19248 23740 19300 23792
rect 19616 23740 19668 23792
rect 19892 23740 19944 23792
rect 20628 23808 20680 23860
rect 24860 23808 24912 23860
rect 23940 23740 23992 23792
rect 25136 23740 25188 23792
rect 27252 23808 27304 23860
rect 12348 23604 12400 23656
rect 5632 23468 5684 23520
rect 5908 23511 5960 23520
rect 5908 23477 5917 23511
rect 5917 23477 5951 23511
rect 5951 23477 5960 23511
rect 5908 23468 5960 23477
rect 6276 23468 6328 23520
rect 6460 23536 6512 23588
rect 6644 23536 6696 23588
rect 7380 23536 7432 23588
rect 14740 23536 14792 23588
rect 17040 23536 17092 23588
rect 17776 23536 17828 23588
rect 18696 23672 18748 23724
rect 19340 23672 19392 23724
rect 18972 23647 19024 23656
rect 18972 23613 18981 23647
rect 18981 23613 19015 23647
rect 19015 23613 19024 23647
rect 18972 23604 19024 23613
rect 19248 23604 19300 23656
rect 20628 23672 20680 23724
rect 20720 23672 20772 23724
rect 22100 23672 22152 23724
rect 22376 23672 22428 23724
rect 28356 23740 28408 23792
rect 31852 23808 31904 23860
rect 32128 23808 32180 23860
rect 32404 23808 32456 23860
rect 20996 23647 21048 23656
rect 20996 23613 21005 23647
rect 21005 23613 21039 23647
rect 21039 23613 21048 23647
rect 20996 23604 21048 23613
rect 21088 23647 21140 23656
rect 21088 23613 21097 23647
rect 21097 23613 21131 23647
rect 21131 23613 21140 23647
rect 21088 23604 21140 23613
rect 21364 23604 21416 23656
rect 7196 23468 7248 23520
rect 7564 23468 7616 23520
rect 8116 23468 8168 23520
rect 11336 23468 11388 23520
rect 11704 23511 11756 23520
rect 11704 23477 11713 23511
rect 11713 23477 11747 23511
rect 11747 23477 11756 23511
rect 11704 23468 11756 23477
rect 12256 23468 12308 23520
rect 13084 23468 13136 23520
rect 13544 23468 13596 23520
rect 17408 23468 17460 23520
rect 17868 23511 17920 23520
rect 17868 23477 17877 23511
rect 17877 23477 17911 23511
rect 17911 23477 17920 23511
rect 17868 23468 17920 23477
rect 18144 23468 18196 23520
rect 19156 23536 19208 23588
rect 18972 23511 19024 23520
rect 18972 23477 18981 23511
rect 18981 23477 19015 23511
rect 19015 23477 19024 23511
rect 18972 23468 19024 23477
rect 25044 23604 25096 23656
rect 25596 23672 25648 23724
rect 22100 23536 22152 23588
rect 20720 23468 20772 23520
rect 21640 23468 21692 23520
rect 25780 23604 25832 23656
rect 26516 23672 26568 23724
rect 28540 23715 28592 23724
rect 28540 23681 28549 23715
rect 28549 23681 28583 23715
rect 28583 23681 28592 23715
rect 28540 23672 28592 23681
rect 28816 23715 28868 23724
rect 28816 23681 28825 23715
rect 28825 23681 28859 23715
rect 28859 23681 28868 23715
rect 28816 23672 28868 23681
rect 28264 23604 28316 23656
rect 29184 23715 29236 23724
rect 29184 23681 29193 23715
rect 29193 23681 29227 23715
rect 29227 23681 29236 23715
rect 29184 23672 29236 23681
rect 30564 23740 30616 23792
rect 26608 23536 26660 23588
rect 26884 23536 26936 23588
rect 29644 23604 29696 23656
rect 31024 23715 31076 23724
rect 31024 23681 31033 23715
rect 31033 23681 31067 23715
rect 31067 23681 31076 23715
rect 31024 23672 31076 23681
rect 31116 23672 31168 23724
rect 31300 23604 31352 23656
rect 31484 23672 31536 23724
rect 34152 23740 34204 23792
rect 32864 23604 32916 23656
rect 33048 23647 33100 23656
rect 33048 23613 33057 23647
rect 33057 23613 33091 23647
rect 33091 23613 33100 23647
rect 33048 23604 33100 23613
rect 34428 23715 34480 23724
rect 34428 23681 34437 23715
rect 34437 23681 34471 23715
rect 34471 23681 34480 23715
rect 34428 23672 34480 23681
rect 34612 23715 34664 23724
rect 34612 23681 34621 23715
rect 34621 23681 34655 23715
rect 34655 23681 34664 23715
rect 34612 23672 34664 23681
rect 34796 23604 34848 23656
rect 26056 23468 26108 23520
rect 26240 23468 26292 23520
rect 28908 23468 28960 23520
rect 29276 23468 29328 23520
rect 31116 23468 31168 23520
rect 31760 23468 31812 23520
rect 32772 23468 32824 23520
rect 33140 23511 33192 23520
rect 33140 23477 33149 23511
rect 33149 23477 33183 23511
rect 33183 23477 33192 23511
rect 33140 23468 33192 23477
rect 34612 23536 34664 23588
rect 34796 23468 34848 23520
rect 35440 23468 35492 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4252 23264 4304 23316
rect 5908 23264 5960 23316
rect 6000 23264 6052 23316
rect 6368 23264 6420 23316
rect 7196 23264 7248 23316
rect 9128 23264 9180 23316
rect 11980 23264 12032 23316
rect 3884 23196 3936 23248
rect 2412 23128 2464 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 3332 23128 3384 23180
rect 4252 23128 4304 23180
rect 3976 23060 4028 23112
rect 4528 23060 4580 23112
rect 5172 23103 5224 23112
rect 5172 23069 5181 23103
rect 5181 23069 5215 23103
rect 5215 23069 5224 23103
rect 5172 23060 5224 23069
rect 5632 23103 5684 23114
rect 1676 23035 1728 23044
rect 1676 23001 1685 23035
rect 1685 23001 1719 23035
rect 1719 23001 1728 23035
rect 1676 22992 1728 23001
rect 2964 22992 3016 23044
rect 4620 22992 4672 23044
rect 4804 22992 4856 23044
rect 5632 23069 5641 23103
rect 5641 23069 5675 23103
rect 5675 23069 5684 23103
rect 5632 23062 5684 23069
rect 6920 23196 6972 23248
rect 10324 23196 10376 23248
rect 10968 23196 11020 23248
rect 13176 23264 13228 23316
rect 17040 23307 17092 23316
rect 17040 23273 17049 23307
rect 17049 23273 17083 23307
rect 17083 23273 17092 23307
rect 17040 23264 17092 23273
rect 6644 23128 6696 23180
rect 3700 22924 3752 22976
rect 4068 22924 4120 22976
rect 4252 22967 4304 22976
rect 4252 22933 4261 22967
rect 4261 22933 4295 22967
rect 4295 22933 4304 22967
rect 4252 22924 4304 22933
rect 5080 22924 5132 22976
rect 5632 22924 5684 22976
rect 6000 23035 6052 23044
rect 6000 23001 6009 23035
rect 6009 23001 6043 23035
rect 6043 23001 6052 23035
rect 6000 22992 6052 23001
rect 6920 23060 6972 23112
rect 7196 23103 7248 23112
rect 7196 23069 7206 23103
rect 7206 23069 7240 23103
rect 7240 23069 7248 23103
rect 7196 23060 7248 23069
rect 8208 23128 8260 23180
rect 8392 23103 8444 23112
rect 8392 23069 8401 23103
rect 8401 23069 8435 23103
rect 8435 23069 8444 23103
rect 8392 23060 8444 23069
rect 6644 22992 6696 23044
rect 7380 23035 7432 23044
rect 7380 23001 7389 23035
rect 7389 23001 7423 23035
rect 7423 23001 7432 23035
rect 7380 22992 7432 23001
rect 7840 22924 7892 22976
rect 8484 23035 8536 23044
rect 8484 23001 8493 23035
rect 8493 23001 8527 23035
rect 8527 23001 8536 23035
rect 8484 22992 8536 23001
rect 8760 23103 8812 23112
rect 8760 23069 8769 23103
rect 8769 23069 8803 23103
rect 8803 23069 8812 23103
rect 8760 23060 8812 23069
rect 9588 23128 9640 23180
rect 11152 23171 11204 23180
rect 11152 23137 11161 23171
rect 11161 23137 11195 23171
rect 11195 23137 11204 23171
rect 11152 23128 11204 23137
rect 11060 23060 11112 23112
rect 11336 23103 11388 23112
rect 11336 23069 11352 23103
rect 11352 23069 11386 23103
rect 11386 23069 11388 23103
rect 11336 23060 11388 23069
rect 11520 23103 11572 23112
rect 11520 23069 11527 23103
rect 11527 23069 11572 23103
rect 11520 23060 11572 23069
rect 12256 23196 12308 23248
rect 14280 23196 14332 23248
rect 14556 23196 14608 23248
rect 16488 23196 16540 23248
rect 17592 23307 17644 23316
rect 17592 23273 17601 23307
rect 17601 23273 17635 23307
rect 17635 23273 17644 23307
rect 17592 23264 17644 23273
rect 17684 23264 17736 23316
rect 18236 23196 18288 23248
rect 13452 23128 13504 23180
rect 14740 23128 14792 23180
rect 11980 23060 12032 23112
rect 12348 23060 12400 23112
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 11612 23035 11664 23044
rect 11612 23001 11621 23035
rect 11621 23001 11655 23035
rect 11655 23001 11664 23035
rect 11612 22992 11664 23001
rect 8576 22924 8628 22976
rect 8760 22924 8812 22976
rect 9404 22924 9456 22976
rect 9956 22924 10008 22976
rect 10324 22924 10376 22976
rect 11060 22924 11112 22976
rect 11888 22992 11940 23044
rect 12532 22992 12584 23044
rect 12808 22992 12860 23044
rect 13820 22992 13872 23044
rect 14372 23060 14424 23112
rect 14556 23060 14608 23112
rect 15844 23128 15896 23180
rect 17960 23128 18012 23180
rect 19340 23264 19392 23316
rect 20536 23264 20588 23316
rect 20996 23264 21048 23316
rect 21640 23307 21692 23316
rect 21640 23273 21649 23307
rect 21649 23273 21683 23307
rect 21683 23273 21692 23307
rect 21640 23264 21692 23273
rect 23388 23264 23440 23316
rect 25228 23264 25280 23316
rect 27620 23264 27672 23316
rect 29184 23264 29236 23316
rect 32588 23264 32640 23316
rect 33968 23264 34020 23316
rect 25320 23196 25372 23248
rect 25872 23196 25924 23248
rect 26516 23196 26568 23248
rect 18880 23128 18932 23180
rect 19248 23128 19300 23180
rect 19340 23128 19392 23180
rect 20628 23128 20680 23180
rect 21640 23128 21692 23180
rect 15016 23103 15068 23112
rect 15016 23069 15025 23103
rect 15025 23069 15059 23103
rect 15059 23069 15068 23103
rect 15016 23060 15068 23069
rect 15660 23060 15712 23112
rect 15200 22992 15252 23044
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 16304 23060 16356 23112
rect 16856 23103 16908 23112
rect 16856 23069 16865 23103
rect 16865 23069 16899 23103
rect 16899 23069 16908 23103
rect 16856 23060 16908 23069
rect 16948 23103 17000 23112
rect 16948 23069 16957 23103
rect 16957 23069 16991 23103
rect 16991 23069 17000 23103
rect 16948 23060 17000 23069
rect 18696 23060 18748 23112
rect 19616 23060 19668 23112
rect 17040 22992 17092 23044
rect 17776 23035 17828 23044
rect 17776 23001 17785 23035
rect 17785 23001 17819 23035
rect 17819 23001 17828 23035
rect 17776 22992 17828 23001
rect 18604 22992 18656 23044
rect 11980 22967 12032 22976
rect 11980 22933 11989 22967
rect 11989 22933 12023 22967
rect 12023 22933 12032 22967
rect 11980 22924 12032 22933
rect 12072 22924 12124 22976
rect 12164 22967 12216 22976
rect 12164 22933 12173 22967
rect 12173 22933 12207 22967
rect 12207 22933 12216 22967
rect 12164 22924 12216 22933
rect 12900 22967 12952 22976
rect 12900 22933 12909 22967
rect 12909 22933 12943 22967
rect 12943 22933 12952 22967
rect 12900 22924 12952 22933
rect 13728 22924 13780 22976
rect 15752 22924 15804 22976
rect 17684 22924 17736 22976
rect 18144 22967 18196 22976
rect 18144 22933 18153 22967
rect 18153 22933 18187 22967
rect 18187 22933 18196 22967
rect 18144 22924 18196 22933
rect 21916 23060 21968 23112
rect 22008 23035 22060 23044
rect 22008 23001 22017 23035
rect 22017 23001 22051 23035
rect 22051 23001 22060 23035
rect 22008 22992 22060 23001
rect 22100 23035 22152 23044
rect 22100 23001 22109 23035
rect 22109 23001 22143 23035
rect 22143 23001 22152 23035
rect 22100 22992 22152 23001
rect 22560 23060 22612 23112
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 24216 23060 24268 23112
rect 25780 23103 25832 23112
rect 25780 23069 25789 23103
rect 25789 23069 25823 23103
rect 25823 23069 25832 23103
rect 25780 23060 25832 23069
rect 25872 23103 25924 23112
rect 25872 23069 25881 23103
rect 25881 23069 25915 23103
rect 25915 23069 25924 23103
rect 25872 23060 25924 23069
rect 27620 23060 27672 23112
rect 28264 23103 28316 23112
rect 28264 23069 28273 23103
rect 28273 23069 28307 23103
rect 28307 23069 28316 23103
rect 28264 23060 28316 23069
rect 24124 22992 24176 23044
rect 25596 22992 25648 23044
rect 27068 22992 27120 23044
rect 28172 23035 28224 23044
rect 28172 23001 28181 23035
rect 28181 23001 28215 23035
rect 28215 23001 28224 23035
rect 28172 22992 28224 23001
rect 22560 22924 22612 22976
rect 22652 22967 22704 22976
rect 22652 22933 22661 22967
rect 22661 22933 22695 22967
rect 22695 22933 22704 22967
rect 22652 22924 22704 22933
rect 30564 22924 30616 22976
rect 31024 22924 31076 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 1860 22720 1912 22772
rect 4712 22720 4764 22772
rect 4896 22720 4948 22772
rect 4068 22695 4120 22704
rect 4068 22661 4077 22695
rect 4077 22661 4111 22695
rect 4111 22661 4120 22695
rect 4068 22652 4120 22661
rect 4160 22652 4212 22704
rect 6828 22720 6880 22772
rect 6920 22763 6972 22772
rect 6920 22729 6929 22763
rect 6929 22729 6963 22763
rect 6963 22729 6972 22763
rect 6920 22720 6972 22729
rect 8208 22720 8260 22772
rect 6552 22695 6604 22704
rect 2504 22584 2556 22636
rect 2964 22584 3016 22636
rect 4344 22627 4396 22636
rect 4344 22593 4353 22627
rect 4353 22593 4387 22627
rect 4387 22593 4396 22627
rect 4344 22584 4396 22593
rect 5264 22584 5316 22636
rect 3332 22516 3384 22568
rect 3700 22516 3752 22568
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 5816 22627 5868 22636
rect 5816 22593 5825 22627
rect 5825 22593 5859 22627
rect 5859 22593 5868 22627
rect 5816 22584 5868 22593
rect 6552 22661 6561 22695
rect 6561 22661 6595 22695
rect 6595 22661 6604 22695
rect 6552 22652 6604 22661
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 6092 22584 6144 22636
rect 4344 22448 4396 22500
rect 5816 22448 5868 22500
rect 4068 22380 4120 22432
rect 4712 22380 4764 22432
rect 5264 22380 5316 22432
rect 7104 22559 7156 22568
rect 7104 22525 7113 22559
rect 7113 22525 7147 22559
rect 7147 22525 7156 22559
rect 7104 22516 7156 22525
rect 7380 22652 7432 22704
rect 8116 22695 8168 22704
rect 8116 22661 8125 22695
rect 8125 22661 8159 22695
rect 8159 22661 8168 22695
rect 8116 22652 8168 22661
rect 7840 22627 7892 22636
rect 7840 22593 7849 22627
rect 7849 22593 7883 22627
rect 7883 22593 7892 22627
rect 7840 22584 7892 22593
rect 8208 22627 8260 22636
rect 8208 22593 8217 22627
rect 8217 22593 8251 22627
rect 8251 22593 8260 22627
rect 8208 22584 8260 22593
rect 7656 22559 7708 22568
rect 7656 22525 7665 22559
rect 7665 22525 7699 22559
rect 7699 22525 7708 22559
rect 7656 22516 7708 22525
rect 8116 22516 8168 22568
rect 6828 22448 6880 22500
rect 9128 22652 9180 22704
rect 10048 22720 10100 22772
rect 10232 22763 10284 22772
rect 10232 22729 10241 22763
rect 10241 22729 10275 22763
rect 10275 22729 10284 22763
rect 10232 22720 10284 22729
rect 10324 22763 10376 22772
rect 10324 22729 10333 22763
rect 10333 22729 10367 22763
rect 10367 22729 10376 22763
rect 10324 22720 10376 22729
rect 9772 22695 9824 22704
rect 9772 22661 9781 22695
rect 9781 22661 9815 22695
rect 9815 22661 9824 22695
rect 9772 22652 9824 22661
rect 10968 22695 11020 22704
rect 10968 22661 10977 22695
rect 10977 22661 11011 22695
rect 11011 22661 11020 22695
rect 10968 22652 11020 22661
rect 11336 22720 11388 22772
rect 11704 22720 11756 22772
rect 11888 22695 11940 22704
rect 11888 22661 11897 22695
rect 11897 22661 11931 22695
rect 11931 22661 11940 22695
rect 11888 22652 11940 22661
rect 12164 22720 12216 22772
rect 14648 22720 14700 22772
rect 15292 22763 15344 22772
rect 15292 22729 15301 22763
rect 15301 22729 15335 22763
rect 15335 22729 15344 22763
rect 15292 22720 15344 22729
rect 15936 22720 15988 22772
rect 16948 22720 17000 22772
rect 17500 22720 17552 22772
rect 19708 22720 19760 22772
rect 12624 22652 12676 22704
rect 12808 22652 12860 22704
rect 13176 22695 13228 22704
rect 13176 22661 13185 22695
rect 13185 22661 13219 22695
rect 13219 22661 13228 22695
rect 13176 22652 13228 22661
rect 13360 22652 13412 22704
rect 9036 22627 9088 22636
rect 9036 22593 9050 22627
rect 9050 22593 9084 22627
rect 9084 22593 9088 22627
rect 9036 22584 9088 22593
rect 9404 22516 9456 22568
rect 8576 22448 8628 22500
rect 9128 22448 9180 22500
rect 9680 22584 9732 22636
rect 11704 22584 11756 22636
rect 12164 22627 12216 22636
rect 12164 22593 12172 22627
rect 12172 22593 12206 22627
rect 12206 22593 12216 22627
rect 12164 22584 12216 22593
rect 13452 22627 13504 22636
rect 10416 22559 10468 22568
rect 10416 22525 10425 22559
rect 10425 22525 10459 22559
rect 10459 22525 10468 22559
rect 10416 22516 10468 22525
rect 10692 22559 10744 22568
rect 10692 22525 10701 22559
rect 10701 22525 10735 22559
rect 10735 22525 10744 22559
rect 10692 22516 10744 22525
rect 10968 22516 11020 22568
rect 11980 22516 12032 22568
rect 13452 22593 13460 22627
rect 13460 22593 13494 22627
rect 13494 22593 13504 22627
rect 13452 22584 13504 22593
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 13728 22516 13780 22568
rect 14280 22627 14332 22636
rect 14280 22593 14289 22627
rect 14289 22593 14323 22627
rect 14323 22593 14332 22627
rect 14280 22584 14332 22593
rect 14740 22652 14792 22704
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 15752 22584 15804 22636
rect 17868 22652 17920 22704
rect 19340 22652 19392 22704
rect 14832 22516 14884 22568
rect 15292 22516 15344 22568
rect 17960 22584 18012 22636
rect 18236 22627 18288 22636
rect 18236 22593 18245 22627
rect 18245 22593 18279 22627
rect 18279 22593 18288 22627
rect 18236 22584 18288 22593
rect 18420 22627 18472 22636
rect 18420 22593 18429 22627
rect 18429 22593 18463 22627
rect 18463 22593 18472 22627
rect 18420 22584 18472 22593
rect 19432 22584 19484 22636
rect 22836 22720 22888 22772
rect 25412 22763 25464 22772
rect 25412 22729 25421 22763
rect 25421 22729 25455 22763
rect 25455 22729 25464 22763
rect 25412 22720 25464 22729
rect 25596 22720 25648 22772
rect 10508 22448 10560 22500
rect 6092 22423 6144 22432
rect 6092 22389 6101 22423
rect 6101 22389 6135 22423
rect 6135 22389 6144 22423
rect 6092 22380 6144 22389
rect 6368 22380 6420 22432
rect 8208 22380 8260 22432
rect 11520 22380 11572 22432
rect 11612 22423 11664 22432
rect 11612 22389 11621 22423
rect 11621 22389 11655 22423
rect 11655 22389 11664 22423
rect 11612 22380 11664 22389
rect 12348 22448 12400 22500
rect 12532 22491 12584 22500
rect 12532 22457 12541 22491
rect 12541 22457 12575 22491
rect 12575 22457 12584 22491
rect 12532 22448 12584 22457
rect 15016 22448 15068 22500
rect 16488 22516 16540 22568
rect 18328 22516 18380 22568
rect 18604 22516 18656 22568
rect 18236 22448 18288 22500
rect 20904 22652 20956 22704
rect 22560 22695 22612 22704
rect 22560 22661 22569 22695
rect 22569 22661 22603 22695
rect 22603 22661 22612 22695
rect 22560 22652 22612 22661
rect 23204 22652 23256 22704
rect 32588 22720 32640 22772
rect 32680 22720 32732 22772
rect 20536 22627 20588 22636
rect 20536 22593 20545 22627
rect 20545 22593 20579 22627
rect 20579 22593 20588 22627
rect 20536 22584 20588 22593
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 22652 22584 22704 22636
rect 23480 22584 23532 22636
rect 23756 22627 23808 22636
rect 23756 22593 23765 22627
rect 23765 22593 23799 22627
rect 23799 22593 23808 22627
rect 23756 22584 23808 22593
rect 23940 22584 23992 22636
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24216 22627 24268 22636
rect 24216 22593 24225 22627
rect 24225 22593 24259 22627
rect 24259 22593 24268 22627
rect 24216 22584 24268 22593
rect 24400 22627 24452 22636
rect 24400 22593 24408 22627
rect 24408 22593 24442 22627
rect 24442 22593 24452 22627
rect 24400 22584 24452 22593
rect 24308 22516 24360 22568
rect 36268 22720 36320 22772
rect 33048 22652 33100 22704
rect 25596 22627 25648 22636
rect 25596 22593 25605 22627
rect 25605 22593 25639 22627
rect 25639 22593 25648 22627
rect 25596 22584 25648 22593
rect 25688 22584 25740 22636
rect 28080 22584 28132 22636
rect 28724 22584 28776 22636
rect 31852 22584 31904 22636
rect 25412 22516 25464 22568
rect 25872 22516 25924 22568
rect 27804 22559 27856 22568
rect 27804 22525 27813 22559
rect 27813 22525 27847 22559
rect 27847 22525 27856 22559
rect 27804 22516 27856 22525
rect 30840 22516 30892 22568
rect 25688 22448 25740 22500
rect 30748 22448 30800 22500
rect 32772 22584 32824 22636
rect 34704 22584 34756 22636
rect 34796 22627 34848 22636
rect 34796 22593 34805 22627
rect 34805 22593 34839 22627
rect 34839 22593 34848 22627
rect 34796 22584 34848 22593
rect 36084 22627 36136 22636
rect 36084 22593 36093 22627
rect 36093 22593 36127 22627
rect 36127 22593 36136 22627
rect 36084 22584 36136 22593
rect 34612 22559 34664 22568
rect 34612 22525 34621 22559
rect 34621 22525 34655 22559
rect 34655 22525 34664 22559
rect 34612 22516 34664 22525
rect 13084 22380 13136 22432
rect 15568 22380 15620 22432
rect 16488 22380 16540 22432
rect 19892 22380 19944 22432
rect 20352 22380 20404 22432
rect 22468 22423 22520 22432
rect 22468 22389 22477 22423
rect 22477 22389 22511 22423
rect 22511 22389 22520 22423
rect 22468 22380 22520 22389
rect 23756 22423 23808 22432
rect 23756 22389 23765 22423
rect 23765 22389 23799 22423
rect 23799 22389 23808 22423
rect 23756 22380 23808 22389
rect 23940 22380 23992 22432
rect 27620 22380 27672 22432
rect 30288 22380 30340 22432
rect 33692 22423 33744 22432
rect 33692 22389 33701 22423
rect 33701 22389 33735 22423
rect 33735 22389 33744 22423
rect 33692 22380 33744 22389
rect 34796 22380 34848 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1676 22176 1728 22228
rect 4620 22176 4672 22228
rect 5724 22176 5776 22228
rect 6552 22176 6604 22228
rect 9680 22176 9732 22228
rect 9956 22176 10008 22228
rect 11796 22176 11848 22228
rect 12348 22176 12400 22228
rect 13544 22176 13596 22228
rect 2688 22108 2740 22160
rect 2780 22083 2832 22092
rect 2780 22049 2789 22083
rect 2789 22049 2823 22083
rect 2823 22049 2832 22083
rect 2780 22040 2832 22049
rect 5080 22108 5132 22160
rect 5540 22108 5592 22160
rect 7932 22108 7984 22160
rect 8760 22108 8812 22160
rect 3332 22040 3384 22092
rect 4068 22040 4120 22092
rect 5172 22040 5224 22092
rect 4620 21972 4672 22024
rect 5264 22015 5316 22024
rect 5264 21981 5273 22015
rect 5273 21981 5307 22015
rect 5307 21981 5316 22015
rect 5264 21972 5316 21981
rect 4712 21904 4764 21956
rect 4804 21904 4856 21956
rect 5908 22040 5960 22092
rect 8208 22083 8260 22092
rect 8208 22049 8217 22083
rect 8217 22049 8251 22083
rect 8251 22049 8260 22083
rect 8208 22040 8260 22049
rect 8484 22040 8536 22092
rect 8944 22040 8996 22092
rect 12808 22108 12860 22160
rect 13820 22219 13872 22228
rect 13820 22185 13829 22219
rect 13829 22185 13863 22219
rect 13863 22185 13872 22219
rect 13820 22176 13872 22185
rect 14832 22151 14884 22160
rect 14832 22117 14841 22151
rect 14841 22117 14875 22151
rect 14875 22117 14884 22151
rect 14832 22108 14884 22117
rect 7104 21972 7156 22024
rect 7472 22015 7524 22024
rect 7472 21981 7481 22015
rect 7481 21981 7515 22015
rect 7515 21981 7524 22015
rect 7472 21972 7524 21981
rect 7932 21972 7984 22024
rect 8300 21972 8352 22024
rect 10968 21972 11020 22024
rect 6460 21904 6512 21956
rect 5264 21836 5316 21888
rect 6552 21836 6604 21888
rect 8024 21904 8076 21956
rect 8576 21904 8628 21956
rect 9772 21904 9824 21956
rect 10600 21836 10652 21888
rect 11152 21836 11204 21888
rect 11336 22015 11388 22024
rect 11336 21981 11345 22015
rect 11345 21981 11379 22015
rect 11379 21981 11388 22015
rect 11336 21972 11388 21981
rect 11520 22015 11572 22024
rect 11520 21981 11529 22015
rect 11529 21981 11563 22015
rect 11563 21981 11572 22015
rect 11520 21972 11572 21981
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 11612 21972 11664 21981
rect 11796 22015 11848 22024
rect 11796 21981 11805 22015
rect 11805 21981 11839 22015
rect 11839 21981 11848 22015
rect 11796 21972 11848 21981
rect 11980 22015 12032 22024
rect 11980 21981 11989 22015
rect 11989 21981 12023 22015
rect 12023 21981 12032 22015
rect 11980 21972 12032 21981
rect 12164 21904 12216 21956
rect 12348 21904 12400 21956
rect 12900 21972 12952 22024
rect 13360 21972 13412 22024
rect 13452 22015 13504 22024
rect 13452 21981 13461 22015
rect 13461 21981 13495 22015
rect 13495 21981 13504 22015
rect 13452 21972 13504 21981
rect 13268 21904 13320 21956
rect 14740 21972 14792 22024
rect 15568 22108 15620 22160
rect 15752 22083 15804 22092
rect 15752 22049 15761 22083
rect 15761 22049 15795 22083
rect 15795 22049 15804 22083
rect 15752 22040 15804 22049
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 17224 22219 17276 22228
rect 17224 22185 17233 22219
rect 17233 22185 17267 22219
rect 17267 22185 17276 22219
rect 17224 22176 17276 22185
rect 17960 22176 18012 22228
rect 17316 22108 17368 22160
rect 19892 22108 19944 22160
rect 20720 22108 20772 22160
rect 21088 22108 21140 22160
rect 22468 22176 22520 22228
rect 23204 22176 23256 22228
rect 23756 22176 23808 22228
rect 24584 22176 24636 22228
rect 23020 22151 23072 22160
rect 23020 22117 23029 22151
rect 23029 22117 23063 22151
rect 23063 22117 23072 22151
rect 23020 22108 23072 22117
rect 21916 22040 21968 22092
rect 25136 22108 25188 22160
rect 26056 22083 26108 22092
rect 26056 22049 26065 22083
rect 26065 22049 26099 22083
rect 26099 22049 26108 22083
rect 26056 22040 26108 22049
rect 26332 22040 26384 22092
rect 27068 22040 27120 22092
rect 32128 22108 32180 22160
rect 32680 22108 32732 22160
rect 35348 22108 35400 22160
rect 27620 22040 27672 22092
rect 30288 22040 30340 22092
rect 30656 22040 30708 22092
rect 14832 21904 14884 21956
rect 15752 21904 15804 21956
rect 13820 21836 13872 21888
rect 15844 21836 15896 21888
rect 16488 21972 16540 22024
rect 18420 21972 18472 22024
rect 16396 21904 16448 21956
rect 19340 21904 19392 21956
rect 16212 21836 16264 21888
rect 18788 21836 18840 21888
rect 19800 21972 19852 22024
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 22100 21972 22152 22024
rect 22744 21972 22796 22024
rect 23112 21972 23164 22024
rect 20260 21904 20312 21956
rect 20996 21904 21048 21956
rect 26240 22015 26292 22024
rect 26240 21981 26249 22015
rect 26249 21981 26283 22015
rect 26283 21981 26292 22015
rect 26240 21972 26292 21981
rect 27160 21972 27212 22024
rect 28172 21972 28224 22024
rect 23756 21904 23808 21956
rect 26976 21904 27028 21956
rect 20168 21836 20220 21888
rect 22008 21836 22060 21888
rect 22468 21836 22520 21888
rect 25780 21836 25832 21888
rect 26240 21836 26292 21888
rect 26424 21879 26476 21888
rect 26424 21845 26433 21879
rect 26433 21845 26467 21879
rect 26467 21845 26476 21879
rect 26424 21836 26476 21845
rect 27804 21904 27856 21956
rect 29000 21972 29052 22024
rect 28540 21904 28592 21956
rect 30380 21947 30432 21956
rect 30380 21913 30389 21947
rect 30389 21913 30423 21947
rect 30423 21913 30432 21947
rect 30380 21904 30432 21913
rect 33324 21972 33376 22024
rect 34796 21972 34848 22024
rect 35992 21972 36044 22024
rect 36084 22015 36136 22024
rect 36084 21981 36093 22015
rect 36093 21981 36127 22015
rect 36127 21981 36136 22015
rect 36084 21972 36136 21981
rect 30748 21904 30800 21956
rect 27712 21836 27764 21888
rect 28172 21836 28224 21888
rect 30012 21879 30064 21888
rect 30012 21845 30021 21879
rect 30021 21845 30055 21879
rect 30055 21845 30064 21879
rect 30012 21836 30064 21845
rect 34244 21836 34296 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 2964 21564 3016 21616
rect 3424 21564 3476 21616
rect 4988 21632 5040 21684
rect 5816 21632 5868 21684
rect 4068 21539 4120 21548
rect 4068 21505 4077 21539
rect 4077 21505 4111 21539
rect 4111 21505 4120 21539
rect 4068 21496 4120 21505
rect 4712 21496 4764 21548
rect 5356 21496 5408 21548
rect 8576 21632 8628 21684
rect 6552 21564 6604 21616
rect 7104 21564 7156 21616
rect 8300 21564 8352 21616
rect 8392 21539 8444 21548
rect 8392 21505 8396 21539
rect 8396 21505 8430 21539
rect 8430 21505 8444 21539
rect 8392 21496 8444 21505
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 2136 21428 2188 21480
rect 5264 21428 5316 21480
rect 5540 21428 5592 21480
rect 8668 21496 8720 21548
rect 8760 21539 8812 21548
rect 8760 21505 8768 21539
rect 8768 21505 8802 21539
rect 8802 21505 8812 21539
rect 8760 21496 8812 21505
rect 9772 21564 9824 21616
rect 11152 21632 11204 21684
rect 11336 21632 11388 21684
rect 12716 21632 12768 21684
rect 13268 21632 13320 21684
rect 17224 21632 17276 21684
rect 11244 21564 11296 21616
rect 13084 21564 13136 21616
rect 14924 21564 14976 21616
rect 17316 21564 17368 21616
rect 8024 21360 8076 21412
rect 2780 21292 2832 21344
rect 4804 21292 4856 21344
rect 6736 21292 6788 21344
rect 7656 21292 7708 21344
rect 9772 21428 9824 21480
rect 11060 21428 11112 21480
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 11796 21539 11848 21548
rect 11796 21505 11805 21539
rect 11805 21505 11839 21539
rect 11839 21505 11848 21539
rect 11796 21496 11848 21505
rect 11980 21496 12032 21548
rect 14648 21496 14700 21548
rect 15568 21496 15620 21548
rect 16580 21496 16632 21548
rect 17684 21564 17736 21616
rect 17868 21564 17920 21616
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 12348 21428 12400 21480
rect 15200 21428 15252 21480
rect 18512 21539 18564 21548
rect 18512 21505 18521 21539
rect 18521 21505 18555 21539
rect 18555 21505 18564 21539
rect 18512 21496 18564 21505
rect 19524 21632 19576 21684
rect 20352 21675 20404 21684
rect 20352 21641 20361 21675
rect 20361 21641 20395 21675
rect 20395 21641 20404 21675
rect 20352 21632 20404 21641
rect 21640 21632 21692 21684
rect 24492 21632 24544 21684
rect 26332 21632 26384 21684
rect 29920 21632 29972 21684
rect 36452 21632 36504 21684
rect 19156 21496 19208 21548
rect 19248 21496 19300 21548
rect 19708 21539 19760 21548
rect 19708 21505 19717 21539
rect 19717 21505 19751 21539
rect 19751 21505 19760 21539
rect 19708 21496 19760 21505
rect 21088 21564 21140 21616
rect 20352 21496 20404 21548
rect 22008 21496 22060 21548
rect 24032 21607 24084 21616
rect 24032 21573 24041 21607
rect 24041 21573 24075 21607
rect 24075 21573 24084 21607
rect 24032 21564 24084 21573
rect 24216 21564 24268 21616
rect 28448 21564 28500 21616
rect 25504 21496 25556 21548
rect 28816 21539 28868 21548
rect 28816 21505 28825 21539
rect 28825 21505 28859 21539
rect 28859 21505 28868 21539
rect 28816 21496 28868 21505
rect 31208 21564 31260 21616
rect 29184 21539 29236 21548
rect 29184 21505 29193 21539
rect 29193 21505 29227 21539
rect 29227 21505 29236 21539
rect 29184 21496 29236 21505
rect 10324 21360 10376 21412
rect 11704 21360 11756 21412
rect 13268 21360 13320 21412
rect 14096 21360 14148 21412
rect 20076 21428 20128 21480
rect 20628 21428 20680 21480
rect 22376 21428 22428 21480
rect 24492 21428 24544 21480
rect 25136 21428 25188 21480
rect 11244 21292 11296 21344
rect 11336 21335 11388 21344
rect 11336 21301 11345 21335
rect 11345 21301 11379 21335
rect 11379 21301 11388 21335
rect 11336 21292 11388 21301
rect 11520 21335 11572 21344
rect 11520 21301 11529 21335
rect 11529 21301 11563 21335
rect 11563 21301 11572 21335
rect 11520 21292 11572 21301
rect 12532 21292 12584 21344
rect 13544 21292 13596 21344
rect 14464 21292 14516 21344
rect 17316 21335 17368 21344
rect 17316 21301 17325 21335
rect 17325 21301 17359 21335
rect 17359 21301 17368 21335
rect 17316 21292 17368 21301
rect 19340 21292 19392 21344
rect 22652 21360 22704 21412
rect 20904 21292 20956 21344
rect 23112 21292 23164 21344
rect 23664 21335 23716 21344
rect 23664 21301 23673 21335
rect 23673 21301 23707 21335
rect 23707 21301 23716 21335
rect 23664 21292 23716 21301
rect 26056 21360 26108 21412
rect 28540 21360 28592 21412
rect 27712 21292 27764 21344
rect 29552 21539 29604 21548
rect 29552 21505 29561 21539
rect 29561 21505 29595 21539
rect 29595 21505 29604 21539
rect 29552 21496 29604 21505
rect 30104 21496 30156 21548
rect 32772 21496 32824 21548
rect 36084 21539 36136 21548
rect 36084 21505 36093 21539
rect 36093 21505 36127 21539
rect 36127 21505 36136 21539
rect 36084 21496 36136 21505
rect 31208 21360 31260 21412
rect 30748 21292 30800 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2136 21131 2188 21140
rect 2136 21097 2145 21131
rect 2145 21097 2179 21131
rect 2179 21097 2188 21131
rect 2136 21088 2188 21097
rect 3056 21088 3108 21140
rect 6828 21088 6880 21140
rect 9772 21131 9824 21140
rect 9772 21097 9781 21131
rect 9781 21097 9815 21131
rect 9815 21097 9824 21131
rect 9772 21088 9824 21097
rect 10600 21088 10652 21140
rect 10784 21088 10836 21140
rect 11336 21088 11388 21140
rect 2872 21020 2924 21072
rect 2228 20952 2280 21004
rect 2688 20995 2740 21004
rect 2688 20961 2697 20995
rect 2697 20961 2731 20995
rect 2731 20961 2740 20995
rect 2688 20952 2740 20961
rect 2780 20884 2832 20936
rect 3056 20884 3108 20936
rect 6368 21020 6420 21072
rect 6920 21020 6972 21072
rect 4712 20952 4764 21004
rect 4620 20927 4672 20936
rect 4620 20893 4629 20927
rect 4629 20893 4663 20927
rect 4663 20893 4672 20927
rect 4620 20884 4672 20893
rect 5264 20952 5316 21004
rect 5356 20952 5408 21004
rect 7472 21063 7524 21072
rect 7472 21029 7481 21063
rect 7481 21029 7515 21063
rect 7515 21029 7524 21063
rect 7472 21020 7524 21029
rect 7656 21020 7708 21072
rect 9036 21020 9088 21072
rect 11060 21020 11112 21072
rect 4988 20927 5040 20936
rect 4988 20893 4997 20927
rect 4997 20893 5031 20927
rect 5031 20893 5040 20927
rect 4988 20884 5040 20893
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 7840 20884 7892 20936
rect 8392 20952 8444 21004
rect 8944 20952 8996 21004
rect 9404 20995 9456 21004
rect 9404 20961 9413 20995
rect 9413 20961 9447 20995
rect 9447 20961 9456 20995
rect 9404 20952 9456 20961
rect 8576 20816 8628 20868
rect 8760 20816 8812 20868
rect 9404 20816 9456 20868
rect 3240 20748 3292 20800
rect 4528 20748 4580 20800
rect 5264 20748 5316 20800
rect 7564 20748 7616 20800
rect 7748 20748 7800 20800
rect 8116 20791 8168 20800
rect 8116 20757 8125 20791
rect 8125 20757 8159 20791
rect 8159 20757 8168 20791
rect 8116 20748 8168 20757
rect 8944 20791 8996 20800
rect 8944 20757 8953 20791
rect 8953 20757 8987 20791
rect 8987 20757 8996 20791
rect 8944 20748 8996 20757
rect 9128 20748 9180 20800
rect 10508 20952 10560 21004
rect 11520 21063 11572 21072
rect 11520 21029 11529 21063
rect 11529 21029 11563 21063
rect 11563 21029 11572 21063
rect 11520 21020 11572 21029
rect 12072 21088 12124 21140
rect 12256 21088 12308 21140
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 11060 20884 11112 20936
rect 11704 20927 11756 20936
rect 11704 20893 11713 20927
rect 11713 20893 11747 20927
rect 11747 20893 11756 20927
rect 11704 20884 11756 20893
rect 10784 20816 10836 20868
rect 12256 20952 12308 21004
rect 12624 21020 12676 21072
rect 13360 21020 13412 21072
rect 13452 21020 13504 21072
rect 12624 20927 12676 20936
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 12532 20816 12584 20868
rect 12808 20816 12860 20868
rect 13268 20884 13320 20936
rect 13084 20859 13136 20868
rect 13084 20825 13093 20859
rect 13093 20825 13127 20859
rect 13127 20825 13136 20859
rect 13084 20816 13136 20825
rect 13360 20859 13412 20868
rect 13360 20825 13369 20859
rect 13369 20825 13403 20859
rect 13403 20825 13412 20859
rect 13360 20816 13412 20825
rect 13176 20748 13228 20800
rect 17132 21088 17184 21140
rect 17316 21088 17368 21140
rect 18512 21088 18564 21140
rect 19156 21088 19208 21140
rect 19708 21088 19760 21140
rect 20628 21088 20680 21140
rect 21916 21088 21968 21140
rect 22928 21131 22980 21140
rect 22928 21097 22937 21131
rect 22937 21097 22971 21131
rect 22971 21097 22980 21131
rect 22928 21088 22980 21097
rect 23572 21131 23624 21140
rect 23572 21097 23581 21131
rect 23581 21097 23615 21131
rect 23615 21097 23624 21131
rect 23572 21088 23624 21097
rect 23940 21131 23992 21140
rect 23940 21097 23949 21131
rect 23949 21097 23983 21131
rect 23983 21097 23992 21131
rect 23940 21088 23992 21097
rect 14188 20884 14240 20936
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 16396 21020 16448 21072
rect 19892 21020 19944 21072
rect 26332 21088 26384 21140
rect 26976 21088 27028 21140
rect 29000 21088 29052 21140
rect 29552 21088 29604 21140
rect 32772 21131 32824 21140
rect 32772 21097 32781 21131
rect 32781 21097 32815 21131
rect 32815 21097 32824 21131
rect 32772 21088 32824 21097
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 19524 20952 19576 21004
rect 19984 20952 20036 21004
rect 14096 20748 14148 20800
rect 15660 20884 15712 20936
rect 15936 20884 15988 20936
rect 17040 20927 17092 20936
rect 17040 20893 17049 20927
rect 17049 20893 17083 20927
rect 17083 20893 17092 20927
rect 17040 20884 17092 20893
rect 17960 20884 18012 20936
rect 16396 20816 16448 20868
rect 18236 20816 18288 20868
rect 19616 20816 19668 20868
rect 15660 20748 15712 20800
rect 15752 20791 15804 20800
rect 15752 20757 15761 20791
rect 15761 20757 15795 20791
rect 15795 20757 15804 20791
rect 15752 20748 15804 20757
rect 17868 20748 17920 20800
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 21456 20927 21508 20936
rect 21456 20893 21465 20927
rect 21465 20893 21499 20927
rect 21499 20893 21508 20927
rect 21456 20884 21508 20893
rect 21548 20927 21600 20936
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 21088 20816 21140 20868
rect 22192 20859 22244 20868
rect 22192 20825 22201 20859
rect 22201 20825 22235 20859
rect 22235 20825 22244 20859
rect 22192 20816 22244 20825
rect 23112 20859 23164 20868
rect 23112 20825 23121 20859
rect 23121 20825 23155 20859
rect 23155 20825 23164 20859
rect 23112 20816 23164 20825
rect 22100 20748 22152 20800
rect 22284 20748 22336 20800
rect 22836 20748 22888 20800
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 23664 20927 23716 20936
rect 23664 20893 23673 20927
rect 23673 20893 23707 20927
rect 23707 20893 23716 20927
rect 23664 20884 23716 20893
rect 24492 21020 24544 21072
rect 24584 21020 24636 21072
rect 24032 20927 24084 20936
rect 24032 20893 24041 20927
rect 24041 20893 24075 20927
rect 24075 20893 24084 20927
rect 24032 20884 24084 20893
rect 23480 20748 23532 20800
rect 23664 20748 23716 20800
rect 24492 20927 24544 20936
rect 24492 20893 24501 20927
rect 24501 20893 24535 20927
rect 24535 20893 24544 20927
rect 24492 20884 24544 20893
rect 24768 20927 24820 20936
rect 24768 20893 24777 20927
rect 24777 20893 24811 20927
rect 24811 20893 24820 20927
rect 24768 20884 24820 20893
rect 24952 20952 25004 21004
rect 25504 20927 25556 20936
rect 25504 20893 25513 20927
rect 25513 20893 25547 20927
rect 25547 20893 25556 20927
rect 25504 20884 25556 20893
rect 25320 20816 25372 20868
rect 26056 20816 26108 20868
rect 29368 21020 29420 21072
rect 31668 21020 31720 21072
rect 33140 21020 33192 21072
rect 27252 20952 27304 21004
rect 27988 20927 28040 20936
rect 27988 20893 27997 20927
rect 27997 20893 28031 20927
rect 28031 20893 28040 20927
rect 27988 20884 28040 20893
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 31208 20952 31260 21004
rect 31484 20927 31536 20936
rect 31484 20893 31493 20927
rect 31493 20893 31527 20927
rect 31527 20893 31536 20927
rect 31484 20884 31536 20893
rect 31668 20927 31720 20936
rect 31668 20893 31677 20927
rect 31677 20893 31711 20927
rect 31711 20893 31720 20927
rect 31668 20884 31720 20893
rect 31944 20884 31996 20936
rect 33048 20927 33100 20936
rect 33048 20893 33057 20927
rect 33057 20893 33091 20927
rect 33091 20893 33100 20927
rect 33048 20884 33100 20893
rect 27252 20816 27304 20868
rect 28172 20859 28224 20868
rect 28172 20825 28189 20859
rect 28189 20825 28224 20859
rect 28172 20816 28224 20825
rect 28264 20859 28316 20868
rect 28264 20825 28273 20859
rect 28273 20825 28307 20859
rect 28307 20825 28316 20859
rect 28264 20816 28316 20825
rect 32036 20816 32088 20868
rect 25780 20748 25832 20800
rect 26792 20748 26844 20800
rect 27712 20748 27764 20800
rect 28356 20748 28408 20800
rect 30288 20748 30340 20800
rect 31300 20791 31352 20800
rect 31300 20757 31309 20791
rect 31309 20757 31343 20791
rect 31343 20757 31352 20791
rect 31300 20748 31352 20757
rect 34612 20748 34664 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 2964 20544 3016 20596
rect 7104 20544 7156 20596
rect 7472 20544 7524 20596
rect 8116 20544 8168 20596
rect 9404 20544 9456 20596
rect 12072 20544 12124 20596
rect 13084 20587 13136 20596
rect 13084 20553 13093 20587
rect 13093 20553 13127 20587
rect 13127 20553 13136 20587
rect 13084 20544 13136 20553
rect 13360 20544 13412 20596
rect 4528 20451 4580 20460
rect 4528 20417 4537 20451
rect 4537 20417 4571 20451
rect 4571 20417 4580 20451
rect 4528 20408 4580 20417
rect 4896 20451 4948 20460
rect 4896 20417 4905 20451
rect 4905 20417 4939 20451
rect 4939 20417 4948 20451
rect 4896 20408 4948 20417
rect 5816 20408 5868 20460
rect 7288 20476 7340 20528
rect 8024 20476 8076 20528
rect 8944 20476 8996 20528
rect 9680 20476 9732 20528
rect 11428 20476 11480 20528
rect 14280 20476 14332 20528
rect 15016 20544 15068 20596
rect 21272 20544 21324 20596
rect 22192 20544 22244 20596
rect 24768 20544 24820 20596
rect 24952 20587 25004 20596
rect 24952 20553 24961 20587
rect 24961 20553 24995 20587
rect 24995 20553 25004 20587
rect 24952 20544 25004 20553
rect 25136 20544 25188 20596
rect 25780 20544 25832 20596
rect 7012 20451 7064 20460
rect 7012 20417 7021 20451
rect 7021 20417 7055 20451
rect 7055 20417 7064 20451
rect 7012 20408 7064 20417
rect 8208 20408 8260 20460
rect 4620 20340 4672 20392
rect 5632 20383 5684 20392
rect 5632 20349 5641 20383
rect 5641 20349 5675 20383
rect 5675 20349 5684 20383
rect 5632 20340 5684 20349
rect 7288 20383 7340 20392
rect 7288 20349 7297 20383
rect 7297 20349 7331 20383
rect 7331 20349 7340 20383
rect 7288 20340 7340 20349
rect 7656 20340 7708 20392
rect 7932 20340 7984 20392
rect 8116 20340 8168 20392
rect 6920 20272 6972 20324
rect 9680 20340 9732 20392
rect 10692 20408 10744 20460
rect 15752 20476 15804 20528
rect 15936 20519 15988 20528
rect 15936 20485 15945 20519
rect 15945 20485 15979 20519
rect 15979 20485 15988 20519
rect 15936 20476 15988 20485
rect 16120 20519 16172 20528
rect 16120 20485 16145 20519
rect 16145 20485 16172 20519
rect 16120 20476 16172 20485
rect 16488 20476 16540 20528
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 17592 20476 17644 20528
rect 18420 20408 18472 20460
rect 20352 20519 20404 20528
rect 20352 20485 20361 20519
rect 20361 20485 20395 20519
rect 20395 20485 20404 20519
rect 20352 20476 20404 20485
rect 20904 20519 20956 20528
rect 20904 20485 20913 20519
rect 20913 20485 20947 20519
rect 20947 20485 20956 20519
rect 20904 20476 20956 20485
rect 21364 20476 21416 20528
rect 21548 20476 21600 20528
rect 23388 20476 23440 20528
rect 24124 20476 24176 20528
rect 20076 20408 20128 20460
rect 12072 20340 12124 20392
rect 12532 20383 12584 20392
rect 12532 20349 12541 20383
rect 12541 20349 12575 20383
rect 12575 20349 12584 20383
rect 12532 20340 12584 20349
rect 14096 20340 14148 20392
rect 15016 20383 15068 20392
rect 15016 20349 15025 20383
rect 15025 20349 15059 20383
rect 15059 20349 15068 20383
rect 15016 20340 15068 20349
rect 15660 20383 15712 20392
rect 15660 20349 15669 20383
rect 15669 20349 15703 20383
rect 15703 20349 15712 20383
rect 15660 20340 15712 20349
rect 16764 20383 16816 20392
rect 16764 20349 16773 20383
rect 16773 20349 16807 20383
rect 16807 20349 16816 20383
rect 16764 20340 16816 20349
rect 17040 20340 17092 20392
rect 16396 20272 16448 20324
rect 7012 20204 7064 20256
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 7380 20247 7432 20256
rect 7380 20213 7389 20247
rect 7389 20213 7423 20247
rect 7423 20213 7432 20247
rect 7380 20204 7432 20213
rect 7472 20204 7524 20256
rect 9772 20204 9824 20256
rect 12900 20204 12952 20256
rect 13268 20247 13320 20256
rect 13268 20213 13277 20247
rect 13277 20213 13311 20247
rect 13311 20213 13320 20247
rect 13268 20204 13320 20213
rect 14556 20204 14608 20256
rect 15200 20204 15252 20256
rect 16028 20204 16080 20256
rect 16120 20247 16172 20256
rect 16120 20213 16129 20247
rect 16129 20213 16163 20247
rect 16163 20213 16172 20247
rect 16120 20204 16172 20213
rect 16304 20247 16356 20256
rect 16304 20213 16313 20247
rect 16313 20213 16347 20247
rect 16347 20213 16356 20247
rect 16304 20204 16356 20213
rect 18144 20272 18196 20324
rect 19340 20272 19392 20324
rect 20444 20408 20496 20460
rect 21456 20408 21508 20460
rect 22376 20408 22428 20460
rect 22836 20451 22888 20460
rect 22836 20417 22845 20451
rect 22845 20417 22879 20451
rect 22879 20417 22888 20451
rect 22836 20408 22888 20417
rect 22928 20408 22980 20460
rect 23664 20408 23716 20460
rect 24216 20408 24268 20460
rect 21824 20340 21876 20392
rect 23572 20340 23624 20392
rect 24308 20340 24360 20392
rect 24768 20340 24820 20392
rect 21456 20272 21508 20324
rect 16948 20204 17000 20256
rect 17224 20204 17276 20256
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 21088 20247 21140 20256
rect 21088 20213 21097 20247
rect 21097 20213 21131 20247
rect 21131 20213 21140 20247
rect 21088 20204 21140 20213
rect 22008 20272 22060 20324
rect 25688 20451 25740 20460
rect 25688 20417 25697 20451
rect 25697 20417 25731 20451
rect 25731 20417 25740 20451
rect 25688 20408 25740 20417
rect 25780 20451 25832 20460
rect 25780 20417 25789 20451
rect 25789 20417 25823 20451
rect 25823 20417 25832 20451
rect 25780 20408 25832 20417
rect 25964 20408 26016 20460
rect 26332 20451 26384 20460
rect 26332 20417 26349 20451
rect 26349 20417 26384 20451
rect 26332 20408 26384 20417
rect 26424 20451 26476 20460
rect 26424 20417 26433 20451
rect 26433 20417 26467 20451
rect 26467 20417 26476 20451
rect 26424 20408 26476 20417
rect 26516 20451 26568 20460
rect 26516 20417 26525 20451
rect 26525 20417 26559 20451
rect 26559 20417 26568 20451
rect 26516 20408 26568 20417
rect 26792 20476 26844 20528
rect 28172 20544 28224 20596
rect 33876 20544 33928 20596
rect 27068 20408 27120 20460
rect 27252 20451 27304 20460
rect 27252 20417 27261 20451
rect 27261 20417 27295 20451
rect 27295 20417 27304 20451
rect 27252 20408 27304 20417
rect 26516 20272 26568 20324
rect 29368 20476 29420 20528
rect 32588 20476 32640 20528
rect 27712 20204 27764 20256
rect 30288 20451 30340 20460
rect 30288 20417 30297 20451
rect 30297 20417 30331 20451
rect 30331 20417 30340 20451
rect 30288 20408 30340 20417
rect 30656 20408 30708 20460
rect 30748 20408 30800 20460
rect 31116 20451 31168 20460
rect 31116 20417 31125 20451
rect 31125 20417 31159 20451
rect 31159 20417 31168 20451
rect 31116 20408 31168 20417
rect 31300 20451 31352 20460
rect 31300 20417 31309 20451
rect 31309 20417 31343 20451
rect 31343 20417 31352 20451
rect 31300 20408 31352 20417
rect 31392 20408 31444 20460
rect 35532 20408 35584 20460
rect 28448 20340 28500 20392
rect 28816 20340 28868 20392
rect 34612 20383 34664 20392
rect 34612 20349 34621 20383
rect 34621 20349 34655 20383
rect 34655 20349 34664 20383
rect 34612 20340 34664 20349
rect 34796 20272 34848 20324
rect 29552 20204 29604 20256
rect 30472 20247 30524 20256
rect 30472 20213 30481 20247
rect 30481 20213 30515 20247
rect 30515 20213 30524 20247
rect 30472 20204 30524 20213
rect 31208 20204 31260 20256
rect 33968 20204 34020 20256
rect 34520 20247 34572 20256
rect 34520 20213 34529 20247
rect 34529 20213 34563 20247
rect 34563 20213 34572 20247
rect 34520 20204 34572 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4896 20000 4948 20052
rect 6368 20000 6420 20052
rect 6644 20000 6696 20052
rect 7380 20000 7432 20052
rect 8392 20043 8444 20052
rect 8392 20009 8401 20043
rect 8401 20009 8435 20043
rect 8435 20009 8444 20043
rect 8392 20000 8444 20009
rect 8484 20000 8536 20052
rect 9128 20000 9180 20052
rect 9588 20000 9640 20052
rect 9956 20000 10008 20052
rect 11060 20000 11112 20052
rect 11796 20000 11848 20052
rect 12532 20000 12584 20052
rect 13636 20043 13688 20052
rect 13636 20009 13645 20043
rect 13645 20009 13679 20043
rect 13679 20009 13688 20043
rect 13636 20000 13688 20009
rect 14280 20000 14332 20052
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 3700 19796 3752 19848
rect 4436 19864 4488 19916
rect 5080 19907 5132 19916
rect 5080 19873 5089 19907
rect 5089 19873 5123 19907
rect 5123 19873 5132 19907
rect 5080 19864 5132 19873
rect 8208 19932 8260 19984
rect 4252 19796 4304 19848
rect 6368 19864 6420 19916
rect 6920 19864 6972 19916
rect 7288 19864 7340 19916
rect 8852 19864 8904 19916
rect 12256 19864 12308 19916
rect 12532 19864 12584 19916
rect 6184 19839 6236 19848
rect 6184 19805 6193 19839
rect 6193 19805 6227 19839
rect 6227 19805 6236 19839
rect 6184 19796 6236 19805
rect 8484 19839 8536 19848
rect 8484 19805 8493 19839
rect 8493 19805 8527 19839
rect 8527 19805 8536 19839
rect 8484 19796 8536 19805
rect 1676 19771 1728 19780
rect 1676 19737 1685 19771
rect 1685 19737 1719 19771
rect 1719 19737 1728 19771
rect 1676 19728 1728 19737
rect 2964 19728 3016 19780
rect 3424 19660 3476 19712
rect 4344 19728 4396 19780
rect 5540 19703 5592 19712
rect 5540 19669 5549 19703
rect 5549 19669 5583 19703
rect 5583 19669 5592 19703
rect 5540 19660 5592 19669
rect 6828 19728 6880 19780
rect 6552 19660 6604 19712
rect 7104 19660 7156 19712
rect 7288 19660 7340 19712
rect 8944 19796 8996 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 8852 19728 8904 19780
rect 9312 19796 9364 19848
rect 15016 19864 15068 19916
rect 15936 20043 15988 20052
rect 15936 20009 15945 20043
rect 15945 20009 15979 20043
rect 15979 20009 15988 20043
rect 15936 20000 15988 20009
rect 16580 20043 16632 20052
rect 16580 20009 16589 20043
rect 16589 20009 16623 20043
rect 16623 20009 16632 20043
rect 16580 20000 16632 20009
rect 17408 20000 17460 20052
rect 20260 20000 20312 20052
rect 22100 20000 22152 20052
rect 26056 20043 26108 20052
rect 26056 20009 26065 20043
rect 26065 20009 26099 20043
rect 26099 20009 26108 20043
rect 26056 20000 26108 20009
rect 27252 20000 27304 20052
rect 28816 20000 28868 20052
rect 29552 20043 29604 20052
rect 29552 20009 29561 20043
rect 29561 20009 29595 20043
rect 29595 20009 29604 20043
rect 29552 20000 29604 20009
rect 31392 20000 31444 20052
rect 33692 20000 33744 20052
rect 15660 19932 15712 19984
rect 19984 19932 20036 19984
rect 21548 19932 21600 19984
rect 26424 19932 26476 19984
rect 31024 19932 31076 19984
rect 9404 19728 9456 19780
rect 10232 19728 10284 19780
rect 8944 19703 8996 19712
rect 8944 19669 8953 19703
rect 8953 19669 8987 19703
rect 8987 19669 8996 19703
rect 8944 19660 8996 19669
rect 9220 19660 9272 19712
rect 10048 19660 10100 19712
rect 14556 19728 14608 19780
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 15936 19796 15988 19848
rect 16396 19839 16448 19848
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 17132 19796 17184 19848
rect 17868 19864 17920 19916
rect 18144 19864 18196 19916
rect 19064 19864 19116 19916
rect 20812 19864 20864 19916
rect 20904 19864 20956 19916
rect 16764 19728 16816 19780
rect 17040 19771 17092 19780
rect 17040 19737 17049 19771
rect 17049 19737 17083 19771
rect 17083 19737 17092 19771
rect 17040 19728 17092 19737
rect 17684 19728 17736 19780
rect 18328 19796 18380 19848
rect 18512 19796 18564 19848
rect 20996 19796 21048 19848
rect 22652 19864 22704 19916
rect 12072 19660 12124 19712
rect 14372 19660 14424 19712
rect 15108 19660 15160 19712
rect 16028 19660 16080 19712
rect 16672 19660 16724 19712
rect 17132 19660 17184 19712
rect 18972 19728 19024 19780
rect 19248 19771 19300 19780
rect 19248 19737 19257 19771
rect 19257 19737 19291 19771
rect 19291 19737 19300 19771
rect 19248 19728 19300 19737
rect 19708 19728 19760 19780
rect 20260 19728 20312 19780
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 26516 19864 26568 19916
rect 21456 19796 21508 19805
rect 25964 19796 26016 19848
rect 27804 19839 27856 19848
rect 27804 19805 27813 19839
rect 27813 19805 27847 19839
rect 27847 19805 27856 19839
rect 27804 19796 27856 19805
rect 29368 19864 29420 19916
rect 29736 19907 29788 19916
rect 29736 19873 29745 19907
rect 29745 19873 29779 19907
rect 29779 19873 29788 19907
rect 29736 19864 29788 19873
rect 33968 19907 34020 19916
rect 33968 19873 33977 19907
rect 33977 19873 34011 19907
rect 34011 19873 34020 19907
rect 33968 19864 34020 19873
rect 35256 19864 35308 19916
rect 35532 19864 35584 19916
rect 28172 19839 28224 19848
rect 28172 19805 28181 19839
rect 28181 19805 28215 19839
rect 28215 19805 28224 19839
rect 28172 19796 28224 19805
rect 29276 19796 29328 19848
rect 34152 19839 34204 19848
rect 34152 19805 34161 19839
rect 34161 19805 34195 19839
rect 34195 19805 34204 19839
rect 34152 19796 34204 19805
rect 23480 19728 23532 19780
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 18696 19660 18748 19712
rect 23388 19660 23440 19712
rect 26792 19660 26844 19712
rect 28540 19728 28592 19780
rect 33968 19728 34020 19780
rect 34152 19660 34204 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 1676 19456 1728 19508
rect 2136 19456 2188 19508
rect 2596 19456 2648 19508
rect 3516 19456 3568 19508
rect 4068 19456 4120 19508
rect 4344 19456 4396 19508
rect 4436 19456 4488 19508
rect 4896 19456 4948 19508
rect 7288 19456 7340 19508
rect 7564 19456 7616 19508
rect 3332 19388 3384 19440
rect 4712 19388 4764 19440
rect 5816 19431 5868 19440
rect 5816 19397 5825 19431
rect 5825 19397 5859 19431
rect 5859 19397 5868 19431
rect 5816 19388 5868 19397
rect 3424 19363 3476 19372
rect 3424 19329 3433 19363
rect 3433 19329 3467 19363
rect 3467 19329 3476 19363
rect 3424 19320 3476 19329
rect 3608 19363 3660 19372
rect 3608 19329 3617 19363
rect 3617 19329 3651 19363
rect 3651 19329 3660 19363
rect 3608 19320 3660 19329
rect 3884 19363 3936 19372
rect 3884 19329 3893 19363
rect 3893 19329 3927 19363
rect 3927 19329 3936 19363
rect 3884 19320 3936 19329
rect 4252 19320 4304 19372
rect 4988 19320 5040 19372
rect 5448 19363 5500 19372
rect 5448 19329 5457 19363
rect 5457 19329 5491 19363
rect 5491 19329 5500 19363
rect 5448 19320 5500 19329
rect 6920 19388 6972 19440
rect 7932 19388 7984 19440
rect 2596 19295 2648 19304
rect 2596 19261 2605 19295
rect 2605 19261 2639 19295
rect 2639 19261 2648 19295
rect 2596 19252 2648 19261
rect 5724 19252 5776 19304
rect 6736 19252 6788 19304
rect 8392 19388 8444 19440
rect 8208 19363 8260 19372
rect 8208 19329 8217 19363
rect 8217 19329 8251 19363
rect 8251 19329 8260 19363
rect 8208 19320 8260 19329
rect 8300 19363 8352 19372
rect 8300 19329 8310 19363
rect 8310 19329 8344 19363
rect 8344 19329 8352 19363
rect 8300 19320 8352 19329
rect 10232 19499 10284 19508
rect 10232 19465 10241 19499
rect 10241 19465 10275 19499
rect 10275 19465 10284 19499
rect 10232 19456 10284 19465
rect 8300 19184 8352 19236
rect 9404 19363 9456 19372
rect 9404 19329 9413 19363
rect 9413 19329 9447 19363
rect 9447 19329 9456 19363
rect 9404 19320 9456 19329
rect 9680 19320 9732 19372
rect 9220 19252 9272 19304
rect 9772 19295 9824 19304
rect 9772 19261 9781 19295
rect 9781 19261 9815 19295
rect 9815 19261 9824 19295
rect 9772 19252 9824 19261
rect 10324 19388 10376 19440
rect 10048 19363 10100 19372
rect 10048 19329 10057 19363
rect 10057 19329 10091 19363
rect 10091 19329 10100 19363
rect 12440 19456 12492 19508
rect 10784 19388 10836 19440
rect 14188 19456 14240 19508
rect 14372 19456 14424 19508
rect 16396 19456 16448 19508
rect 18420 19456 18472 19508
rect 18788 19456 18840 19508
rect 19340 19456 19392 19508
rect 19892 19456 19944 19508
rect 19984 19456 20036 19508
rect 22560 19456 22612 19508
rect 23204 19456 23256 19508
rect 24676 19456 24728 19508
rect 13544 19388 13596 19440
rect 13636 19431 13688 19440
rect 13636 19397 13645 19431
rect 13645 19397 13679 19431
rect 13679 19397 13688 19431
rect 13636 19388 13688 19397
rect 13912 19388 13964 19440
rect 10048 19320 10100 19329
rect 11796 19320 11848 19372
rect 12624 19320 12676 19372
rect 13176 19363 13228 19372
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 13268 19320 13320 19372
rect 10692 19252 10744 19304
rect 10876 19295 10928 19304
rect 10876 19261 10885 19295
rect 10885 19261 10919 19295
rect 10919 19261 10928 19295
rect 10876 19252 10928 19261
rect 12808 19252 12860 19304
rect 8760 19184 8812 19236
rect 4620 19116 4672 19168
rect 7196 19116 7248 19168
rect 8668 19116 8720 19168
rect 11888 19184 11940 19236
rect 13452 19184 13504 19236
rect 13820 19184 13872 19236
rect 14280 19388 14332 19440
rect 14096 19363 14148 19372
rect 14096 19329 14105 19363
rect 14105 19329 14139 19363
rect 14139 19329 14148 19363
rect 14096 19320 14148 19329
rect 14556 19320 14608 19372
rect 15200 19320 15252 19372
rect 16212 19388 16264 19440
rect 15568 19320 15620 19372
rect 14280 19295 14332 19304
rect 14280 19261 14289 19295
rect 14289 19261 14323 19295
rect 14323 19261 14332 19295
rect 14280 19252 14332 19261
rect 16764 19252 16816 19304
rect 18604 19388 18656 19440
rect 17132 19363 17184 19372
rect 17132 19329 17141 19363
rect 17141 19329 17175 19363
rect 17175 19329 17184 19363
rect 17132 19320 17184 19329
rect 17684 19320 17736 19372
rect 18604 19252 18656 19304
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19064 19320 19116 19372
rect 20628 19388 20680 19440
rect 19708 19320 19760 19372
rect 19340 19252 19392 19304
rect 19984 19320 20036 19372
rect 20260 19363 20312 19372
rect 20260 19329 20269 19363
rect 20269 19329 20303 19363
rect 20303 19329 20312 19363
rect 20260 19320 20312 19329
rect 20904 19320 20956 19372
rect 22652 19363 22704 19372
rect 22652 19329 22661 19363
rect 22661 19329 22695 19363
rect 22695 19329 22704 19363
rect 22652 19320 22704 19329
rect 22836 19388 22888 19440
rect 23296 19388 23348 19440
rect 24768 19388 24820 19440
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 24400 19320 24452 19372
rect 19248 19184 19300 19236
rect 12348 19116 12400 19168
rect 12716 19116 12768 19168
rect 12992 19159 13044 19168
rect 12992 19125 13001 19159
rect 13001 19125 13035 19159
rect 13035 19125 13044 19159
rect 12992 19116 13044 19125
rect 13268 19116 13320 19168
rect 16396 19116 16448 19168
rect 16764 19116 16816 19168
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 21364 19184 21416 19236
rect 23296 19295 23348 19304
rect 23296 19261 23305 19295
rect 23305 19261 23339 19295
rect 23339 19261 23348 19295
rect 23296 19252 23348 19261
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 25228 19363 25280 19372
rect 25228 19329 25237 19363
rect 25237 19329 25271 19363
rect 25271 19329 25280 19363
rect 25228 19320 25280 19329
rect 30380 19456 30432 19508
rect 33968 19456 34020 19508
rect 27804 19388 27856 19440
rect 27896 19363 27948 19372
rect 27896 19329 27905 19363
rect 27905 19329 27939 19363
rect 27939 19329 27948 19363
rect 27896 19320 27948 19329
rect 29644 19388 29696 19440
rect 28264 19363 28316 19372
rect 28264 19329 28273 19363
rect 28273 19329 28307 19363
rect 28307 19329 28316 19363
rect 28264 19320 28316 19329
rect 29000 19320 29052 19372
rect 32772 19363 32824 19372
rect 32772 19329 32781 19363
rect 32781 19329 32815 19363
rect 32815 19329 32824 19363
rect 32772 19320 32824 19329
rect 34428 19320 34480 19372
rect 29092 19252 29144 19304
rect 29828 19252 29880 19304
rect 30196 19252 30248 19304
rect 32864 19295 32916 19304
rect 32864 19261 32873 19295
rect 32873 19261 32907 19295
rect 32907 19261 32916 19295
rect 32864 19252 32916 19261
rect 32956 19252 33008 19304
rect 26700 19184 26752 19236
rect 30472 19184 30524 19236
rect 24308 19116 24360 19168
rect 24400 19116 24452 19168
rect 25780 19116 25832 19168
rect 27988 19116 28040 19168
rect 28172 19116 28224 19168
rect 28540 19159 28592 19168
rect 28540 19125 28549 19159
rect 28549 19125 28583 19159
rect 28583 19125 28592 19159
rect 28540 19116 28592 19125
rect 30012 19116 30064 19168
rect 30564 19116 30616 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3516 18912 3568 18964
rect 3884 18912 3936 18964
rect 5448 18912 5500 18964
rect 6736 18955 6788 18964
rect 6736 18921 6745 18955
rect 6745 18921 6779 18955
rect 6779 18921 6788 18955
rect 6736 18912 6788 18921
rect 4620 18844 4672 18896
rect 6644 18844 6696 18896
rect 8760 18912 8812 18964
rect 9404 18912 9456 18964
rect 9864 18912 9916 18964
rect 10692 18955 10744 18964
rect 10692 18921 10701 18955
rect 10701 18921 10735 18955
rect 10735 18921 10744 18955
rect 10692 18912 10744 18921
rect 6920 18844 6972 18896
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 2780 18708 2832 18760
rect 4988 18776 5040 18828
rect 5448 18776 5500 18828
rect 7012 18776 7064 18828
rect 4436 18751 4488 18760
rect 4436 18717 4445 18751
rect 4445 18717 4479 18751
rect 4479 18717 4488 18751
rect 4436 18708 4488 18717
rect 1676 18683 1728 18692
rect 1676 18649 1685 18683
rect 1685 18649 1719 18683
rect 1719 18649 1728 18683
rect 1676 18640 1728 18649
rect 4896 18708 4948 18760
rect 5356 18640 5408 18692
rect 8024 18708 8076 18760
rect 8392 18776 8444 18828
rect 9220 18776 9272 18828
rect 9588 18776 9640 18828
rect 10692 18776 10744 18828
rect 11152 18776 11204 18828
rect 12072 18912 12124 18964
rect 8760 18708 8812 18760
rect 11060 18708 11112 18760
rect 12440 18844 12492 18896
rect 12716 18844 12768 18896
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 11888 18708 11940 18760
rect 12072 18751 12124 18760
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 8392 18572 8444 18624
rect 8852 18572 8904 18624
rect 9220 18683 9272 18692
rect 9220 18649 9229 18683
rect 9229 18649 9263 18683
rect 9263 18649 9272 18683
rect 9220 18640 9272 18649
rect 9772 18640 9824 18692
rect 10508 18640 10560 18692
rect 11244 18640 11296 18692
rect 12256 18683 12308 18692
rect 12256 18649 12265 18683
rect 12265 18649 12299 18683
rect 12299 18649 12308 18683
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 13452 18751 13504 18760
rect 13452 18717 13461 18751
rect 13461 18717 13495 18751
rect 13495 18717 13504 18751
rect 13452 18708 13504 18717
rect 13636 18912 13688 18964
rect 14096 18912 14148 18964
rect 15384 18912 15436 18964
rect 16764 18912 16816 18964
rect 20904 18912 20956 18964
rect 21824 18912 21876 18964
rect 23112 18955 23164 18964
rect 23112 18921 23121 18955
rect 23121 18921 23155 18955
rect 23155 18921 23164 18955
rect 23112 18912 23164 18921
rect 24308 18912 24360 18964
rect 28724 18912 28776 18964
rect 29184 18912 29236 18964
rect 30196 18955 30248 18964
rect 30196 18921 30205 18955
rect 30205 18921 30239 18955
rect 30239 18921 30248 18955
rect 30196 18912 30248 18921
rect 30656 18955 30708 18964
rect 30656 18921 30665 18955
rect 30665 18921 30699 18955
rect 30699 18921 30708 18955
rect 30656 18912 30708 18921
rect 33692 18912 33744 18964
rect 16672 18844 16724 18896
rect 15936 18776 15988 18828
rect 16580 18776 16632 18828
rect 21272 18776 21324 18828
rect 22008 18776 22060 18828
rect 12256 18640 12308 18649
rect 13176 18640 13228 18692
rect 9864 18572 9916 18624
rect 10876 18572 10928 18624
rect 12348 18572 12400 18624
rect 15752 18751 15804 18760
rect 15752 18717 15758 18751
rect 15758 18717 15792 18751
rect 15792 18717 15804 18751
rect 15752 18708 15804 18717
rect 16120 18751 16172 18760
rect 16120 18717 16129 18751
rect 16129 18717 16163 18751
rect 16163 18717 16172 18751
rect 16120 18708 16172 18717
rect 16672 18708 16724 18760
rect 17040 18751 17092 18760
rect 17040 18717 17049 18751
rect 17049 18717 17083 18751
rect 17083 18717 17092 18751
rect 17040 18708 17092 18717
rect 14188 18640 14240 18692
rect 14556 18640 14608 18692
rect 17684 18640 17736 18692
rect 18144 18708 18196 18760
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 21548 18751 21600 18760
rect 21548 18717 21557 18751
rect 21557 18717 21591 18751
rect 21591 18717 21600 18751
rect 21548 18708 21600 18717
rect 21916 18751 21968 18760
rect 21916 18717 21925 18751
rect 21925 18717 21959 18751
rect 21959 18717 21968 18751
rect 21916 18708 21968 18717
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 18604 18640 18656 18692
rect 23296 18751 23348 18760
rect 23296 18717 23305 18751
rect 23305 18717 23339 18751
rect 23339 18717 23348 18751
rect 23296 18708 23348 18717
rect 23480 18751 23532 18760
rect 23480 18717 23489 18751
rect 23489 18717 23523 18751
rect 23523 18717 23532 18751
rect 23480 18708 23532 18717
rect 23664 18640 23716 18692
rect 16212 18572 16264 18624
rect 16856 18615 16908 18624
rect 16856 18581 16865 18615
rect 16865 18581 16899 18615
rect 16899 18581 16908 18615
rect 16856 18572 16908 18581
rect 21272 18572 21324 18624
rect 23296 18572 23348 18624
rect 24308 18708 24360 18760
rect 24216 18640 24268 18692
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 25228 18708 25280 18760
rect 25596 18640 25648 18692
rect 25872 18751 25924 18760
rect 25872 18717 25881 18751
rect 25881 18717 25915 18751
rect 25915 18717 25924 18751
rect 25872 18708 25924 18717
rect 26056 18776 26108 18828
rect 26700 18751 26752 18760
rect 26700 18717 26709 18751
rect 26709 18717 26743 18751
rect 26743 18717 26752 18751
rect 26700 18708 26752 18717
rect 27068 18708 27120 18760
rect 27528 18751 27580 18760
rect 27528 18717 27537 18751
rect 27537 18717 27571 18751
rect 27571 18717 27580 18751
rect 27528 18708 27580 18717
rect 27620 18751 27672 18760
rect 27620 18717 27630 18751
rect 27630 18717 27664 18751
rect 27664 18717 27672 18751
rect 27620 18708 27672 18717
rect 28172 18844 28224 18896
rect 28908 18844 28960 18896
rect 27988 18751 28040 18760
rect 27988 18717 28002 18751
rect 28002 18717 28036 18751
rect 28036 18717 28040 18751
rect 27988 18708 28040 18717
rect 29552 18751 29604 18760
rect 29552 18717 29561 18751
rect 29561 18717 29595 18751
rect 29595 18717 29604 18751
rect 29552 18708 29604 18717
rect 29644 18751 29696 18760
rect 29644 18717 29654 18751
rect 29654 18717 29688 18751
rect 29688 18717 29696 18751
rect 29644 18708 29696 18717
rect 29828 18751 29880 18760
rect 29828 18717 29837 18751
rect 29837 18717 29871 18751
rect 29871 18717 29880 18751
rect 29828 18708 29880 18717
rect 30748 18708 30800 18760
rect 26056 18640 26108 18692
rect 27436 18640 27488 18692
rect 24952 18572 25004 18624
rect 25504 18615 25556 18624
rect 25504 18581 25513 18615
rect 25513 18581 25547 18615
rect 25547 18581 25556 18615
rect 25504 18572 25556 18581
rect 25872 18572 25924 18624
rect 28264 18640 28316 18692
rect 28908 18572 28960 18624
rect 30472 18640 30524 18692
rect 33600 18844 33652 18896
rect 32864 18776 32916 18828
rect 33232 18708 33284 18760
rect 35348 18708 35400 18760
rect 33692 18640 33744 18692
rect 30104 18572 30156 18624
rect 33324 18572 33376 18624
rect 35348 18572 35400 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 1676 18368 1728 18420
rect 5448 18368 5500 18420
rect 3516 18275 3568 18284
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 7564 18368 7616 18420
rect 7748 18411 7800 18420
rect 7748 18377 7757 18411
rect 7757 18377 7791 18411
rect 7791 18377 7800 18411
rect 7748 18368 7800 18377
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 8484 18368 8536 18420
rect 9220 18368 9272 18420
rect 10508 18368 10560 18420
rect 7104 18300 7156 18352
rect 2504 18207 2556 18216
rect 2504 18173 2513 18207
rect 2513 18173 2547 18207
rect 2547 18173 2556 18207
rect 2504 18164 2556 18173
rect 2596 18207 2648 18216
rect 2596 18173 2605 18207
rect 2605 18173 2639 18207
rect 2639 18173 2648 18207
rect 2596 18164 2648 18173
rect 5724 18164 5776 18216
rect 8392 18275 8444 18284
rect 8392 18241 8401 18275
rect 8401 18241 8435 18275
rect 8435 18241 8444 18275
rect 8392 18232 8444 18241
rect 8576 18232 8628 18284
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 9496 18343 9548 18352
rect 9496 18309 9505 18343
rect 9505 18309 9539 18343
rect 9539 18309 9548 18343
rect 9496 18300 9548 18309
rect 10048 18343 10100 18352
rect 10048 18309 10057 18343
rect 10057 18309 10091 18343
rect 10091 18309 10100 18343
rect 10048 18300 10100 18309
rect 10140 18300 10192 18352
rect 11888 18368 11940 18420
rect 8944 18232 8996 18284
rect 8852 18164 8904 18216
rect 9864 18164 9916 18216
rect 10232 18164 10284 18216
rect 10692 18232 10744 18284
rect 11428 18300 11480 18352
rect 10968 18232 11020 18284
rect 11888 18232 11940 18284
rect 12072 18232 12124 18284
rect 12164 18275 12216 18284
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12808 18368 12860 18420
rect 13084 18368 13136 18420
rect 13820 18411 13872 18420
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 15752 18368 15804 18420
rect 21456 18368 21508 18420
rect 12164 18232 12216 18241
rect 12716 18275 12768 18284
rect 12716 18241 12725 18275
rect 12725 18241 12759 18275
rect 12759 18241 12768 18275
rect 12716 18232 12768 18241
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 16856 18300 16908 18352
rect 22008 18300 22060 18352
rect 23020 18411 23072 18420
rect 23020 18377 23029 18411
rect 23029 18377 23063 18411
rect 23063 18377 23072 18411
rect 23020 18368 23072 18377
rect 24584 18368 24636 18420
rect 25780 18368 25832 18420
rect 26700 18368 26752 18420
rect 27620 18368 27672 18420
rect 27896 18368 27948 18420
rect 30748 18368 30800 18420
rect 31576 18368 31628 18420
rect 31852 18368 31904 18420
rect 12992 18232 13044 18241
rect 9128 18096 9180 18148
rect 7380 18071 7432 18080
rect 7380 18037 7389 18071
rect 7389 18037 7423 18071
rect 7423 18037 7432 18071
rect 7380 18028 7432 18037
rect 8392 18028 8444 18080
rect 9220 18028 9272 18080
rect 9680 18028 9732 18080
rect 10048 18028 10100 18080
rect 10692 18028 10744 18080
rect 11152 18164 11204 18216
rect 12256 18207 12308 18216
rect 12256 18173 12265 18207
rect 12265 18173 12299 18207
rect 12299 18173 12308 18207
rect 12256 18164 12308 18173
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 13544 18232 13596 18284
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 21364 18275 21416 18284
rect 21364 18241 21373 18275
rect 21373 18241 21407 18275
rect 21407 18241 21416 18275
rect 21364 18232 21416 18241
rect 23480 18300 23532 18352
rect 24216 18300 24268 18352
rect 27068 18300 27120 18352
rect 23664 18275 23716 18284
rect 23664 18241 23673 18275
rect 23673 18241 23707 18275
rect 23707 18241 23716 18275
rect 23664 18232 23716 18241
rect 23756 18232 23808 18284
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 24124 18232 24176 18284
rect 13176 18164 13228 18173
rect 15660 18164 15712 18216
rect 21732 18164 21784 18216
rect 25412 18275 25464 18284
rect 25412 18241 25421 18275
rect 25421 18241 25455 18275
rect 25455 18241 25464 18275
rect 25412 18232 25464 18241
rect 24860 18164 24912 18216
rect 25044 18164 25096 18216
rect 25596 18232 25648 18284
rect 26056 18232 26108 18284
rect 26148 18275 26200 18284
rect 26148 18241 26157 18275
rect 26157 18241 26191 18275
rect 26191 18241 26200 18275
rect 26148 18232 26200 18241
rect 28172 18300 28224 18352
rect 27344 18232 27396 18284
rect 27528 18275 27580 18284
rect 27528 18241 27537 18275
rect 27537 18241 27571 18275
rect 27571 18241 27580 18275
rect 27528 18232 27580 18241
rect 27804 18232 27856 18284
rect 28172 18164 28224 18216
rect 12532 18096 12584 18148
rect 13084 18096 13136 18148
rect 18052 18096 18104 18148
rect 21180 18096 21232 18148
rect 24676 18096 24728 18148
rect 11152 18028 11204 18080
rect 11336 18028 11388 18080
rect 20628 18071 20680 18080
rect 20628 18037 20637 18071
rect 20637 18037 20671 18071
rect 20671 18037 20680 18071
rect 20628 18028 20680 18037
rect 22008 18028 22060 18080
rect 24400 18028 24452 18080
rect 25412 18028 25464 18080
rect 25688 18096 25740 18148
rect 29000 18232 29052 18284
rect 29644 18232 29696 18284
rect 33600 18300 33652 18352
rect 33692 18343 33744 18352
rect 33692 18309 33701 18343
rect 33701 18309 33735 18343
rect 33735 18309 33744 18343
rect 33692 18300 33744 18309
rect 32772 18275 32824 18284
rect 32772 18241 32781 18275
rect 32781 18241 32815 18275
rect 32815 18241 32824 18275
rect 32772 18232 32824 18241
rect 32956 18275 33008 18284
rect 32956 18241 32965 18275
rect 32965 18241 32999 18275
rect 32999 18241 33008 18275
rect 32956 18232 33008 18241
rect 33324 18232 33376 18284
rect 33784 18275 33836 18284
rect 33784 18241 33793 18275
rect 33793 18241 33827 18275
rect 33827 18241 33836 18275
rect 33784 18232 33836 18241
rect 35256 18411 35308 18420
rect 35256 18377 35265 18411
rect 35265 18377 35299 18411
rect 35299 18377 35308 18411
rect 35256 18368 35308 18377
rect 34336 18300 34388 18352
rect 35348 18343 35400 18352
rect 35348 18309 35357 18343
rect 35357 18309 35391 18343
rect 35391 18309 35400 18343
rect 35348 18300 35400 18309
rect 31944 18096 31996 18148
rect 35440 18232 35492 18284
rect 29828 18028 29880 18080
rect 31208 18028 31260 18080
rect 34612 18028 34664 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2320 17620 2372 17672
rect 3332 17824 3384 17876
rect 4620 17824 4672 17876
rect 4344 17688 4396 17740
rect 5816 17824 5868 17876
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 11244 17824 11296 17876
rect 11428 17824 11480 17876
rect 12164 17824 12216 17876
rect 12440 17867 12492 17876
rect 12440 17833 12449 17867
rect 12449 17833 12483 17867
rect 12483 17833 12492 17867
rect 12440 17824 12492 17833
rect 14004 17824 14056 17876
rect 14648 17824 14700 17876
rect 15108 17824 15160 17876
rect 18604 17824 18656 17876
rect 18880 17824 18932 17876
rect 20720 17824 20772 17876
rect 21640 17824 21692 17876
rect 22376 17824 22428 17876
rect 23664 17867 23716 17876
rect 23664 17833 23673 17867
rect 23673 17833 23707 17867
rect 23707 17833 23716 17867
rect 23664 17824 23716 17833
rect 24676 17824 24728 17876
rect 24952 17824 25004 17876
rect 25780 17824 25832 17876
rect 28908 17824 28960 17876
rect 31484 17824 31536 17876
rect 31668 17824 31720 17876
rect 34336 17867 34388 17876
rect 34336 17833 34345 17867
rect 34345 17833 34379 17867
rect 34379 17833 34388 17867
rect 34336 17824 34388 17833
rect 34520 17867 34572 17876
rect 34520 17833 34529 17867
rect 34529 17833 34563 17867
rect 34563 17833 34572 17867
rect 34520 17824 34572 17833
rect 9036 17756 9088 17808
rect 10232 17756 10284 17808
rect 10692 17756 10744 17808
rect 3424 17620 3476 17672
rect 3792 17620 3844 17672
rect 3056 17552 3108 17604
rect 3240 17552 3292 17604
rect 3608 17552 3660 17604
rect 4160 17595 4212 17604
rect 4160 17561 4169 17595
rect 4169 17561 4203 17595
rect 4203 17561 4212 17595
rect 4160 17552 4212 17561
rect 4528 17620 4580 17672
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 8576 17688 8628 17740
rect 9680 17688 9732 17740
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 4896 17663 4948 17672
rect 4896 17629 4905 17663
rect 4905 17629 4939 17663
rect 4939 17629 4948 17663
rect 4896 17620 4948 17629
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 6644 17620 6696 17672
rect 7932 17620 7984 17672
rect 4804 17484 4856 17536
rect 5540 17552 5592 17604
rect 5632 17595 5684 17604
rect 5632 17561 5641 17595
rect 5641 17561 5675 17595
rect 5675 17561 5684 17595
rect 5632 17552 5684 17561
rect 7748 17552 7800 17604
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 9036 17552 9088 17604
rect 9496 17552 9548 17604
rect 5908 17484 5960 17536
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 7564 17484 7616 17536
rect 9312 17484 9364 17536
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 10416 17688 10468 17740
rect 10692 17620 10744 17672
rect 10048 17484 10100 17536
rect 10140 17484 10192 17536
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 10692 17484 10744 17536
rect 11428 17620 11480 17672
rect 11520 17620 11572 17672
rect 11888 17663 11940 17672
rect 11888 17629 11892 17663
rect 11892 17629 11926 17663
rect 11926 17629 11940 17663
rect 11888 17620 11940 17629
rect 11152 17595 11204 17604
rect 11152 17561 11161 17595
rect 11161 17561 11195 17595
rect 11195 17561 11204 17595
rect 11152 17552 11204 17561
rect 11796 17552 11848 17604
rect 14740 17756 14792 17808
rect 14924 17756 14976 17808
rect 21824 17756 21876 17808
rect 23020 17756 23072 17808
rect 24492 17756 24544 17808
rect 25136 17756 25188 17808
rect 12164 17663 12216 17672
rect 12164 17629 12209 17663
rect 12209 17629 12216 17663
rect 12164 17620 12216 17629
rect 12440 17620 12492 17672
rect 12624 17663 12676 17672
rect 12624 17629 12633 17663
rect 12633 17629 12667 17663
rect 12667 17629 12676 17663
rect 12624 17620 12676 17629
rect 12992 17620 13044 17672
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 15016 17620 15068 17672
rect 15384 17620 15436 17672
rect 15752 17663 15804 17672
rect 15752 17629 15761 17663
rect 15761 17629 15795 17663
rect 15795 17629 15804 17663
rect 15752 17620 15804 17629
rect 17592 17688 17644 17740
rect 16028 17663 16080 17672
rect 16028 17629 16037 17663
rect 16037 17629 16071 17663
rect 16071 17629 16080 17663
rect 16028 17620 16080 17629
rect 17408 17663 17460 17672
rect 17408 17629 17417 17663
rect 17417 17629 17451 17663
rect 17451 17629 17460 17663
rect 17408 17620 17460 17629
rect 13176 17552 13228 17604
rect 16948 17552 17000 17604
rect 17684 17663 17736 17672
rect 17684 17629 17693 17663
rect 17693 17629 17727 17663
rect 17727 17629 17736 17663
rect 17684 17620 17736 17629
rect 20536 17688 20588 17740
rect 22008 17688 22060 17740
rect 17960 17552 18012 17604
rect 18972 17620 19024 17672
rect 20260 17663 20312 17672
rect 20260 17629 20269 17663
rect 20269 17629 20303 17663
rect 20303 17629 20312 17663
rect 20260 17620 20312 17629
rect 21180 17620 21232 17672
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 11428 17484 11480 17536
rect 15108 17484 15160 17536
rect 15384 17484 15436 17536
rect 17040 17484 17092 17536
rect 19892 17552 19944 17604
rect 22560 17620 22612 17672
rect 22836 17663 22888 17672
rect 22836 17629 22845 17663
rect 22845 17629 22879 17663
rect 22879 17629 22888 17663
rect 22836 17620 22888 17629
rect 23020 17620 23072 17672
rect 23112 17620 23164 17672
rect 26976 17688 27028 17740
rect 29552 17688 29604 17740
rect 31668 17688 31720 17740
rect 23756 17620 23808 17672
rect 22100 17552 22152 17604
rect 27436 17620 27488 17672
rect 28816 17663 28868 17672
rect 28816 17629 28825 17663
rect 28825 17629 28859 17663
rect 28859 17629 28868 17663
rect 28816 17620 28868 17629
rect 21088 17484 21140 17536
rect 21824 17527 21876 17536
rect 21824 17493 21833 17527
rect 21833 17493 21867 17527
rect 21867 17493 21876 17527
rect 21824 17484 21876 17493
rect 22008 17484 22060 17536
rect 22836 17484 22888 17536
rect 29276 17552 29328 17604
rect 29644 17620 29696 17672
rect 30104 17663 30156 17672
rect 30104 17629 30113 17663
rect 30113 17629 30147 17663
rect 30147 17629 30156 17663
rect 30104 17620 30156 17629
rect 29828 17595 29880 17604
rect 29828 17561 29837 17595
rect 29837 17561 29871 17595
rect 29871 17561 29880 17595
rect 29828 17552 29880 17561
rect 30012 17552 30064 17604
rect 30564 17620 30616 17672
rect 32772 17620 32824 17672
rect 29644 17484 29696 17536
rect 30472 17552 30524 17604
rect 30288 17484 30340 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 3056 17280 3108 17332
rect 2780 17144 2832 17196
rect 4252 17280 4304 17332
rect 3608 17212 3660 17264
rect 5540 17280 5592 17332
rect 5632 17280 5684 17332
rect 7196 17280 7248 17332
rect 7932 17280 7984 17332
rect 4804 17212 4856 17264
rect 3976 17187 4028 17196
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 1676 17119 1728 17128
rect 1676 17085 1685 17119
rect 1685 17085 1719 17119
rect 1719 17085 1728 17119
rect 1676 17076 1728 17085
rect 4344 17187 4396 17196
rect 4344 17153 4353 17187
rect 4353 17153 4387 17187
rect 4387 17153 4396 17187
rect 4344 17144 4396 17153
rect 4528 17144 4580 17196
rect 5356 17212 5408 17264
rect 6920 17212 6972 17264
rect 5724 17144 5776 17196
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 5908 17187 5960 17196
rect 5908 17153 5917 17187
rect 5917 17153 5951 17187
rect 5951 17153 5960 17187
rect 5908 17144 5960 17153
rect 7564 17255 7616 17264
rect 7564 17221 7573 17255
rect 7573 17221 7607 17255
rect 7607 17221 7616 17255
rect 7564 17212 7616 17221
rect 9312 17280 9364 17332
rect 9772 17280 9824 17332
rect 9956 17323 10008 17332
rect 9956 17289 9965 17323
rect 9965 17289 9999 17323
rect 9999 17289 10008 17323
rect 9956 17280 10008 17289
rect 10048 17280 10100 17332
rect 10600 17280 10652 17332
rect 11336 17280 11388 17332
rect 11704 17280 11756 17332
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 12624 17323 12676 17332
rect 12624 17289 12633 17323
rect 12633 17289 12667 17323
rect 12667 17289 12676 17323
rect 12624 17280 12676 17289
rect 15292 17323 15344 17332
rect 15292 17289 15301 17323
rect 15301 17289 15335 17323
rect 15335 17289 15344 17323
rect 15292 17280 15344 17289
rect 21364 17280 21416 17332
rect 30656 17280 30708 17332
rect 8852 17144 8904 17196
rect 4804 17076 4856 17128
rect 5264 17076 5316 17128
rect 6460 17076 6512 17128
rect 7012 17119 7064 17128
rect 7012 17085 7021 17119
rect 7021 17085 7055 17119
rect 7055 17085 7064 17119
rect 7012 17076 7064 17085
rect 2320 16940 2372 16992
rect 4068 17008 4120 17060
rect 9956 17144 10008 17196
rect 10416 17212 10468 17264
rect 10692 17212 10744 17264
rect 10508 17144 10560 17196
rect 12532 17212 12584 17264
rect 13544 17212 13596 17264
rect 9496 17076 9548 17128
rect 10324 17008 10376 17060
rect 11060 17076 11112 17128
rect 11244 17076 11296 17128
rect 12808 17144 12860 17196
rect 12992 17076 13044 17128
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 15660 17144 15712 17196
rect 17592 17212 17644 17264
rect 17960 17212 18012 17264
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 21916 17212 21968 17264
rect 19892 17144 19944 17196
rect 15200 17008 15252 17060
rect 18052 17076 18104 17128
rect 19340 17076 19392 17128
rect 16396 17008 16448 17060
rect 19892 17008 19944 17060
rect 4160 16940 4212 16992
rect 4804 16940 4856 16992
rect 10140 16940 10192 16992
rect 13820 16940 13872 16992
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 19340 16940 19392 16949
rect 20996 17144 21048 17196
rect 20720 17076 20772 17128
rect 21088 17076 21140 17128
rect 20168 17008 20220 17060
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 26332 17212 26384 17264
rect 30012 17212 30064 17264
rect 30288 17255 30340 17264
rect 30288 17221 30297 17255
rect 30297 17221 30331 17255
rect 30331 17221 30340 17255
rect 30288 17212 30340 17221
rect 32036 17280 32088 17332
rect 32956 17280 33008 17332
rect 22652 17144 22704 17196
rect 23388 17187 23440 17196
rect 23388 17153 23397 17187
rect 23397 17153 23431 17187
rect 23431 17153 23440 17187
rect 23388 17144 23440 17153
rect 24400 17144 24452 17196
rect 25136 17187 25188 17196
rect 25136 17153 25145 17187
rect 25145 17153 25179 17187
rect 25179 17153 25188 17187
rect 25136 17144 25188 17153
rect 25320 17144 25372 17196
rect 25504 17144 25556 17196
rect 27344 17187 27396 17196
rect 27344 17153 27353 17187
rect 27353 17153 27387 17187
rect 27387 17153 27396 17187
rect 27344 17144 27396 17153
rect 27620 17187 27672 17196
rect 27620 17153 27629 17187
rect 27629 17153 27663 17187
rect 27663 17153 27672 17187
rect 27620 17144 27672 17153
rect 27804 17144 27856 17196
rect 27988 17187 28040 17196
rect 27988 17153 27997 17187
rect 27997 17153 28031 17187
rect 28031 17153 28040 17187
rect 27988 17144 28040 17153
rect 30196 17144 30248 17196
rect 30564 17187 30616 17196
rect 30564 17153 30573 17187
rect 30573 17153 30607 17187
rect 30607 17153 30616 17187
rect 30564 17144 30616 17153
rect 31484 17187 31536 17196
rect 31484 17153 31491 17187
rect 31491 17153 31536 17187
rect 31484 17144 31536 17153
rect 22560 17076 22612 17128
rect 28816 17119 28868 17128
rect 28816 17085 28825 17119
rect 28825 17085 28859 17119
rect 28859 17085 28868 17119
rect 28816 17076 28868 17085
rect 25964 17008 26016 17060
rect 30656 17076 30708 17128
rect 31208 17076 31260 17128
rect 31668 17187 31720 17196
rect 31668 17153 31677 17187
rect 31677 17153 31711 17187
rect 31711 17153 31720 17187
rect 31668 17144 31720 17153
rect 31852 17144 31904 17196
rect 32220 17187 32272 17196
rect 32220 17153 32229 17187
rect 32229 17153 32263 17187
rect 32263 17153 32272 17187
rect 32220 17144 32272 17153
rect 32312 17144 32364 17196
rect 32496 17144 32548 17196
rect 32036 17076 32088 17128
rect 31944 17008 31996 17060
rect 21272 16940 21324 16992
rect 22560 16940 22612 16992
rect 27252 16940 27304 16992
rect 28448 16940 28500 16992
rect 29644 16940 29696 16992
rect 29736 16940 29788 16992
rect 34704 17008 34756 17060
rect 32312 16940 32364 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1676 16736 1728 16788
rect 3700 16736 3752 16788
rect 4436 16736 4488 16788
rect 5724 16736 5776 16788
rect 6092 16779 6144 16788
rect 6092 16745 6101 16779
rect 6101 16745 6135 16779
rect 6135 16745 6144 16779
rect 6092 16736 6144 16745
rect 9772 16779 9824 16788
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 10324 16779 10376 16788
rect 10324 16745 10333 16779
rect 10333 16745 10367 16779
rect 10367 16745 10376 16779
rect 10324 16736 10376 16745
rect 11612 16736 11664 16788
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 20628 16736 20680 16788
rect 20996 16736 21048 16788
rect 24032 16736 24084 16788
rect 25228 16736 25280 16788
rect 25596 16736 25648 16788
rect 26240 16736 26292 16788
rect 26332 16736 26384 16788
rect 2228 16668 2280 16720
rect 2412 16643 2464 16652
rect 2412 16609 2421 16643
rect 2421 16609 2455 16643
rect 2455 16609 2464 16643
rect 2412 16600 2464 16609
rect 2596 16600 2648 16652
rect 2320 16575 2372 16584
rect 2320 16541 2329 16575
rect 2329 16541 2363 16575
rect 2363 16541 2372 16575
rect 2320 16532 2372 16541
rect 3332 16575 3384 16584
rect 3332 16541 3341 16575
rect 3341 16541 3375 16575
rect 3375 16541 3384 16575
rect 3332 16532 3384 16541
rect 4344 16643 4396 16652
rect 4344 16609 4353 16643
rect 4353 16609 4387 16643
rect 4387 16609 4396 16643
rect 4344 16600 4396 16609
rect 4896 16600 4948 16652
rect 4436 16532 4488 16584
rect 5908 16668 5960 16720
rect 8392 16668 8444 16720
rect 6460 16600 6512 16652
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 9312 16600 9364 16652
rect 3700 16464 3752 16516
rect 4528 16507 4580 16516
rect 4528 16473 4537 16507
rect 4537 16473 4571 16507
rect 4571 16473 4580 16507
rect 4528 16464 4580 16473
rect 4620 16464 4672 16516
rect 5632 16507 5684 16516
rect 5632 16473 5641 16507
rect 5641 16473 5675 16507
rect 5675 16473 5684 16507
rect 5632 16464 5684 16473
rect 7104 16532 7156 16584
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 8944 16575 8996 16584
rect 8944 16541 8953 16575
rect 8953 16541 8987 16575
rect 8987 16541 8996 16575
rect 8944 16532 8996 16541
rect 12532 16668 12584 16720
rect 12716 16668 12768 16720
rect 18880 16668 18932 16720
rect 22008 16668 22060 16720
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 3608 16396 3660 16448
rect 4804 16396 4856 16448
rect 8576 16464 8628 16516
rect 7564 16396 7616 16448
rect 8300 16396 8352 16448
rect 9496 16464 9548 16516
rect 9680 16507 9732 16516
rect 9680 16473 9689 16507
rect 9689 16473 9723 16507
rect 9723 16473 9732 16507
rect 9680 16464 9732 16473
rect 8944 16396 8996 16448
rect 11060 16575 11112 16584
rect 11060 16541 11069 16575
rect 11069 16541 11103 16575
rect 11103 16541 11112 16575
rect 11060 16532 11112 16541
rect 11612 16575 11664 16584
rect 11612 16541 11621 16575
rect 11621 16541 11655 16575
rect 11655 16541 11664 16575
rect 11612 16532 11664 16541
rect 11704 16532 11756 16584
rect 12716 16532 12768 16584
rect 19340 16600 19392 16652
rect 23204 16668 23256 16720
rect 24216 16668 24268 16720
rect 25320 16668 25372 16720
rect 18328 16532 18380 16584
rect 22652 16643 22704 16652
rect 22652 16609 22661 16643
rect 22661 16609 22695 16643
rect 22695 16609 22704 16643
rect 22652 16600 22704 16609
rect 23388 16600 23440 16652
rect 22192 16532 22244 16584
rect 10600 16464 10652 16516
rect 13544 16464 13596 16516
rect 14188 16464 14240 16516
rect 15660 16464 15712 16516
rect 18052 16464 18104 16516
rect 21640 16464 21692 16516
rect 12072 16396 12124 16448
rect 23112 16396 23164 16448
rect 23940 16532 23992 16584
rect 24492 16532 24544 16584
rect 24860 16575 24912 16584
rect 25136 16600 25188 16652
rect 27620 16736 27672 16788
rect 28816 16736 28868 16788
rect 27160 16668 27212 16720
rect 27436 16668 27488 16720
rect 24860 16541 24905 16575
rect 24905 16541 24912 16575
rect 24860 16532 24912 16541
rect 25228 16532 25280 16584
rect 25688 16575 25740 16584
rect 25688 16541 25697 16575
rect 25697 16541 25731 16575
rect 25731 16541 25740 16575
rect 25688 16532 25740 16541
rect 26516 16575 26568 16584
rect 26516 16541 26525 16575
rect 26525 16541 26559 16575
rect 26559 16541 26568 16575
rect 26516 16532 26568 16541
rect 26608 16575 26660 16584
rect 26608 16541 26617 16575
rect 26617 16541 26651 16575
rect 26651 16541 26660 16575
rect 26608 16532 26660 16541
rect 26792 16575 26844 16584
rect 26792 16541 26801 16575
rect 26801 16541 26835 16575
rect 26835 16541 26844 16575
rect 26792 16532 26844 16541
rect 26976 16532 27028 16584
rect 27620 16600 27672 16652
rect 34060 16736 34112 16788
rect 32312 16643 32364 16652
rect 32312 16609 32321 16643
rect 32321 16609 32355 16643
rect 32355 16609 32364 16643
rect 32312 16600 32364 16609
rect 35256 16643 35308 16652
rect 35256 16609 35265 16643
rect 35265 16609 35299 16643
rect 35299 16609 35308 16643
rect 35256 16600 35308 16609
rect 27436 16532 27488 16584
rect 24676 16507 24728 16516
rect 24676 16473 24685 16507
rect 24685 16473 24719 16507
rect 24719 16473 24728 16507
rect 24676 16464 24728 16473
rect 26332 16464 26384 16516
rect 29184 16532 29236 16584
rect 33876 16532 33928 16584
rect 36084 16532 36136 16584
rect 27988 16396 28040 16448
rect 28264 16464 28316 16516
rect 30380 16464 30432 16516
rect 31300 16464 31352 16516
rect 33600 16464 33652 16516
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 3608 16235 3660 16244
rect 3608 16201 3617 16235
rect 3617 16201 3651 16235
rect 3651 16201 3660 16235
rect 3608 16192 3660 16201
rect 3884 16192 3936 16244
rect 8484 16192 8536 16244
rect 8668 16192 8720 16244
rect 9036 16235 9088 16244
rect 9036 16201 9045 16235
rect 9045 16201 9079 16235
rect 9079 16201 9088 16235
rect 9036 16192 9088 16201
rect 9680 16192 9732 16244
rect 11336 16235 11388 16244
rect 11336 16201 11345 16235
rect 11345 16201 11379 16235
rect 11379 16201 11388 16235
rect 11336 16192 11388 16201
rect 12992 16192 13044 16244
rect 4344 16124 4396 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 2780 16056 2832 16108
rect 4896 16056 4948 16108
rect 3884 16031 3936 16040
rect 3884 15997 3893 16031
rect 3893 15997 3927 16031
rect 3927 15997 3936 16031
rect 3884 15988 3936 15997
rect 2412 15852 2464 15904
rect 5080 15988 5132 16040
rect 6736 16124 6788 16176
rect 5356 16056 5408 16108
rect 5540 15988 5592 16040
rect 5816 15988 5868 16040
rect 7196 15988 7248 16040
rect 5724 15920 5776 15972
rect 4068 15852 4120 15904
rect 5448 15852 5500 15904
rect 12256 16167 12308 16176
rect 12256 16133 12265 16167
rect 12265 16133 12299 16167
rect 12299 16133 12308 16167
rect 12256 16124 12308 16133
rect 9312 16056 9364 16108
rect 10968 16056 11020 16108
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 12072 16099 12124 16108
rect 12072 16065 12081 16099
rect 12081 16065 12115 16099
rect 12115 16065 12124 16099
rect 12072 16056 12124 16065
rect 12440 16056 12492 16108
rect 12808 16056 12860 16108
rect 13820 16124 13872 16176
rect 8116 15852 8168 15904
rect 8760 15852 8812 15904
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 10600 15988 10652 16040
rect 12808 15963 12860 15972
rect 12808 15929 12817 15963
rect 12817 15929 12851 15963
rect 12851 15929 12860 15963
rect 12808 15920 12860 15929
rect 13544 16056 13596 16108
rect 17132 16235 17184 16244
rect 17132 16201 17141 16235
rect 17141 16201 17175 16235
rect 17175 16201 17184 16235
rect 17132 16192 17184 16201
rect 19340 16192 19392 16244
rect 19616 16192 19668 16244
rect 17224 16124 17276 16176
rect 21640 16124 21692 16176
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 14372 15920 14424 15972
rect 11244 15852 11296 15904
rect 13636 15852 13688 15904
rect 14188 15852 14240 15904
rect 14464 15852 14516 15904
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 15476 16056 15528 16108
rect 17592 16099 17644 16108
rect 17592 16065 17601 16099
rect 17601 16065 17635 16099
rect 17635 16065 17644 16099
rect 17592 16056 17644 16065
rect 17224 15988 17276 16040
rect 18696 15988 18748 16040
rect 19892 15988 19944 16040
rect 21548 15988 21600 16040
rect 16948 15920 17000 15972
rect 15200 15852 15252 15904
rect 15936 15852 15988 15904
rect 19156 15920 19208 15972
rect 19064 15852 19116 15904
rect 20536 15852 20588 15904
rect 21916 16056 21968 16108
rect 22284 16099 22336 16108
rect 22284 16065 22293 16099
rect 22293 16065 22327 16099
rect 22327 16065 22336 16099
rect 22284 16056 22336 16065
rect 23664 16124 23716 16176
rect 24216 16167 24268 16176
rect 24216 16133 24225 16167
rect 24225 16133 24259 16167
rect 24259 16133 24268 16167
rect 24216 16124 24268 16133
rect 24308 16167 24360 16176
rect 24308 16133 24317 16167
rect 24317 16133 24351 16167
rect 24351 16133 24360 16167
rect 24308 16124 24360 16133
rect 24952 16192 25004 16244
rect 25688 16192 25740 16244
rect 29736 16192 29788 16244
rect 32036 16192 32088 16244
rect 32588 16192 32640 16244
rect 33416 16192 33468 16244
rect 22100 15988 22152 16040
rect 22192 16031 22244 16040
rect 22192 15997 22201 16031
rect 22201 15997 22235 16031
rect 22235 15997 22244 16031
rect 22192 15988 22244 15997
rect 23480 15988 23532 16040
rect 23940 16099 23992 16108
rect 23940 16065 23949 16099
rect 23949 16065 23983 16099
rect 23983 16065 23992 16099
rect 23940 16056 23992 16065
rect 24032 16099 24084 16108
rect 24032 16065 24042 16099
rect 24042 16065 24076 16099
rect 24076 16065 24084 16099
rect 24032 16056 24084 16065
rect 24584 16056 24636 16108
rect 24768 16056 24820 16108
rect 24952 16099 25004 16108
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 26332 16124 26384 16176
rect 30472 16124 30524 16176
rect 31484 16124 31536 16176
rect 25228 16099 25280 16108
rect 25228 16065 25237 16099
rect 25237 16065 25271 16099
rect 25271 16065 25280 16099
rect 25228 16056 25280 16065
rect 26056 16099 26108 16108
rect 26056 16065 26065 16099
rect 26065 16065 26099 16099
rect 26099 16065 26108 16099
rect 26056 16056 26108 16065
rect 27896 16099 27948 16108
rect 27896 16065 27905 16099
rect 27905 16065 27939 16099
rect 27939 16065 27948 16099
rect 27896 16056 27948 16065
rect 28080 16099 28132 16108
rect 28080 16065 28089 16099
rect 28089 16065 28123 16099
rect 28123 16065 28132 16099
rect 28080 16056 28132 16065
rect 28264 16099 28316 16108
rect 28264 16065 28273 16099
rect 28273 16065 28307 16099
rect 28307 16065 28316 16099
rect 28264 16056 28316 16065
rect 26148 15988 26200 16040
rect 29276 16099 29328 16108
rect 29276 16065 29285 16099
rect 29285 16065 29319 16099
rect 29319 16065 29328 16099
rect 29276 16056 29328 16065
rect 29460 16056 29512 16108
rect 31024 16056 31076 16108
rect 30104 15988 30156 16040
rect 31760 16056 31812 16108
rect 31484 15988 31536 16040
rect 31576 15988 31628 16040
rect 22652 15920 22704 15972
rect 29368 15920 29420 15972
rect 23020 15852 23072 15904
rect 25320 15852 25372 15904
rect 27620 15852 27672 15904
rect 30748 15852 30800 15904
rect 31024 15852 31076 15904
rect 31668 15920 31720 15972
rect 34796 15852 34848 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4804 15648 4856 15700
rect 1400 15512 1452 15564
rect 1860 15555 1912 15564
rect 1860 15521 1869 15555
rect 1869 15521 1903 15555
rect 1903 15521 1912 15555
rect 1860 15512 1912 15521
rect 5080 15512 5132 15564
rect 5448 15648 5500 15700
rect 5632 15648 5684 15700
rect 3240 15444 3292 15496
rect 5356 15555 5408 15564
rect 5356 15521 5365 15555
rect 5365 15521 5399 15555
rect 5399 15521 5408 15555
rect 5356 15512 5408 15521
rect 6092 15512 6144 15564
rect 7104 15691 7156 15700
rect 7104 15657 7113 15691
rect 7113 15657 7147 15691
rect 7147 15657 7156 15691
rect 7104 15648 7156 15657
rect 7196 15691 7248 15700
rect 7196 15657 7205 15691
rect 7205 15657 7239 15691
rect 7239 15657 7248 15691
rect 7196 15648 7248 15657
rect 8208 15648 8260 15700
rect 9312 15691 9364 15700
rect 9312 15657 9321 15691
rect 9321 15657 9355 15691
rect 9355 15657 9364 15691
rect 9312 15648 9364 15657
rect 10600 15691 10652 15700
rect 10600 15657 10609 15691
rect 10609 15657 10643 15691
rect 10643 15657 10652 15691
rect 10600 15648 10652 15657
rect 16028 15648 16080 15700
rect 6736 15580 6788 15632
rect 8760 15580 8812 15632
rect 9128 15580 9180 15632
rect 12808 15580 12860 15632
rect 4804 15376 4856 15428
rect 2136 15308 2188 15360
rect 5264 15308 5316 15360
rect 6644 15308 6696 15360
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 7472 15376 7524 15428
rect 8024 15444 8076 15496
rect 8392 15512 8444 15564
rect 9496 15512 9548 15564
rect 8484 15444 8536 15496
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 9404 15444 9456 15496
rect 10232 15512 10284 15564
rect 11244 15555 11296 15564
rect 11244 15521 11253 15555
rect 11253 15521 11287 15555
rect 11287 15521 11296 15555
rect 11244 15512 11296 15521
rect 11336 15512 11388 15564
rect 14832 15580 14884 15632
rect 15108 15580 15160 15632
rect 14280 15512 14332 15564
rect 14648 15512 14700 15564
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 12532 15444 12584 15496
rect 12624 15487 12676 15496
rect 12624 15453 12633 15487
rect 12633 15453 12667 15487
rect 12667 15453 12676 15487
rect 12624 15444 12676 15453
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 14832 15487 14884 15496
rect 14832 15453 14842 15487
rect 14842 15453 14876 15487
rect 14876 15453 14884 15487
rect 14832 15444 14884 15453
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 15476 15444 15528 15496
rect 10876 15376 10928 15428
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 10232 15351 10284 15360
rect 10232 15317 10241 15351
rect 10241 15317 10275 15351
rect 10275 15317 10284 15351
rect 10232 15308 10284 15317
rect 10784 15308 10836 15360
rect 12164 15308 12216 15360
rect 13360 15308 13412 15360
rect 14924 15308 14976 15360
rect 15384 15351 15436 15360
rect 15384 15317 15393 15351
rect 15393 15317 15427 15351
rect 15427 15317 15436 15351
rect 15384 15308 15436 15317
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 19524 15648 19576 15700
rect 19800 15648 19852 15700
rect 18696 15580 18748 15632
rect 18420 15512 18472 15564
rect 19064 15487 19116 15496
rect 19064 15453 19073 15487
rect 19073 15453 19107 15487
rect 19107 15453 19116 15487
rect 19064 15444 19116 15453
rect 19616 15512 19668 15564
rect 19432 15444 19484 15496
rect 21364 15691 21416 15700
rect 21364 15657 21373 15691
rect 21373 15657 21407 15691
rect 21407 15657 21416 15691
rect 21364 15648 21416 15657
rect 30564 15648 30616 15700
rect 31208 15648 31260 15700
rect 32772 15648 32824 15700
rect 33968 15691 34020 15700
rect 33968 15657 33977 15691
rect 33977 15657 34011 15691
rect 34011 15657 34020 15691
rect 33968 15648 34020 15657
rect 34704 15691 34756 15700
rect 34704 15657 34713 15691
rect 34713 15657 34747 15691
rect 34747 15657 34756 15691
rect 34704 15648 34756 15657
rect 34796 15648 34848 15700
rect 21916 15580 21968 15632
rect 23112 15623 23164 15632
rect 23112 15589 23121 15623
rect 23121 15589 23155 15623
rect 23155 15589 23164 15623
rect 23112 15580 23164 15589
rect 26240 15580 26292 15632
rect 21548 15512 21600 15564
rect 25136 15512 25188 15564
rect 30472 15555 30524 15564
rect 30472 15521 30481 15555
rect 30481 15521 30515 15555
rect 30515 15521 30524 15555
rect 30472 15512 30524 15521
rect 15660 15376 15712 15428
rect 16948 15376 17000 15428
rect 17500 15376 17552 15428
rect 20628 15444 20680 15496
rect 20352 15376 20404 15428
rect 17316 15308 17368 15360
rect 17868 15308 17920 15360
rect 23020 15487 23072 15496
rect 23020 15453 23029 15487
rect 23029 15453 23063 15487
rect 23063 15453 23072 15487
rect 23020 15444 23072 15453
rect 23204 15444 23256 15496
rect 30656 15487 30708 15496
rect 30656 15453 30673 15487
rect 30673 15453 30708 15487
rect 30656 15444 30708 15453
rect 30748 15487 30800 15496
rect 30748 15453 30757 15487
rect 30757 15453 30791 15487
rect 30791 15453 30800 15487
rect 30748 15444 30800 15453
rect 31024 15444 31076 15496
rect 31208 15487 31260 15496
rect 31208 15453 31217 15487
rect 31217 15453 31251 15487
rect 31251 15453 31260 15487
rect 31208 15444 31260 15453
rect 21272 15376 21324 15428
rect 21180 15308 21232 15360
rect 24952 15376 25004 15428
rect 27344 15376 27396 15428
rect 28080 15308 28132 15360
rect 29828 15308 29880 15360
rect 30380 15376 30432 15428
rect 30564 15308 30616 15360
rect 30748 15308 30800 15360
rect 32864 15580 32916 15632
rect 32956 15580 33008 15632
rect 31576 15512 31628 15564
rect 31760 15512 31812 15564
rect 33140 15512 33192 15564
rect 34244 15580 34296 15632
rect 34612 15512 34664 15564
rect 31668 15487 31720 15496
rect 31668 15453 31682 15487
rect 31682 15453 31716 15487
rect 31716 15453 31720 15487
rect 31668 15444 31720 15453
rect 32956 15444 33008 15496
rect 34520 15444 34572 15496
rect 33140 15419 33192 15428
rect 33140 15385 33149 15419
rect 33149 15385 33183 15419
rect 33183 15385 33192 15419
rect 33140 15376 33192 15385
rect 31760 15308 31812 15360
rect 35532 15444 35584 15496
rect 34428 15351 34480 15360
rect 34428 15317 34437 15351
rect 34437 15317 34471 15351
rect 34471 15317 34480 15351
rect 34428 15308 34480 15317
rect 34612 15308 34664 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 1860 14968 1912 15020
rect 3240 15036 3292 15088
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 4068 15079 4120 15088
rect 4068 15045 4077 15079
rect 4077 15045 4111 15079
rect 4111 15045 4120 15079
rect 4068 15036 4120 15045
rect 4804 15036 4856 15088
rect 5724 14968 5776 15020
rect 6276 15036 6328 15088
rect 2228 14943 2280 14952
rect 2228 14909 2237 14943
rect 2237 14909 2271 14943
rect 2271 14909 2280 14943
rect 2228 14900 2280 14909
rect 2044 14764 2096 14816
rect 3700 14875 3752 14884
rect 3700 14841 3709 14875
rect 3709 14841 3743 14875
rect 3743 14841 3752 14875
rect 3700 14832 3752 14841
rect 5540 14900 5592 14952
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 9588 15104 9640 15156
rect 10140 15104 10192 15156
rect 8116 15079 8168 15088
rect 8116 15045 8125 15079
rect 8125 15045 8159 15079
rect 8159 15045 8168 15079
rect 8116 15036 8168 15045
rect 9772 15036 9824 15088
rect 9128 14900 9180 14952
rect 9312 14900 9364 14952
rect 9496 14900 9548 14952
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 10232 14900 10284 14952
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 14924 15036 14976 15088
rect 17684 15104 17736 15156
rect 18052 15104 18104 15156
rect 19064 15104 19116 15156
rect 19524 15104 19576 15156
rect 21456 15104 21508 15156
rect 23020 15104 23072 15156
rect 24676 15104 24728 15156
rect 26976 15104 27028 15156
rect 32128 15104 32180 15156
rect 32772 15147 32824 15156
rect 32772 15113 32781 15147
rect 32781 15113 32815 15147
rect 32815 15113 32824 15147
rect 32772 15104 32824 15113
rect 10876 14968 10928 15020
rect 20352 15036 20404 15088
rect 20812 15036 20864 15088
rect 23572 15036 23624 15088
rect 15200 14900 15252 14952
rect 15476 14968 15528 15020
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 17408 14968 17460 15020
rect 18604 14968 18656 15020
rect 19340 15011 19392 15020
rect 19340 14977 19349 15011
rect 19349 14977 19383 15011
rect 19383 14977 19392 15011
rect 19340 14968 19392 14977
rect 20536 15011 20588 15020
rect 20536 14977 20545 15011
rect 20545 14977 20579 15011
rect 20579 14977 20588 15011
rect 20536 14968 20588 14977
rect 16212 14900 16264 14952
rect 9404 14832 9456 14884
rect 10876 14832 10928 14884
rect 12532 14832 12584 14884
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 18052 14900 18104 14909
rect 18144 14943 18196 14952
rect 18144 14909 18153 14943
rect 18153 14909 18187 14943
rect 18187 14909 18196 14943
rect 18144 14900 18196 14909
rect 18328 14900 18380 14952
rect 19248 14900 19300 14952
rect 19432 14900 19484 14952
rect 20996 14900 21048 14952
rect 6092 14764 6144 14816
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 6644 14764 6696 14773
rect 7656 14764 7708 14816
rect 11060 14764 11112 14816
rect 15476 14764 15528 14816
rect 18972 14832 19024 14884
rect 20076 14832 20128 14884
rect 21364 14832 21416 14884
rect 23480 14968 23532 15020
rect 24032 14968 24084 15020
rect 25504 15036 25556 15088
rect 31852 15036 31904 15088
rect 32680 15036 32732 15088
rect 26240 14968 26292 15020
rect 27252 14968 27304 15020
rect 27712 15011 27764 15020
rect 27712 14977 27721 15011
rect 27721 14977 27755 15011
rect 27755 14977 27764 15011
rect 27712 14968 27764 14977
rect 31760 14968 31812 15020
rect 32312 15011 32364 15020
rect 32312 14977 32329 15011
rect 32329 14977 32364 15011
rect 32312 14968 32364 14977
rect 32956 14968 33008 15020
rect 24216 14943 24268 14952
rect 24216 14909 24225 14943
rect 24225 14909 24259 14943
rect 24259 14909 24268 14943
rect 24216 14900 24268 14909
rect 25228 14900 25280 14952
rect 25596 14900 25648 14952
rect 25780 14900 25832 14952
rect 22744 14832 22796 14884
rect 21548 14764 21600 14816
rect 30380 14832 30432 14884
rect 31392 14832 31444 14884
rect 33784 14832 33836 14884
rect 24584 14807 24636 14816
rect 24584 14773 24593 14807
rect 24593 14773 24627 14807
rect 24627 14773 24636 14807
rect 24584 14764 24636 14773
rect 24676 14807 24728 14816
rect 24676 14773 24685 14807
rect 24685 14773 24719 14807
rect 24719 14773 24728 14807
rect 24676 14764 24728 14773
rect 24768 14764 24820 14816
rect 25228 14764 25280 14816
rect 27436 14764 27488 14816
rect 34060 14764 34112 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2228 14560 2280 14612
rect 4712 14492 4764 14544
rect 1860 14467 1912 14476
rect 1860 14433 1869 14467
rect 1869 14433 1903 14467
rect 1903 14433 1912 14467
rect 1860 14424 1912 14433
rect 3792 14424 3844 14476
rect 4252 14467 4304 14476
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 5356 14424 5408 14476
rect 8484 14492 8536 14544
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 9772 14560 9824 14612
rect 10508 14560 10560 14612
rect 10692 14560 10744 14612
rect 13268 14560 13320 14612
rect 14924 14560 14976 14612
rect 18420 14560 18472 14612
rect 23020 14560 23072 14612
rect 24676 14560 24728 14612
rect 26148 14560 26200 14612
rect 27436 14603 27488 14612
rect 27436 14569 27445 14603
rect 27445 14569 27479 14603
rect 27479 14569 27488 14603
rect 27436 14560 27488 14569
rect 35256 14560 35308 14612
rect 35440 14560 35492 14612
rect 7288 14424 7340 14476
rect 8208 14424 8260 14476
rect 3240 14356 3292 14408
rect 3700 14356 3752 14408
rect 6000 14356 6052 14408
rect 2412 14288 2464 14340
rect 6828 14356 6880 14408
rect 8300 14356 8352 14408
rect 8668 14467 8720 14476
rect 8668 14433 8677 14467
rect 8677 14433 8711 14467
rect 8711 14433 8720 14467
rect 8668 14424 8720 14433
rect 10140 14492 10192 14544
rect 16212 14492 16264 14544
rect 19432 14492 19484 14544
rect 9772 14424 9824 14476
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 2504 14220 2556 14272
rect 3700 14220 3752 14272
rect 5356 14263 5408 14272
rect 5356 14229 5365 14263
rect 5365 14229 5399 14263
rect 5399 14229 5408 14263
rect 5356 14220 5408 14229
rect 5908 14263 5960 14272
rect 5908 14229 5917 14263
rect 5917 14229 5951 14263
rect 5951 14229 5960 14263
rect 5908 14220 5960 14229
rect 6368 14263 6420 14272
rect 6368 14229 6377 14263
rect 6377 14229 6411 14263
rect 6411 14229 6420 14263
rect 6368 14220 6420 14229
rect 7472 14288 7524 14340
rect 8484 14356 8536 14408
rect 9312 14356 9364 14408
rect 10508 14424 10560 14476
rect 12348 14424 12400 14476
rect 12900 14424 12952 14476
rect 13176 14424 13228 14476
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 13268 14399 13320 14408
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 18696 14424 18748 14476
rect 20720 14492 20772 14544
rect 21640 14492 21692 14544
rect 24492 14492 24544 14544
rect 25412 14535 25464 14544
rect 25412 14501 25421 14535
rect 25421 14501 25455 14535
rect 25455 14501 25464 14535
rect 25412 14492 25464 14501
rect 25964 14535 26016 14544
rect 25964 14501 25973 14535
rect 25973 14501 26007 14535
rect 26007 14501 26016 14535
rect 25964 14492 26016 14501
rect 27160 14492 27212 14544
rect 34244 14492 34296 14544
rect 13544 14399 13596 14408
rect 13544 14365 13553 14399
rect 13553 14365 13587 14399
rect 13587 14365 13596 14399
rect 13544 14356 13596 14365
rect 13912 14356 13964 14408
rect 17684 14356 17736 14408
rect 17960 14399 18012 14408
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 22560 14424 22612 14476
rect 23204 14424 23256 14476
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 8300 14220 8352 14272
rect 8852 14288 8904 14340
rect 9404 14220 9456 14272
rect 10048 14220 10100 14272
rect 13728 14288 13780 14340
rect 10416 14220 10468 14272
rect 14740 14220 14792 14272
rect 18052 14220 18104 14272
rect 18696 14220 18748 14272
rect 20076 14356 20128 14408
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 20720 14399 20772 14408
rect 20720 14365 20729 14399
rect 20729 14365 20763 14399
rect 20763 14365 20772 14399
rect 20720 14356 20772 14365
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 23388 14399 23440 14408
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 23572 14399 23624 14408
rect 23572 14365 23581 14399
rect 23581 14365 23615 14399
rect 23615 14365 23624 14399
rect 23572 14356 23624 14365
rect 23756 14399 23808 14408
rect 23756 14365 23765 14399
rect 23765 14365 23799 14399
rect 23799 14365 23808 14399
rect 23756 14356 23808 14365
rect 20904 14288 20956 14340
rect 22652 14288 22704 14340
rect 22928 14288 22980 14340
rect 25504 14399 25556 14408
rect 25504 14365 25513 14399
rect 25513 14365 25547 14399
rect 25547 14365 25556 14399
rect 25504 14356 25556 14365
rect 25872 14399 25924 14408
rect 25872 14365 25881 14399
rect 25881 14365 25915 14399
rect 25915 14365 25924 14399
rect 25872 14356 25924 14365
rect 26884 14424 26936 14476
rect 25596 14288 25648 14340
rect 26976 14399 27028 14408
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 27252 14356 27304 14408
rect 27068 14288 27120 14340
rect 27528 14288 27580 14340
rect 26148 14220 26200 14272
rect 26608 14220 26660 14272
rect 27712 14399 27764 14408
rect 27712 14365 27721 14399
rect 27721 14365 27755 14399
rect 27755 14365 27764 14399
rect 27712 14356 27764 14365
rect 27896 14399 27948 14408
rect 27896 14365 27905 14399
rect 27905 14365 27939 14399
rect 27939 14365 27948 14399
rect 27896 14356 27948 14365
rect 29644 14399 29696 14408
rect 29644 14365 29653 14399
rect 29653 14365 29687 14399
rect 29687 14365 29696 14399
rect 29644 14356 29696 14365
rect 30840 14424 30892 14476
rect 33508 14424 33560 14476
rect 31668 14356 31720 14408
rect 34060 14399 34112 14408
rect 34060 14365 34069 14399
rect 34069 14365 34103 14399
rect 34103 14365 34112 14399
rect 34060 14356 34112 14365
rect 28356 14288 28408 14340
rect 29092 14288 29144 14340
rect 28816 14220 28868 14272
rect 30012 14331 30064 14340
rect 30012 14297 30021 14331
rect 30021 14297 30055 14331
rect 30055 14297 30064 14331
rect 30012 14288 30064 14297
rect 30380 14288 30432 14340
rect 30472 14288 30524 14340
rect 30656 14288 30708 14340
rect 31208 14288 31260 14340
rect 31392 14288 31444 14340
rect 32312 14288 32364 14340
rect 33508 14288 33560 14340
rect 33692 14288 33744 14340
rect 34612 14288 34664 14340
rect 30196 14220 30248 14272
rect 33324 14220 33376 14272
rect 34520 14220 34572 14272
rect 34980 14220 35032 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 1860 14016 1912 14068
rect 2412 14016 2464 14068
rect 3700 14059 3752 14068
rect 3700 14025 3709 14059
rect 3709 14025 3743 14059
rect 3743 14025 3752 14059
rect 3700 14016 3752 14025
rect 6368 14016 6420 14068
rect 6828 14016 6880 14068
rect 2780 13880 2832 13932
rect 3240 13880 3292 13932
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 2044 13812 2096 13864
rect 6644 13948 6696 14000
rect 4252 13880 4304 13932
rect 4436 13812 4488 13864
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 4896 13880 4948 13932
rect 5540 13880 5592 13932
rect 5632 13923 5684 13932
rect 5632 13889 5641 13923
rect 5641 13889 5675 13923
rect 5675 13889 5684 13923
rect 5632 13880 5684 13889
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 7472 14016 7524 14068
rect 7840 14016 7892 14068
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 9036 14016 9088 14068
rect 8208 13948 8260 14000
rect 9404 13948 9456 14000
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 8024 13880 8076 13932
rect 2872 13744 2924 13796
rect 3976 13744 4028 13796
rect 4804 13744 4856 13796
rect 3056 13676 3108 13728
rect 5448 13787 5500 13796
rect 5448 13753 5457 13787
rect 5457 13753 5491 13787
rect 5491 13753 5500 13787
rect 5448 13744 5500 13753
rect 5724 13744 5776 13796
rect 6276 13812 6328 13864
rect 6736 13744 6788 13796
rect 8484 13855 8536 13864
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 8944 13923 8996 13932
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 9128 13880 9180 13932
rect 10784 14016 10836 14068
rect 11520 14016 11572 14068
rect 13912 14059 13964 14068
rect 13912 14025 13921 14059
rect 13921 14025 13955 14059
rect 13955 14025 13964 14059
rect 13912 14016 13964 14025
rect 15752 14016 15804 14068
rect 16948 14016 17000 14068
rect 17684 14016 17736 14068
rect 21364 14059 21416 14068
rect 21364 14025 21373 14059
rect 21373 14025 21407 14059
rect 21407 14025 21416 14059
rect 21364 14016 21416 14025
rect 21548 14016 21600 14068
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 10968 13880 11020 13932
rect 12900 13948 12952 14000
rect 12716 13880 12768 13932
rect 14004 13880 14056 13932
rect 14740 13880 14792 13932
rect 8852 13812 8904 13864
rect 9036 13812 9088 13864
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 13084 13812 13136 13864
rect 15016 13812 15068 13864
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 17868 13948 17920 14000
rect 16948 13923 17000 13932
rect 16948 13889 16957 13923
rect 16957 13889 16991 13923
rect 16991 13889 17000 13923
rect 16948 13880 17000 13889
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 17316 13880 17368 13932
rect 19156 13880 19208 13932
rect 21824 13948 21876 14000
rect 25872 14016 25924 14068
rect 26148 14059 26200 14068
rect 26148 14025 26157 14059
rect 26157 14025 26191 14059
rect 26191 14025 26200 14059
rect 26148 14016 26200 14025
rect 27896 14016 27948 14068
rect 30656 14016 30708 14068
rect 30840 14016 30892 14068
rect 17592 13812 17644 13864
rect 8668 13676 8720 13728
rect 8852 13719 8904 13728
rect 8852 13685 8861 13719
rect 8861 13685 8895 13719
rect 8895 13685 8904 13719
rect 8852 13676 8904 13685
rect 9496 13676 9548 13728
rect 12440 13744 12492 13796
rect 12716 13744 12768 13796
rect 19800 13812 19852 13864
rect 20536 13812 20588 13864
rect 21640 13880 21692 13932
rect 22560 13923 22612 13932
rect 22560 13889 22569 13923
rect 22569 13889 22603 13923
rect 22603 13889 22612 13923
rect 22560 13880 22612 13889
rect 22652 13880 22704 13932
rect 23204 13880 23256 13932
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24492 13923 24544 13932
rect 24492 13889 24501 13923
rect 24501 13889 24535 13923
rect 24535 13889 24544 13923
rect 24492 13880 24544 13889
rect 24952 13880 25004 13932
rect 25320 13812 25372 13864
rect 27160 13948 27212 14000
rect 26700 13880 26752 13932
rect 27804 13948 27856 14000
rect 29092 13948 29144 14000
rect 29828 13948 29880 14000
rect 26332 13812 26384 13864
rect 27528 13812 27580 13864
rect 28816 13880 28868 13932
rect 28908 13923 28960 13932
rect 28908 13889 28917 13923
rect 28917 13889 28951 13923
rect 28951 13889 28960 13923
rect 28908 13880 28960 13889
rect 29000 13923 29052 13932
rect 29000 13889 29009 13923
rect 29009 13889 29043 13923
rect 29043 13889 29052 13923
rect 29000 13880 29052 13889
rect 30932 13880 30984 13932
rect 32496 14016 32548 14068
rect 33232 14016 33284 14068
rect 33784 14016 33836 14068
rect 34336 14016 34388 14068
rect 34520 14016 34572 14068
rect 31208 13948 31260 14000
rect 33324 13948 33376 14000
rect 29920 13812 29972 13864
rect 31668 13880 31720 13932
rect 32772 13880 32824 13932
rect 33968 13880 34020 13932
rect 34152 13880 34204 13932
rect 35072 13923 35124 13932
rect 35072 13889 35081 13923
rect 35081 13889 35115 13923
rect 35115 13889 35124 13923
rect 35072 13880 35124 13889
rect 35440 14016 35492 14068
rect 31760 13812 31812 13864
rect 32496 13855 32548 13864
rect 32496 13821 32505 13855
rect 32505 13821 32539 13855
rect 32539 13821 32548 13855
rect 32496 13812 32548 13821
rect 33232 13812 33284 13864
rect 19892 13744 19944 13796
rect 21364 13744 21416 13796
rect 22376 13744 22428 13796
rect 22928 13744 22980 13796
rect 23388 13744 23440 13796
rect 25688 13744 25740 13796
rect 29460 13744 29512 13796
rect 30932 13744 30984 13796
rect 35256 13812 35308 13864
rect 10416 13676 10468 13728
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 15016 13676 15068 13728
rect 15292 13676 15344 13728
rect 18236 13676 18288 13728
rect 18328 13676 18380 13728
rect 22468 13676 22520 13728
rect 25412 13719 25464 13728
rect 25412 13685 25421 13719
rect 25421 13685 25455 13719
rect 25455 13685 25464 13719
rect 25412 13676 25464 13685
rect 26424 13676 26476 13728
rect 31116 13676 31168 13728
rect 31484 13676 31536 13728
rect 33692 13676 33744 13728
rect 34796 13676 34848 13728
rect 34980 13676 35032 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1676 13472 1728 13524
rect 4436 13515 4488 13524
rect 4436 13481 4445 13515
rect 4445 13481 4479 13515
rect 4479 13481 4488 13515
rect 4436 13472 4488 13481
rect 4712 13472 4764 13524
rect 5356 13472 5408 13524
rect 5816 13472 5868 13524
rect 6736 13472 6788 13524
rect 9772 13472 9824 13524
rect 9864 13472 9916 13524
rect 12532 13472 12584 13524
rect 14740 13515 14792 13524
rect 14740 13481 14749 13515
rect 14749 13481 14783 13515
rect 14783 13481 14792 13515
rect 14740 13472 14792 13481
rect 5264 13404 5316 13456
rect 6552 13404 6604 13456
rect 2872 13379 2924 13388
rect 2872 13345 2881 13379
rect 2881 13345 2915 13379
rect 2915 13345 2924 13379
rect 2872 13336 2924 13345
rect 3056 13379 3108 13388
rect 3056 13345 3065 13379
rect 3065 13345 3099 13379
rect 3099 13345 3108 13379
rect 3056 13336 3108 13345
rect 4988 13336 5040 13388
rect 5816 13336 5868 13388
rect 7748 13404 7800 13456
rect 3240 13200 3292 13252
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 4160 13243 4212 13252
rect 4160 13209 4169 13243
rect 4169 13209 4203 13243
rect 4203 13209 4212 13243
rect 4160 13200 4212 13209
rect 5724 13268 5776 13320
rect 7104 13336 7156 13388
rect 7380 13379 7432 13388
rect 7380 13345 7389 13379
rect 7389 13345 7423 13379
rect 7423 13345 7432 13379
rect 7380 13336 7432 13345
rect 4528 13132 4580 13184
rect 4712 13132 4764 13184
rect 6000 13200 6052 13252
rect 6184 13200 6236 13252
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 7012 13268 7064 13320
rect 7472 13268 7524 13320
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 6828 13200 6880 13252
rect 7748 13200 7800 13252
rect 7932 13200 7984 13252
rect 5356 13175 5408 13184
rect 5356 13141 5365 13175
rect 5365 13141 5399 13175
rect 5399 13141 5408 13175
rect 5356 13132 5408 13141
rect 5448 13132 5500 13184
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 8024 13132 8076 13184
rect 8208 13175 8260 13184
rect 8208 13141 8217 13175
rect 8217 13141 8251 13175
rect 8251 13141 8260 13175
rect 8208 13132 8260 13141
rect 9220 13404 9272 13456
rect 10692 13404 10744 13456
rect 8668 13268 8720 13320
rect 9404 13268 9456 13320
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10324 13243 10376 13252
rect 10324 13209 10333 13243
rect 10333 13209 10367 13243
rect 10367 13209 10376 13243
rect 10324 13200 10376 13209
rect 9956 13132 10008 13184
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 14648 13379 14700 13388
rect 14648 13345 14657 13379
rect 14657 13345 14691 13379
rect 14691 13345 14700 13379
rect 14648 13336 14700 13345
rect 17132 13472 17184 13524
rect 19340 13472 19392 13524
rect 20168 13472 20220 13524
rect 22744 13472 22796 13524
rect 24492 13472 24544 13524
rect 26424 13515 26476 13524
rect 26424 13481 26433 13515
rect 26433 13481 26467 13515
rect 26467 13481 26476 13515
rect 26424 13472 26476 13481
rect 29000 13472 29052 13524
rect 30288 13515 30340 13524
rect 30288 13481 30297 13515
rect 30297 13481 30331 13515
rect 30331 13481 30340 13515
rect 30288 13472 30340 13481
rect 30564 13472 30616 13524
rect 31392 13472 31444 13524
rect 33232 13472 33284 13524
rect 34612 13472 34664 13524
rect 34796 13472 34848 13524
rect 35256 13472 35308 13524
rect 35808 13472 35860 13524
rect 17592 13404 17644 13456
rect 19524 13447 19576 13456
rect 19524 13413 19533 13447
rect 19533 13413 19567 13447
rect 19567 13413 19576 13447
rect 19524 13404 19576 13413
rect 19892 13404 19944 13456
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 12900 13268 12952 13320
rect 13636 13268 13688 13320
rect 14004 13268 14056 13320
rect 11520 13200 11572 13252
rect 14280 13200 14332 13252
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 15752 13268 15804 13320
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 16580 13268 16632 13320
rect 17960 13336 18012 13388
rect 17408 13268 17460 13320
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 17500 13200 17552 13252
rect 18328 13268 18380 13320
rect 19156 13200 19208 13252
rect 19340 13200 19392 13252
rect 21548 13404 21600 13456
rect 20536 13336 20588 13388
rect 29644 13336 29696 13388
rect 31852 13404 31904 13456
rect 30288 13336 30340 13388
rect 30656 13336 30708 13388
rect 31576 13336 31628 13388
rect 34060 13404 34112 13456
rect 32496 13379 32548 13388
rect 32496 13345 32505 13379
rect 32505 13345 32539 13379
rect 32539 13345 32548 13379
rect 32496 13336 32548 13345
rect 19892 13268 19944 13320
rect 20168 13268 20220 13320
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 20444 13200 20496 13252
rect 12808 13132 12860 13184
rect 13176 13132 13228 13184
rect 15016 13132 15068 13184
rect 18880 13132 18932 13184
rect 19708 13132 19760 13184
rect 20812 13132 20864 13184
rect 28816 13200 28868 13252
rect 29644 13200 29696 13252
rect 30104 13200 30156 13252
rect 30288 13200 30340 13252
rect 26976 13132 27028 13184
rect 27344 13132 27396 13184
rect 30656 13243 30708 13252
rect 30656 13209 30665 13243
rect 30665 13209 30699 13243
rect 30699 13209 30708 13243
rect 30656 13200 30708 13209
rect 30840 13311 30892 13320
rect 30840 13277 30849 13311
rect 30849 13277 30883 13311
rect 30883 13277 30892 13311
rect 30840 13268 30892 13277
rect 32312 13268 32364 13320
rect 32956 13311 33008 13320
rect 32956 13277 32965 13311
rect 32965 13277 32999 13311
rect 32999 13277 33008 13311
rect 32956 13268 33008 13277
rect 33600 13268 33652 13320
rect 34520 13268 34572 13320
rect 31024 13200 31076 13252
rect 31760 13200 31812 13252
rect 32772 13243 32824 13252
rect 32772 13209 32781 13243
rect 32781 13209 32815 13243
rect 32815 13209 32824 13243
rect 32772 13200 32824 13209
rect 32864 13243 32916 13252
rect 32864 13209 32873 13243
rect 32873 13209 32907 13243
rect 32907 13209 32916 13243
rect 32864 13200 32916 13209
rect 31484 13132 31536 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 3148 12971 3200 12980
rect 3148 12937 3157 12971
rect 3157 12937 3191 12971
rect 3191 12937 3200 12971
rect 3148 12928 3200 12937
rect 3240 12971 3292 12980
rect 3240 12937 3249 12971
rect 3249 12937 3283 12971
rect 3283 12937 3292 12971
rect 3240 12928 3292 12937
rect 5264 12928 5316 12980
rect 5816 12971 5868 12980
rect 4436 12860 4488 12912
rect 2780 12792 2832 12844
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 4068 12792 4120 12844
rect 4804 12835 4856 12844
rect 4804 12801 4808 12835
rect 4808 12801 4842 12835
rect 4842 12801 4856 12835
rect 4804 12792 4856 12801
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 3700 12767 3752 12776
rect 3700 12733 3709 12767
rect 3709 12733 3743 12767
rect 3743 12733 3752 12767
rect 3700 12724 3752 12733
rect 3056 12656 3108 12708
rect 4712 12724 4764 12776
rect 4528 12656 4580 12708
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5172 12835 5224 12844
rect 5172 12801 5180 12835
rect 5180 12801 5214 12835
rect 5214 12801 5224 12835
rect 5172 12792 5224 12801
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 6920 12928 6972 12980
rect 7196 12928 7248 12980
rect 8208 12928 8260 12980
rect 8576 12928 8628 12980
rect 8944 12928 8996 12980
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 10324 12928 10376 12980
rect 11428 12928 11480 12980
rect 14280 12971 14332 12980
rect 14280 12937 14289 12971
rect 14289 12937 14323 12971
rect 14323 12937 14332 12971
rect 14280 12928 14332 12937
rect 19340 12928 19392 12980
rect 6644 12860 6696 12912
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 6460 12792 6512 12844
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 6368 12724 6420 12776
rect 8024 12860 8076 12912
rect 7288 12792 7340 12844
rect 7196 12724 7248 12776
rect 3884 12588 3936 12640
rect 6920 12656 6972 12708
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 8300 12792 8352 12801
rect 8484 12860 8536 12912
rect 9588 12860 9640 12912
rect 10508 12860 10560 12912
rect 14188 12860 14240 12912
rect 16488 12860 16540 12912
rect 9128 12792 9180 12844
rect 10048 12792 10100 12844
rect 10692 12792 10744 12844
rect 7748 12724 7800 12776
rect 8760 12724 8812 12776
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 14372 12724 14424 12776
rect 14832 12792 14884 12844
rect 15844 12792 15896 12844
rect 19708 12835 19760 12844
rect 19708 12801 19717 12835
rect 19717 12801 19751 12835
rect 19751 12801 19760 12835
rect 19708 12792 19760 12801
rect 20168 12792 20220 12844
rect 21732 12792 21784 12844
rect 21916 12792 21968 12844
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 14924 12724 14976 12776
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 17500 12724 17552 12776
rect 22284 12971 22336 12980
rect 22284 12937 22293 12971
rect 22293 12937 22327 12971
rect 22327 12937 22336 12971
rect 22284 12928 22336 12937
rect 23020 12903 23072 12912
rect 23020 12869 23045 12903
rect 23045 12869 23072 12903
rect 24400 12928 24452 12980
rect 29460 12928 29512 12980
rect 32864 12928 32916 12980
rect 23020 12860 23072 12869
rect 23480 12860 23532 12912
rect 22928 12792 22980 12844
rect 32680 12792 32732 12844
rect 32864 12792 32916 12844
rect 8300 12656 8352 12708
rect 8852 12656 8904 12708
rect 5448 12588 5500 12640
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 6184 12588 6236 12640
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 7932 12588 7984 12640
rect 8208 12588 8260 12640
rect 9680 12656 9732 12708
rect 10416 12656 10468 12708
rect 17408 12656 17460 12708
rect 19340 12656 19392 12708
rect 25044 12724 25096 12776
rect 22468 12656 22520 12708
rect 9128 12588 9180 12640
rect 9956 12588 10008 12640
rect 10784 12588 10836 12640
rect 14648 12631 14700 12640
rect 14648 12597 14657 12631
rect 14657 12597 14691 12631
rect 14691 12597 14700 12631
rect 14648 12588 14700 12597
rect 20076 12588 20128 12640
rect 20352 12588 20404 12640
rect 20536 12588 20588 12640
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 22100 12588 22152 12640
rect 22376 12588 22428 12640
rect 26608 12656 26660 12708
rect 23204 12631 23256 12640
rect 23204 12597 23213 12631
rect 23213 12597 23247 12631
rect 23247 12597 23256 12631
rect 23204 12588 23256 12597
rect 23572 12588 23624 12640
rect 24308 12588 24360 12640
rect 26424 12588 26476 12640
rect 28816 12588 28868 12640
rect 29828 12588 29880 12640
rect 32680 12588 32732 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1676 12384 1728 12436
rect 3608 12384 3660 12436
rect 3884 12384 3936 12436
rect 4252 12384 4304 12436
rect 2412 12248 2464 12300
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 2228 12180 2280 12232
rect 2964 12316 3016 12368
rect 3148 12316 3200 12368
rect 4712 12359 4764 12368
rect 4712 12325 4721 12359
rect 4721 12325 4755 12359
rect 4755 12325 4764 12359
rect 4712 12316 4764 12325
rect 3056 12223 3108 12232
rect 3056 12189 3064 12223
rect 3064 12189 3098 12223
rect 3098 12189 3108 12223
rect 3056 12180 3108 12189
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 2872 12155 2924 12164
rect 2872 12121 2881 12155
rect 2881 12121 2915 12155
rect 2915 12121 2924 12155
rect 2872 12112 2924 12121
rect 3700 12248 3752 12300
rect 3792 12248 3844 12300
rect 3332 12180 3384 12232
rect 3608 12223 3660 12232
rect 3608 12189 3617 12223
rect 3617 12189 3651 12223
rect 3651 12189 3660 12223
rect 3608 12180 3660 12189
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 4344 12180 4396 12232
rect 4620 12248 4672 12300
rect 5908 12384 5960 12436
rect 6920 12384 6972 12436
rect 7196 12384 7248 12436
rect 8024 12384 8076 12436
rect 5448 12316 5500 12368
rect 5724 12291 5776 12300
rect 5724 12257 5733 12291
rect 5733 12257 5767 12291
rect 5767 12257 5776 12291
rect 5724 12248 5776 12257
rect 7564 12316 7616 12368
rect 6920 12248 6972 12300
rect 7288 12248 7340 12300
rect 7932 12316 7984 12368
rect 8668 12384 8720 12436
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 10048 12384 10100 12436
rect 13084 12427 13136 12436
rect 13084 12393 13093 12427
rect 13093 12393 13127 12427
rect 13127 12393 13136 12427
rect 13084 12384 13136 12393
rect 15384 12427 15436 12436
rect 15384 12393 15393 12427
rect 15393 12393 15427 12427
rect 15427 12393 15436 12427
rect 15384 12384 15436 12393
rect 15568 12384 15620 12436
rect 15936 12384 15988 12436
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 18236 12384 18288 12436
rect 18972 12384 19024 12436
rect 21732 12384 21784 12436
rect 22468 12384 22520 12436
rect 23940 12384 23992 12436
rect 24584 12384 24636 12436
rect 25964 12384 26016 12436
rect 27620 12427 27672 12436
rect 27620 12393 27629 12427
rect 27629 12393 27663 12427
rect 27663 12393 27672 12427
rect 27620 12384 27672 12393
rect 28080 12427 28132 12436
rect 28080 12393 28089 12427
rect 28089 12393 28123 12427
rect 28123 12393 28132 12427
rect 28080 12384 28132 12393
rect 28356 12384 28408 12436
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 8484 12316 8536 12368
rect 4160 12112 4212 12164
rect 3608 12044 3660 12096
rect 4896 12180 4948 12232
rect 4620 12112 4672 12164
rect 5448 12180 5500 12232
rect 5632 12112 5684 12164
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 6736 12180 6788 12232
rect 4804 12044 4856 12096
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 6460 12112 6512 12164
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 8668 12248 8720 12300
rect 9496 12316 9548 12368
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 8208 12180 8260 12232
rect 8576 12155 8628 12164
rect 6644 12044 6696 12096
rect 8576 12121 8585 12155
rect 8585 12121 8619 12155
rect 8619 12121 8628 12155
rect 8576 12112 8628 12121
rect 7472 12087 7524 12096
rect 7472 12053 7481 12087
rect 7481 12053 7515 12087
rect 7515 12053 7524 12087
rect 7472 12044 7524 12053
rect 7564 12087 7616 12096
rect 7564 12053 7573 12087
rect 7573 12053 7607 12087
rect 7607 12053 7616 12087
rect 7564 12044 7616 12053
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 10140 12316 10192 12368
rect 10876 12316 10928 12368
rect 14372 12316 14424 12368
rect 10048 12248 10100 12300
rect 11704 12248 11756 12300
rect 15752 12316 15804 12368
rect 17776 12316 17828 12368
rect 19156 12316 19208 12368
rect 20260 12316 20312 12368
rect 22100 12316 22152 12368
rect 22560 12316 22612 12368
rect 23388 12316 23440 12368
rect 10140 12180 10192 12232
rect 10600 12180 10652 12232
rect 10876 12180 10928 12232
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 12256 12180 12308 12232
rect 10048 12112 10100 12164
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 17224 12248 17276 12300
rect 18328 12291 18380 12300
rect 18328 12257 18337 12291
rect 18337 12257 18371 12291
rect 18371 12257 18380 12291
rect 18328 12248 18380 12257
rect 21088 12248 21140 12300
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 13636 12112 13688 12164
rect 14280 12155 14332 12164
rect 14280 12121 14289 12155
rect 14289 12121 14323 12155
rect 14323 12121 14332 12155
rect 14280 12112 14332 12121
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15200 12180 15252 12189
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 18144 12180 18196 12232
rect 19064 12180 19116 12232
rect 23020 12248 23072 12300
rect 11060 12044 11112 12096
rect 11336 12044 11388 12096
rect 12900 12044 12952 12096
rect 14188 12044 14240 12096
rect 14556 12044 14608 12096
rect 16488 12112 16540 12164
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 21732 12180 21784 12232
rect 22284 12180 22336 12232
rect 16672 12044 16724 12096
rect 17408 12044 17460 12096
rect 18328 12044 18380 12096
rect 18604 12044 18656 12096
rect 19708 12112 19760 12164
rect 22744 12180 22796 12232
rect 23572 12180 23624 12232
rect 24308 12180 24360 12232
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 25044 12223 25096 12232
rect 25044 12189 25053 12223
rect 25053 12189 25087 12223
rect 25087 12189 25096 12223
rect 25044 12180 25096 12189
rect 26608 12316 26660 12368
rect 27528 12316 27580 12368
rect 25688 12248 25740 12300
rect 27068 12248 27120 12300
rect 29184 12316 29236 12368
rect 29736 12316 29788 12368
rect 20812 12044 20864 12096
rect 21088 12044 21140 12096
rect 21180 12044 21232 12096
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 22468 12044 22520 12096
rect 23020 12087 23072 12096
rect 23020 12053 23029 12087
rect 23029 12053 23063 12087
rect 23063 12053 23072 12087
rect 23020 12044 23072 12053
rect 23204 12044 23256 12096
rect 23940 12112 23992 12164
rect 24860 12112 24912 12164
rect 25872 12180 25924 12232
rect 26884 12180 26936 12232
rect 29644 12248 29696 12300
rect 27620 12180 27672 12232
rect 25596 12155 25648 12164
rect 25596 12121 25605 12155
rect 25605 12121 25639 12155
rect 25639 12121 25648 12155
rect 25596 12112 25648 12121
rect 25964 12112 26016 12164
rect 27988 12180 28040 12232
rect 28172 12180 28224 12232
rect 24400 12044 24452 12096
rect 25320 12044 25372 12096
rect 29184 12180 29236 12232
rect 30196 12427 30248 12436
rect 30196 12393 30205 12427
rect 30205 12393 30239 12427
rect 30239 12393 30248 12427
rect 30196 12384 30248 12393
rect 29092 12112 29144 12164
rect 29460 12112 29512 12164
rect 29552 12112 29604 12164
rect 29828 12155 29880 12164
rect 29828 12121 29837 12155
rect 29837 12121 29871 12155
rect 29871 12121 29880 12155
rect 29828 12112 29880 12121
rect 30472 12180 30524 12232
rect 30564 12223 30616 12232
rect 30564 12189 30573 12223
rect 30573 12189 30607 12223
rect 30607 12189 30616 12223
rect 30564 12180 30616 12189
rect 31668 12384 31720 12436
rect 33508 12384 33560 12436
rect 34704 12384 34756 12436
rect 34796 12384 34848 12436
rect 30840 12190 30892 12242
rect 31024 12223 31076 12232
rect 31024 12189 31038 12223
rect 31038 12189 31072 12223
rect 31072 12189 31076 12223
rect 31024 12180 31076 12189
rect 34060 12316 34112 12368
rect 32312 12248 32364 12300
rect 32128 12180 32180 12232
rect 32864 12248 32916 12300
rect 33692 12248 33744 12300
rect 34152 12248 34204 12300
rect 33048 12180 33100 12232
rect 34336 12223 34388 12232
rect 34336 12189 34345 12223
rect 34345 12189 34379 12223
rect 34379 12189 34388 12223
rect 34336 12180 34388 12189
rect 34796 12180 34848 12232
rect 31208 12044 31260 12096
rect 31484 12044 31536 12096
rect 31944 12112 31996 12164
rect 34060 12112 34112 12164
rect 34980 12155 35032 12164
rect 34980 12121 34989 12155
rect 34989 12121 35023 12155
rect 35023 12121 35032 12155
rect 34980 12112 35032 12121
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 2412 11883 2464 11892
rect 2412 11849 2421 11883
rect 2421 11849 2455 11883
rect 2455 11849 2464 11883
rect 2412 11840 2464 11849
rect 3148 11840 3200 11892
rect 3332 11840 3384 11892
rect 4160 11840 4212 11892
rect 4620 11840 4672 11892
rect 5908 11883 5960 11892
rect 5908 11849 5917 11883
rect 5917 11849 5951 11883
rect 5951 11849 5960 11883
rect 5908 11840 5960 11849
rect 6000 11883 6052 11892
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 6552 11840 6604 11892
rect 6736 11840 6788 11892
rect 7472 11840 7524 11892
rect 2504 11704 2556 11756
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 6276 11772 6328 11824
rect 3608 11636 3660 11688
rect 4344 11636 4396 11688
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 5264 11747 5316 11756
rect 5264 11713 5273 11747
rect 5273 11713 5307 11747
rect 5307 11713 5316 11747
rect 5264 11704 5316 11713
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 5632 11704 5684 11756
rect 5816 11704 5868 11756
rect 6184 11747 6236 11756
rect 6184 11713 6193 11747
rect 6193 11713 6227 11747
rect 6227 11713 6236 11747
rect 6184 11704 6236 11713
rect 6644 11747 6696 11756
rect 6644 11713 6648 11747
rect 6648 11713 6682 11747
rect 6682 11713 6696 11747
rect 6644 11704 6696 11713
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 7288 11772 7340 11824
rect 3056 11568 3108 11620
rect 3516 11568 3568 11620
rect 5908 11636 5960 11688
rect 6092 11636 6144 11688
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 8668 11840 8720 11892
rect 9404 11840 9456 11892
rect 9496 11840 9548 11892
rect 9956 11840 10008 11892
rect 10048 11883 10100 11892
rect 10048 11849 10057 11883
rect 10057 11849 10091 11883
rect 10091 11849 10100 11883
rect 10048 11840 10100 11849
rect 10324 11840 10376 11892
rect 10692 11840 10744 11892
rect 8116 11772 8168 11824
rect 7380 11704 7432 11713
rect 8300 11747 8352 11756
rect 8300 11713 8309 11747
rect 8309 11713 8343 11747
rect 8343 11713 8352 11747
rect 8300 11704 8352 11713
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 8576 11636 8628 11688
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 9588 11704 9640 11756
rect 11980 11772 12032 11824
rect 9312 11636 9364 11688
rect 10600 11704 10652 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 14188 11772 14240 11824
rect 15476 11772 15528 11824
rect 16672 11883 16724 11892
rect 16672 11849 16681 11883
rect 16681 11849 16715 11883
rect 16715 11849 16724 11883
rect 16672 11840 16724 11849
rect 16764 11840 16816 11892
rect 10508 11636 10560 11688
rect 11520 11679 11572 11688
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 4896 11500 4948 11552
rect 5724 11568 5776 11620
rect 7380 11568 7432 11620
rect 8852 11568 8904 11620
rect 13176 11704 13228 11756
rect 13452 11704 13504 11756
rect 14556 11704 14608 11756
rect 15200 11704 15252 11756
rect 12440 11636 12492 11688
rect 12808 11636 12860 11688
rect 13360 11636 13412 11688
rect 15752 11704 15804 11756
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 16764 11636 16816 11688
rect 19708 11840 19760 11892
rect 19892 11840 19944 11892
rect 20536 11840 20588 11892
rect 23020 11840 23072 11892
rect 23480 11840 23532 11892
rect 26700 11883 26752 11892
rect 26700 11849 26709 11883
rect 26709 11849 26743 11883
rect 26743 11849 26752 11883
rect 26700 11840 26752 11849
rect 27528 11840 27580 11892
rect 20168 11772 20220 11824
rect 17224 11704 17276 11756
rect 17592 11747 17644 11756
rect 17592 11713 17601 11747
rect 17601 11713 17635 11747
rect 17635 11713 17644 11747
rect 17592 11704 17644 11713
rect 17684 11747 17736 11756
rect 17684 11713 17693 11747
rect 17693 11713 17727 11747
rect 17727 11713 17736 11747
rect 17684 11704 17736 11713
rect 17868 11747 17920 11756
rect 17868 11713 17877 11747
rect 17877 11713 17911 11747
rect 17911 11713 17920 11747
rect 17868 11704 17920 11713
rect 17960 11747 18012 11756
rect 17960 11713 17969 11747
rect 17969 11713 18003 11747
rect 18003 11713 18012 11747
rect 17960 11704 18012 11713
rect 19156 11704 19208 11756
rect 19892 11704 19944 11756
rect 20260 11704 20312 11756
rect 20536 11747 20588 11756
rect 20536 11713 20545 11747
rect 20545 11713 20579 11747
rect 20579 11713 20588 11747
rect 20536 11704 20588 11713
rect 22284 11772 22336 11824
rect 23204 11772 23256 11824
rect 25044 11772 25096 11824
rect 21548 11704 21600 11756
rect 17500 11636 17552 11688
rect 24032 11704 24084 11756
rect 26700 11704 26752 11756
rect 27160 11704 27212 11756
rect 27252 11747 27304 11756
rect 27252 11713 27261 11747
rect 27261 11713 27295 11747
rect 27295 11713 27304 11747
rect 27252 11704 27304 11713
rect 27620 11704 27672 11756
rect 27712 11747 27764 11756
rect 27712 11713 27721 11747
rect 27721 11713 27755 11747
rect 27755 11713 27764 11747
rect 27712 11704 27764 11713
rect 30564 11840 30616 11892
rect 31024 11840 31076 11892
rect 31760 11840 31812 11892
rect 29368 11772 29420 11824
rect 30656 11772 30708 11824
rect 32772 11840 32824 11892
rect 32864 11840 32916 11892
rect 34336 11840 34388 11892
rect 29000 11704 29052 11756
rect 25320 11636 25372 11688
rect 30104 11747 30156 11756
rect 30104 11713 30113 11747
rect 30113 11713 30147 11747
rect 30147 11713 30156 11747
rect 30104 11704 30156 11713
rect 30288 11747 30340 11756
rect 30288 11713 30305 11747
rect 30305 11713 30340 11747
rect 30288 11704 30340 11713
rect 30380 11747 30432 11756
rect 30380 11713 30389 11747
rect 30389 11713 30423 11747
rect 30423 11713 30432 11747
rect 30380 11704 30432 11713
rect 31024 11704 31076 11756
rect 32956 11815 33008 11824
rect 32956 11781 32965 11815
rect 32965 11781 32999 11815
rect 32999 11781 33008 11815
rect 32956 11772 33008 11781
rect 34520 11772 34572 11824
rect 31392 11704 31444 11756
rect 32680 11747 32732 11756
rect 32680 11713 32689 11747
rect 32689 11713 32723 11747
rect 32723 11713 32732 11747
rect 32680 11704 32732 11713
rect 13636 11568 13688 11620
rect 17868 11568 17920 11620
rect 17960 11568 18012 11620
rect 5632 11500 5684 11552
rect 8944 11500 8996 11552
rect 10508 11500 10560 11552
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 16764 11500 16816 11552
rect 18512 11500 18564 11552
rect 19708 11500 19760 11552
rect 20720 11500 20772 11552
rect 21456 11568 21508 11620
rect 22652 11500 22704 11552
rect 25504 11500 25556 11552
rect 27528 11543 27580 11552
rect 27528 11509 27537 11543
rect 27537 11509 27571 11543
rect 27571 11509 27580 11543
rect 27528 11500 27580 11509
rect 28080 11611 28132 11620
rect 28080 11577 28089 11611
rect 28089 11577 28123 11611
rect 28123 11577 28132 11611
rect 28080 11568 28132 11577
rect 32404 11636 32456 11688
rect 35440 11636 35492 11688
rect 36084 11679 36136 11688
rect 36084 11645 36093 11679
rect 36093 11645 36127 11679
rect 36127 11645 36136 11679
rect 36084 11636 36136 11645
rect 29460 11568 29512 11620
rect 29552 11568 29604 11620
rect 34704 11568 34756 11620
rect 29000 11500 29052 11552
rect 33048 11543 33100 11552
rect 33048 11509 33057 11543
rect 33057 11509 33091 11543
rect 33091 11509 33100 11543
rect 33048 11500 33100 11509
rect 34796 11500 34848 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2872 11296 2924 11348
rect 2412 11228 2464 11280
rect 3332 11228 3384 11280
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 2596 11092 2648 11101
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 2504 11024 2556 11076
rect 3148 11092 3200 11144
rect 6460 11296 6512 11348
rect 5264 11228 5316 11280
rect 5540 11228 5592 11280
rect 8484 11228 8536 11280
rect 8668 11228 8720 11280
rect 10876 11296 10928 11348
rect 11152 11296 11204 11348
rect 12440 11296 12492 11348
rect 12532 11339 12584 11348
rect 12532 11305 12541 11339
rect 12541 11305 12575 11339
rect 12575 11305 12584 11339
rect 12532 11296 12584 11305
rect 12900 11339 12952 11348
rect 12900 11305 12909 11339
rect 12909 11305 12943 11339
rect 12943 11305 12952 11339
rect 12900 11296 12952 11305
rect 16856 11296 16908 11348
rect 4804 11160 4856 11212
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 4988 11135 5040 11144
rect 4988 11101 4998 11135
rect 4998 11101 5032 11135
rect 5032 11101 5040 11135
rect 4988 11092 5040 11101
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 5724 11092 5776 11144
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 6736 11160 6788 11212
rect 7380 11203 7432 11212
rect 7380 11169 7389 11203
rect 7389 11169 7423 11203
rect 7423 11169 7432 11203
rect 7380 11160 7432 11169
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 7012 11092 7064 11144
rect 5632 11024 5684 11076
rect 3056 10956 3108 11008
rect 3700 10956 3752 11008
rect 4160 10956 4212 11008
rect 4252 10956 4304 11008
rect 4712 10956 4764 11008
rect 5448 10956 5500 11008
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 5908 11024 5960 11076
rect 6828 10956 6880 11008
rect 7748 11024 7800 11076
rect 8300 11092 8352 11144
rect 9128 11092 9180 11144
rect 9312 11092 9364 11144
rect 9956 11135 10008 11144
rect 9956 11101 9965 11135
rect 9965 11101 9999 11135
rect 9999 11101 10008 11135
rect 9956 11092 10008 11101
rect 11704 11228 11756 11280
rect 17224 11271 17276 11280
rect 17224 11237 17233 11271
rect 17233 11237 17267 11271
rect 17267 11237 17276 11271
rect 17224 11228 17276 11237
rect 8668 11024 8720 11076
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 12532 11160 12584 11212
rect 13728 11160 13780 11212
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 12716 11092 12768 11144
rect 10508 11024 10560 11076
rect 8484 10956 8536 11008
rect 9220 10956 9272 11008
rect 10232 10999 10284 11008
rect 10232 10965 10241 10999
rect 10241 10965 10275 10999
rect 10275 10965 10284 10999
rect 10232 10956 10284 10965
rect 13452 11092 13504 11144
rect 14004 11092 14056 11144
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 14556 11135 14608 11144
rect 14556 11101 14565 11135
rect 14565 11101 14599 11135
rect 14599 11101 14608 11135
rect 14556 11092 14608 11101
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 15292 11160 15344 11212
rect 16488 11160 16540 11212
rect 17684 11228 17736 11280
rect 18144 11228 18196 11280
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 19708 11296 19760 11348
rect 22100 11296 22152 11348
rect 23020 11296 23072 11348
rect 23296 11296 23348 11348
rect 23480 11339 23532 11348
rect 23480 11305 23489 11339
rect 23489 11305 23523 11339
rect 23523 11305 23532 11339
rect 23480 11296 23532 11305
rect 24308 11296 24360 11348
rect 26608 11296 26660 11348
rect 26792 11296 26844 11348
rect 27620 11339 27672 11348
rect 27620 11305 27629 11339
rect 27629 11305 27663 11339
rect 27663 11305 27672 11339
rect 27620 11296 27672 11305
rect 19984 11228 20036 11280
rect 27252 11228 27304 11280
rect 29736 11296 29788 11348
rect 31760 11296 31812 11348
rect 32588 11339 32640 11348
rect 32588 11305 32597 11339
rect 32597 11305 32631 11339
rect 32631 11305 32640 11339
rect 32588 11296 32640 11305
rect 16672 11092 16724 11144
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 12532 10956 12584 11008
rect 15200 11024 15252 11076
rect 17224 11067 17276 11076
rect 17224 11033 17233 11067
rect 17233 11033 17267 11067
rect 17267 11033 17276 11067
rect 19616 11160 19668 11212
rect 19708 11160 19760 11212
rect 20168 11160 20220 11212
rect 20536 11092 20588 11144
rect 17224 11024 17276 11033
rect 20628 11024 20680 11076
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 22744 11135 22796 11144
rect 22744 11101 22753 11135
rect 22753 11101 22787 11135
rect 22787 11101 22796 11135
rect 22744 11092 22796 11101
rect 24768 11160 24820 11212
rect 26516 11160 26568 11212
rect 26792 11160 26844 11212
rect 23020 11135 23072 11144
rect 23020 11101 23029 11135
rect 23029 11101 23063 11135
rect 23063 11101 23072 11135
rect 23020 11092 23072 11101
rect 23388 11092 23440 11144
rect 27804 11160 27856 11212
rect 28540 11228 28592 11280
rect 31300 11228 31352 11280
rect 31668 11228 31720 11280
rect 23112 11024 23164 11076
rect 13452 10956 13504 11008
rect 14648 10956 14700 11008
rect 18052 10956 18104 11008
rect 18236 10999 18288 11008
rect 18236 10965 18245 10999
rect 18245 10965 18279 10999
rect 18279 10965 18288 10999
rect 18236 10956 18288 10965
rect 18512 10956 18564 11008
rect 20260 10956 20312 11008
rect 24400 11067 24452 11076
rect 24400 11033 24409 11067
rect 24409 11033 24443 11067
rect 24443 11033 24452 11067
rect 24400 11024 24452 11033
rect 24860 11024 24912 11076
rect 25320 11024 25372 11076
rect 27160 11024 27212 11076
rect 23572 10956 23624 11008
rect 24216 10956 24268 11008
rect 27988 11135 28040 11144
rect 27988 11101 27997 11135
rect 27997 11101 28031 11135
rect 28031 11101 28040 11135
rect 27988 11092 28040 11101
rect 28172 11135 28224 11144
rect 28172 11101 28181 11135
rect 28181 11101 28215 11135
rect 28215 11101 28224 11135
rect 28172 11092 28224 11101
rect 28356 11135 28408 11144
rect 28356 11101 28365 11135
rect 28365 11101 28399 11135
rect 28399 11101 28408 11135
rect 28356 11092 28408 11101
rect 28816 11092 28868 11144
rect 29000 11135 29052 11144
rect 29000 11101 29009 11135
rect 29009 11101 29043 11135
rect 29043 11101 29052 11135
rect 29000 11092 29052 11101
rect 29092 11135 29144 11144
rect 29092 11101 29101 11135
rect 29101 11101 29135 11135
rect 29135 11101 29144 11135
rect 29092 11092 29144 11101
rect 31944 11203 31996 11212
rect 31944 11169 31953 11203
rect 31953 11169 31987 11203
rect 31987 11169 31996 11203
rect 31944 11160 31996 11169
rect 32404 11228 32456 11280
rect 32772 11228 32824 11280
rect 33048 11296 33100 11348
rect 33140 11296 33192 11348
rect 34520 11296 34572 11348
rect 34704 11296 34756 11348
rect 34888 11339 34940 11348
rect 34888 11305 34897 11339
rect 34897 11305 34931 11339
rect 34931 11305 34940 11339
rect 34888 11296 34940 11305
rect 34980 11228 35032 11280
rect 28540 11024 28592 11076
rect 28448 10956 28500 11008
rect 28724 10999 28776 11008
rect 28724 10965 28733 10999
rect 28733 10965 28767 10999
rect 28767 10965 28776 10999
rect 28724 10956 28776 10965
rect 29000 10956 29052 11008
rect 29552 11135 29604 11144
rect 29552 11101 29561 11135
rect 29561 11101 29595 11135
rect 29595 11101 29604 11135
rect 29552 11092 29604 11101
rect 31392 11092 31444 11144
rect 31576 11067 31628 11076
rect 31576 11033 31603 11067
rect 31603 11033 31628 11067
rect 31576 11024 31628 11033
rect 31668 11024 31720 11076
rect 32036 11092 32088 11144
rect 34520 11160 34572 11212
rect 32312 11135 32364 11144
rect 32312 11101 32321 11135
rect 32321 11101 32355 11135
rect 32355 11101 32364 11135
rect 32312 11092 32364 11101
rect 32864 11092 32916 11144
rect 34796 11135 34848 11144
rect 34796 11101 34805 11135
rect 34805 11101 34839 11135
rect 34839 11101 34848 11135
rect 34796 11092 34848 11101
rect 35348 11135 35400 11144
rect 35348 11101 35357 11135
rect 35357 11101 35391 11135
rect 35391 11101 35400 11135
rect 35348 11092 35400 11101
rect 33048 11067 33100 11076
rect 33048 11033 33057 11067
rect 33057 11033 33091 11067
rect 33091 11033 33100 11067
rect 33048 11024 33100 11033
rect 29552 10956 29604 11008
rect 29736 10999 29788 11008
rect 29736 10965 29745 10999
rect 29745 10965 29779 10999
rect 29779 10965 29788 10999
rect 29736 10956 29788 10965
rect 31852 10956 31904 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 3148 10795 3200 10804
rect 3148 10761 3157 10795
rect 3157 10761 3191 10795
rect 3191 10761 3200 10795
rect 3148 10752 3200 10761
rect 3424 10752 3476 10804
rect 2964 10684 3016 10736
rect 3700 10727 3752 10736
rect 3700 10693 3709 10727
rect 3709 10693 3743 10727
rect 3743 10693 3752 10727
rect 3700 10684 3752 10693
rect 5448 10752 5500 10804
rect 5540 10752 5592 10804
rect 7012 10752 7064 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 3608 10616 3660 10668
rect 3884 10616 3936 10668
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 3792 10548 3844 10600
rect 4804 10659 4856 10668
rect 4804 10625 4813 10659
rect 4813 10625 4847 10659
rect 4847 10625 4856 10659
rect 4804 10616 4856 10625
rect 5816 10684 5868 10736
rect 1676 10412 1728 10464
rect 2320 10412 2372 10464
rect 3332 10412 3384 10464
rect 3608 10412 3660 10464
rect 4712 10591 4764 10600
rect 4712 10557 4721 10591
rect 4721 10557 4755 10591
rect 4755 10557 4764 10591
rect 4712 10548 4764 10557
rect 5264 10480 5316 10532
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 8576 10684 8628 10736
rect 8760 10684 8812 10736
rect 8668 10548 8720 10600
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9128 10616 9180 10668
rect 9404 10659 9456 10668
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 12716 10752 12768 10804
rect 21088 10752 21140 10804
rect 21272 10752 21324 10804
rect 21824 10752 21876 10804
rect 23848 10752 23900 10804
rect 24216 10795 24268 10804
rect 24216 10761 24225 10795
rect 24225 10761 24259 10795
rect 24259 10761 24268 10795
rect 24216 10752 24268 10761
rect 25136 10752 25188 10804
rect 25780 10752 25832 10804
rect 27712 10752 27764 10804
rect 27804 10752 27856 10804
rect 28356 10752 28408 10804
rect 28816 10752 28868 10804
rect 10416 10684 10468 10736
rect 11980 10684 12032 10736
rect 18512 10684 18564 10736
rect 18788 10684 18840 10736
rect 20628 10684 20680 10736
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 10232 10548 10284 10600
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 15568 10548 15620 10600
rect 6644 10480 6696 10532
rect 8116 10480 8168 10532
rect 12072 10480 12124 10532
rect 3976 10412 4028 10464
rect 4068 10412 4120 10464
rect 4896 10412 4948 10464
rect 9496 10412 9548 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 15016 10412 15068 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 17776 10616 17828 10668
rect 17960 10616 18012 10668
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 18972 10616 19024 10668
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 19340 10616 19392 10668
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 20996 10684 21048 10736
rect 17684 10591 17736 10600
rect 17684 10557 17693 10591
rect 17693 10557 17727 10591
rect 17727 10557 17736 10591
rect 17684 10548 17736 10557
rect 18696 10548 18748 10600
rect 19524 10548 19576 10600
rect 19892 10591 19944 10600
rect 19892 10557 19901 10591
rect 19901 10557 19935 10591
rect 19935 10557 19944 10591
rect 19892 10548 19944 10557
rect 17868 10412 17920 10464
rect 18328 10412 18380 10464
rect 18512 10455 18564 10464
rect 18512 10421 18521 10455
rect 18521 10421 18555 10455
rect 18555 10421 18564 10455
rect 18512 10412 18564 10421
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 22928 10727 22980 10736
rect 22928 10693 22937 10727
rect 22937 10693 22971 10727
rect 22971 10693 22980 10727
rect 22928 10684 22980 10693
rect 21272 10616 21324 10668
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 23112 10659 23164 10668
rect 23112 10625 23121 10659
rect 23121 10625 23155 10659
rect 23155 10625 23164 10659
rect 23112 10616 23164 10625
rect 24768 10684 24820 10736
rect 28908 10684 28960 10736
rect 29644 10795 29696 10804
rect 29644 10761 29653 10795
rect 29653 10761 29687 10795
rect 29687 10761 29696 10795
rect 29644 10752 29696 10761
rect 31668 10752 31720 10804
rect 29828 10684 29880 10736
rect 30748 10684 30800 10736
rect 31116 10684 31168 10736
rect 32404 10795 32456 10804
rect 32404 10761 32413 10795
rect 32413 10761 32447 10795
rect 32447 10761 32456 10795
rect 32404 10752 32456 10761
rect 24584 10616 24636 10668
rect 28080 10616 28132 10668
rect 28724 10659 28776 10668
rect 28724 10625 28733 10659
rect 28733 10625 28767 10659
rect 28767 10625 28776 10659
rect 28724 10616 28776 10625
rect 29000 10659 29052 10668
rect 29000 10625 29009 10659
rect 29009 10625 29043 10659
rect 29043 10625 29052 10659
rect 29000 10616 29052 10625
rect 29736 10616 29788 10668
rect 30380 10659 30432 10668
rect 30380 10625 30389 10659
rect 30389 10625 30423 10659
rect 30423 10625 30432 10659
rect 30380 10616 30432 10625
rect 31668 10659 31720 10668
rect 31668 10625 31677 10659
rect 31677 10625 31711 10659
rect 31711 10625 31720 10659
rect 31668 10616 31720 10625
rect 20996 10548 21048 10600
rect 22744 10548 22796 10600
rect 23848 10548 23900 10600
rect 27620 10548 27672 10600
rect 28540 10548 28592 10600
rect 28816 10548 28868 10600
rect 29552 10548 29604 10600
rect 30564 10548 30616 10600
rect 31576 10548 31628 10600
rect 32404 10616 32456 10668
rect 32772 10684 32824 10736
rect 19892 10412 19944 10464
rect 20260 10412 20312 10464
rect 20812 10455 20864 10464
rect 20812 10421 20821 10455
rect 20821 10421 20855 10455
rect 20855 10421 20864 10455
rect 20812 10412 20864 10421
rect 20996 10412 21048 10464
rect 22560 10480 22612 10532
rect 24768 10480 24820 10532
rect 27528 10480 27580 10532
rect 29092 10480 29144 10532
rect 31760 10480 31812 10532
rect 23848 10412 23900 10464
rect 24400 10412 24452 10464
rect 26240 10412 26292 10464
rect 26608 10412 26660 10464
rect 28080 10412 28132 10464
rect 28448 10412 28500 10464
rect 29184 10412 29236 10464
rect 29552 10412 29604 10464
rect 30288 10412 30340 10464
rect 32864 10659 32916 10668
rect 32864 10625 32873 10659
rect 32873 10625 32907 10659
rect 32907 10625 32916 10659
rect 32864 10616 32916 10625
rect 34428 10684 34480 10736
rect 34980 10684 35032 10736
rect 33508 10548 33560 10600
rect 34152 10480 34204 10532
rect 33416 10412 33468 10464
rect 34336 10412 34388 10464
rect 34980 10412 35032 10464
rect 35532 10412 35584 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2596 10208 2648 10260
rect 3792 10251 3844 10260
rect 3792 10217 3801 10251
rect 3801 10217 3835 10251
rect 3835 10217 3844 10251
rect 3792 10208 3844 10217
rect 3884 10208 3936 10260
rect 5908 10208 5960 10260
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2872 10140 2924 10192
rect 3240 10140 3292 10192
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 4896 10140 4948 10192
rect 3608 10072 3660 10124
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 3884 10004 3936 10056
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 5356 10072 5408 10124
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4252 10047 4304 10056
rect 4252 10013 4287 10047
rect 4287 10013 4304 10047
rect 4252 10004 4304 10013
rect 2504 9936 2556 9988
rect 3148 9936 3200 9988
rect 2412 9868 2464 9920
rect 3976 9868 4028 9920
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 4896 10004 4948 10056
rect 6000 10140 6052 10192
rect 5908 10047 5960 10056
rect 5908 10013 5922 10047
rect 5922 10013 5956 10047
rect 5956 10013 5960 10047
rect 6920 10140 6972 10192
rect 8300 10140 8352 10192
rect 12072 10208 12124 10260
rect 6368 10072 6420 10124
rect 5908 10004 5960 10013
rect 5632 9936 5684 9988
rect 5724 9979 5776 9988
rect 5724 9945 5733 9979
rect 5733 9945 5767 9979
rect 5767 9945 5776 9979
rect 5724 9936 5776 9945
rect 6276 9936 6328 9988
rect 7656 10004 7708 10056
rect 7840 10004 7892 10056
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 8760 10072 8812 10124
rect 9036 10115 9088 10124
rect 9036 10081 9045 10115
rect 9045 10081 9079 10115
rect 9079 10081 9088 10115
rect 9036 10072 9088 10081
rect 11888 10140 11940 10192
rect 15476 10208 15528 10260
rect 15568 10208 15620 10260
rect 19616 10208 19668 10260
rect 20076 10208 20128 10260
rect 20812 10251 20864 10260
rect 20812 10217 20821 10251
rect 20821 10217 20855 10251
rect 20855 10217 20864 10251
rect 20812 10208 20864 10217
rect 20996 10251 21048 10260
rect 20996 10217 21005 10251
rect 21005 10217 21039 10251
rect 21039 10217 21048 10251
rect 20996 10208 21048 10217
rect 22652 10208 22704 10260
rect 23204 10251 23256 10260
rect 23204 10217 23213 10251
rect 23213 10217 23247 10251
rect 23247 10217 23256 10251
rect 23204 10208 23256 10217
rect 24400 10208 24452 10260
rect 24492 10251 24544 10260
rect 24492 10217 24501 10251
rect 24501 10217 24535 10251
rect 24535 10217 24544 10251
rect 24492 10208 24544 10217
rect 25044 10251 25096 10260
rect 25044 10217 25053 10251
rect 25053 10217 25087 10251
rect 25087 10217 25096 10251
rect 25044 10208 25096 10217
rect 25504 10251 25556 10260
rect 25504 10217 25513 10251
rect 25513 10217 25547 10251
rect 25547 10217 25556 10251
rect 25504 10208 25556 10217
rect 25780 10208 25832 10260
rect 11612 10072 11664 10124
rect 12532 10072 12584 10124
rect 13912 10072 13964 10124
rect 17040 10140 17092 10192
rect 18604 10140 18656 10192
rect 19984 10140 20036 10192
rect 7196 9936 7248 9988
rect 8944 10004 8996 10056
rect 10692 10004 10744 10056
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 11520 10004 11572 10056
rect 12256 10004 12308 10056
rect 13452 10004 13504 10056
rect 4712 9868 4764 9920
rect 5908 9868 5960 9920
rect 6552 9868 6604 9920
rect 7104 9911 7156 9920
rect 7104 9877 7113 9911
rect 7113 9877 7147 9911
rect 7147 9877 7156 9911
rect 7104 9868 7156 9877
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 8300 9936 8352 9988
rect 8484 9979 8536 9988
rect 8484 9945 8493 9979
rect 8493 9945 8527 9979
rect 8527 9945 8536 9979
rect 8484 9936 8536 9945
rect 9312 9979 9364 9988
rect 9312 9945 9321 9979
rect 9321 9945 9355 9979
rect 9355 9945 9364 9979
rect 9312 9936 9364 9945
rect 12716 9979 12768 9988
rect 12716 9945 12725 9979
rect 12725 9945 12759 9979
rect 12759 9945 12768 9979
rect 12716 9936 12768 9945
rect 12808 9936 12860 9988
rect 15016 10047 15068 10056
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 15384 10004 15436 10056
rect 22468 10072 22520 10124
rect 26056 10072 26108 10124
rect 17776 10004 17828 10056
rect 18236 10004 18288 10056
rect 21180 10047 21232 10056
rect 21180 10013 21189 10047
rect 21189 10013 21223 10047
rect 21223 10013 21232 10047
rect 21180 10004 21232 10013
rect 21548 10004 21600 10056
rect 8116 9868 8168 9920
rect 8944 9868 8996 9920
rect 14556 9868 14608 9920
rect 21456 9936 21508 9988
rect 23848 9936 23900 9988
rect 17408 9868 17460 9920
rect 17868 9868 17920 9920
rect 18052 9868 18104 9920
rect 22928 9868 22980 9920
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 25320 10047 25372 10056
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 25412 10047 25464 10056
rect 25412 10013 25421 10047
rect 25421 10013 25455 10047
rect 25455 10013 25464 10047
rect 25412 10004 25464 10013
rect 24400 9936 24452 9988
rect 25964 10004 26016 10056
rect 26240 10047 26292 10056
rect 26240 10013 26249 10047
rect 26249 10013 26283 10047
rect 26283 10013 26292 10047
rect 26240 10004 26292 10013
rect 26976 10208 27028 10260
rect 27528 10140 27580 10192
rect 26056 9936 26108 9988
rect 26976 10047 27028 10056
rect 26976 10013 26985 10047
rect 26985 10013 27019 10047
rect 27019 10013 27028 10047
rect 26976 10004 27028 10013
rect 27068 10047 27120 10056
rect 27068 10013 27077 10047
rect 27077 10013 27111 10047
rect 27111 10013 27120 10047
rect 27068 10004 27120 10013
rect 26516 9936 26568 9988
rect 27252 10072 27304 10124
rect 27620 10072 27672 10124
rect 27988 10140 28040 10192
rect 29828 10140 29880 10192
rect 31208 10251 31260 10260
rect 31208 10217 31217 10251
rect 31217 10217 31251 10251
rect 31251 10217 31260 10251
rect 31208 10208 31260 10217
rect 31668 10208 31720 10260
rect 32864 10208 32916 10260
rect 34428 10251 34480 10260
rect 34428 10217 34437 10251
rect 34437 10217 34471 10251
rect 34471 10217 34480 10251
rect 34428 10208 34480 10217
rect 31300 10140 31352 10192
rect 31576 10140 31628 10192
rect 33876 10140 33928 10192
rect 27528 10047 27580 10056
rect 27528 10013 27537 10047
rect 27537 10013 27571 10047
rect 27571 10013 27580 10047
rect 27528 10004 27580 10013
rect 27712 10004 27764 10056
rect 28080 10047 28132 10056
rect 28080 10013 28089 10047
rect 28089 10013 28123 10047
rect 28123 10013 28132 10047
rect 28080 10004 28132 10013
rect 28356 10047 28408 10056
rect 28356 10013 28365 10047
rect 28365 10013 28399 10047
rect 28399 10013 28408 10047
rect 28356 10004 28408 10013
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28448 10004 28500 10013
rect 28724 10004 28776 10056
rect 29184 10072 29236 10124
rect 29276 10072 29328 10124
rect 29092 10004 29144 10056
rect 30196 10072 30248 10124
rect 31392 10115 31444 10124
rect 31392 10081 31401 10115
rect 31401 10081 31435 10115
rect 31435 10081 31444 10115
rect 31392 10072 31444 10081
rect 31024 10047 31076 10056
rect 31024 10013 31033 10047
rect 31033 10013 31067 10047
rect 31067 10013 31076 10047
rect 31024 10004 31076 10013
rect 31944 10072 31996 10124
rect 32404 10072 32456 10124
rect 27804 9911 27856 9920
rect 27804 9877 27813 9911
rect 27813 9877 27847 9911
rect 27847 9877 27856 9911
rect 27804 9868 27856 9877
rect 28632 9868 28684 9920
rect 28816 9936 28868 9988
rect 30472 9936 30524 9988
rect 28908 9868 28960 9920
rect 29736 9868 29788 9920
rect 30288 9868 30340 9920
rect 31760 10004 31812 10056
rect 32128 10004 32180 10056
rect 32772 10004 32824 10056
rect 35440 10072 35492 10124
rect 32496 9936 32548 9988
rect 33324 9936 33376 9988
rect 33876 10004 33928 10056
rect 34704 10047 34756 10056
rect 34704 10013 34713 10047
rect 34713 10013 34747 10047
rect 34747 10013 34756 10047
rect 34704 10004 34756 10013
rect 34796 9936 34848 9988
rect 35164 9936 35216 9988
rect 35992 9979 36044 9988
rect 35992 9945 36001 9979
rect 36001 9945 36035 9979
rect 36035 9945 36044 9979
rect 35992 9936 36044 9945
rect 31392 9868 31444 9920
rect 33140 9868 33192 9920
rect 34152 9911 34204 9920
rect 34152 9877 34161 9911
rect 34161 9877 34195 9911
rect 34195 9877 34204 9911
rect 34152 9868 34204 9877
rect 34336 9868 34388 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 3424 9664 3476 9716
rect 2320 9639 2372 9648
rect 2320 9605 2329 9639
rect 2329 9605 2363 9639
rect 2363 9605 2372 9639
rect 2320 9596 2372 9605
rect 2688 9639 2740 9648
rect 2688 9605 2697 9639
rect 2697 9605 2731 9639
rect 2731 9605 2740 9639
rect 2688 9596 2740 9605
rect 2412 9528 2464 9580
rect 4620 9596 4672 9648
rect 5632 9664 5684 9716
rect 7472 9596 7524 9648
rect 8484 9664 8536 9716
rect 8760 9664 8812 9716
rect 9312 9664 9364 9716
rect 7748 9596 7800 9648
rect 10876 9664 10928 9716
rect 12716 9664 12768 9716
rect 11980 9639 12032 9648
rect 4068 9528 4120 9580
rect 3056 9460 3108 9512
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 5264 9528 5316 9580
rect 5448 9571 5500 9580
rect 5448 9537 5454 9571
rect 5454 9537 5488 9571
rect 5488 9537 5500 9571
rect 5448 9528 5500 9537
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 6920 9571 6972 9580
rect 6920 9537 6924 9571
rect 6924 9537 6958 9571
rect 6958 9537 6972 9571
rect 6920 9528 6972 9537
rect 3976 9392 4028 9444
rect 4896 9392 4948 9444
rect 7012 9460 7064 9512
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 7472 9460 7524 9512
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 8208 9392 8260 9444
rect 4804 9324 4856 9376
rect 5172 9324 5224 9376
rect 5908 9324 5960 9376
rect 6644 9324 6696 9376
rect 6736 9367 6788 9376
rect 6736 9333 6745 9367
rect 6745 9333 6779 9367
rect 6779 9333 6788 9367
rect 6736 9324 6788 9333
rect 7748 9324 7800 9376
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 9036 9528 9088 9580
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 9864 9528 9916 9580
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 13360 9664 13412 9716
rect 14648 9664 14700 9716
rect 15016 9664 15068 9716
rect 19064 9664 19116 9716
rect 9588 9460 9640 9512
rect 10600 9460 10652 9512
rect 10968 9528 11020 9580
rect 11704 9528 11756 9580
rect 12900 9639 12952 9648
rect 12900 9605 12909 9639
rect 12909 9605 12943 9639
rect 12943 9605 12952 9639
rect 12900 9596 12952 9605
rect 9404 9392 9456 9444
rect 8576 9367 8628 9376
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 9128 9324 9180 9376
rect 10324 9324 10376 9376
rect 10876 9392 10928 9444
rect 11612 9392 11664 9444
rect 12532 9392 12584 9444
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 12716 9324 12768 9376
rect 13452 9528 13504 9580
rect 13912 9528 13964 9580
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 14832 9571 14884 9580
rect 14832 9537 14841 9571
rect 14841 9537 14875 9571
rect 14875 9537 14884 9571
rect 17868 9596 17920 9648
rect 20904 9664 20956 9716
rect 19432 9596 19484 9648
rect 14832 9528 14884 9537
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 13544 9392 13596 9444
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 15568 9460 15620 9512
rect 17684 9528 17736 9580
rect 18144 9528 18196 9580
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 22468 9664 22520 9716
rect 22560 9707 22612 9716
rect 22560 9673 22569 9707
rect 22569 9673 22603 9707
rect 22603 9673 22612 9707
rect 22560 9664 22612 9673
rect 23848 9664 23900 9716
rect 26332 9664 26384 9716
rect 27068 9664 27120 9716
rect 18052 9460 18104 9512
rect 19892 9460 19944 9512
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 23020 9596 23072 9648
rect 25228 9596 25280 9648
rect 20904 9392 20956 9444
rect 14188 9324 14240 9376
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 15200 9324 15252 9376
rect 15844 9324 15896 9376
rect 18052 9324 18104 9376
rect 22284 9392 22336 9444
rect 23388 9528 23440 9580
rect 23664 9528 23716 9580
rect 26056 9571 26108 9580
rect 26056 9537 26065 9571
rect 26065 9537 26099 9571
rect 26099 9537 26108 9571
rect 26056 9528 26108 9537
rect 26424 9639 26476 9648
rect 26424 9605 26433 9639
rect 26433 9605 26467 9639
rect 26467 9605 26476 9639
rect 26424 9596 26476 9605
rect 23204 9324 23256 9376
rect 23296 9324 23348 9376
rect 25872 9367 25924 9376
rect 25872 9333 25881 9367
rect 25881 9333 25915 9367
rect 25915 9333 25924 9367
rect 25872 9324 25924 9333
rect 26976 9571 27028 9580
rect 26976 9537 26985 9571
rect 26985 9537 27019 9571
rect 27019 9537 27028 9571
rect 26976 9528 27028 9537
rect 26792 9460 26844 9512
rect 28448 9664 28500 9716
rect 28540 9664 28592 9716
rect 31024 9664 31076 9716
rect 32220 9707 32272 9716
rect 32220 9673 32229 9707
rect 32229 9673 32263 9707
rect 32263 9673 32272 9707
rect 32220 9664 32272 9673
rect 34704 9664 34756 9716
rect 28356 9596 28408 9648
rect 31852 9596 31904 9648
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 27252 9571 27304 9580
rect 27252 9537 27261 9571
rect 27261 9537 27295 9571
rect 27295 9537 27304 9571
rect 27252 9528 27304 9537
rect 29828 9571 29880 9580
rect 29828 9537 29837 9571
rect 29837 9537 29871 9571
rect 29871 9537 29880 9571
rect 29828 9528 29880 9537
rect 30288 9528 30340 9580
rect 30472 9571 30524 9580
rect 30472 9537 30481 9571
rect 30481 9537 30515 9571
rect 30515 9537 30524 9571
rect 30472 9528 30524 9537
rect 31024 9528 31076 9580
rect 31392 9571 31444 9580
rect 31392 9537 31401 9571
rect 31401 9537 31435 9571
rect 31435 9537 31444 9571
rect 31392 9528 31444 9537
rect 31576 9571 31628 9580
rect 31576 9537 31585 9571
rect 31585 9537 31619 9571
rect 31619 9537 31628 9571
rect 31576 9528 31628 9537
rect 33692 9596 33744 9648
rect 33784 9639 33836 9648
rect 33784 9605 33793 9639
rect 33793 9605 33827 9639
rect 33827 9605 33836 9639
rect 33784 9596 33836 9605
rect 34428 9596 34480 9648
rect 35164 9596 35216 9648
rect 27528 9460 27580 9512
rect 28172 9460 28224 9512
rect 29552 9460 29604 9512
rect 31760 9503 31812 9512
rect 27068 9392 27120 9444
rect 27620 9392 27672 9444
rect 30932 9392 30984 9444
rect 27344 9324 27396 9376
rect 31760 9469 31769 9503
rect 31769 9469 31803 9503
rect 31803 9469 31812 9503
rect 31760 9460 31812 9469
rect 32404 9571 32456 9580
rect 32404 9537 32413 9571
rect 32413 9537 32447 9571
rect 32447 9537 32456 9571
rect 32404 9528 32456 9537
rect 33048 9528 33100 9580
rect 33508 9571 33560 9580
rect 33508 9537 33517 9571
rect 33517 9537 33551 9571
rect 33551 9537 33560 9571
rect 33508 9528 33560 9537
rect 35072 9528 35124 9580
rect 35348 9460 35400 9512
rect 35532 9571 35584 9580
rect 35532 9537 35541 9571
rect 35541 9537 35575 9571
rect 35575 9537 35584 9571
rect 35532 9528 35584 9537
rect 35624 9460 35676 9512
rect 35256 9392 35308 9444
rect 35440 9392 35492 9444
rect 35716 9392 35768 9444
rect 31392 9324 31444 9376
rect 32588 9324 32640 9376
rect 32772 9324 32824 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4344 9120 4396 9172
rect 6368 9120 6420 9172
rect 8300 9120 8352 9172
rect 10232 9120 10284 9172
rect 2504 9052 2556 9104
rect 4712 8984 4764 9036
rect 4896 8984 4948 9036
rect 6092 8984 6144 9036
rect 6276 8984 6328 9036
rect 6552 8984 6604 9036
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 5632 8916 5684 8968
rect 4620 8848 4672 8900
rect 4528 8780 4580 8832
rect 5356 8848 5408 8900
rect 5540 8848 5592 8900
rect 6000 8848 6052 8900
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 7104 8959 7156 8968
rect 7104 8925 7112 8959
rect 7112 8925 7146 8959
rect 7146 8925 7156 8959
rect 7104 8916 7156 8925
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 8760 9052 8812 9104
rect 8576 8984 8628 9036
rect 8484 8916 8536 8968
rect 8668 8916 8720 8968
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 10508 8984 10560 9036
rect 10968 9120 11020 9172
rect 11704 9163 11756 9172
rect 11704 9129 11713 9163
rect 11713 9129 11747 9163
rect 11747 9129 11756 9163
rect 11704 9120 11756 9129
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 22560 9120 22612 9172
rect 22928 9120 22980 9172
rect 23388 9120 23440 9172
rect 25872 9120 25924 9172
rect 12532 9052 12584 9104
rect 9496 8916 9548 8968
rect 12440 8984 12492 9036
rect 11612 8916 11664 8968
rect 14188 9052 14240 9104
rect 16580 9052 16632 9104
rect 17592 9095 17644 9104
rect 17592 9061 17601 9095
rect 17601 9061 17635 9095
rect 17635 9061 17644 9095
rect 17592 9052 17644 9061
rect 17776 9052 17828 9104
rect 19064 9052 19116 9104
rect 20996 9052 21048 9104
rect 17132 8984 17184 9036
rect 4988 8780 5040 8832
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 6368 8780 6420 8832
rect 6552 8780 6604 8832
rect 8116 8848 8168 8900
rect 11152 8848 11204 8900
rect 8760 8780 8812 8832
rect 9312 8780 9364 8832
rect 10048 8780 10100 8832
rect 10232 8780 10284 8832
rect 11980 8780 12032 8832
rect 12624 8823 12676 8832
rect 12624 8789 12633 8823
rect 12633 8789 12667 8823
rect 12667 8789 12676 8823
rect 12624 8780 12676 8789
rect 12808 8780 12860 8832
rect 17040 8959 17092 8968
rect 17040 8925 17049 8959
rect 17049 8925 17083 8959
rect 17083 8925 17092 8959
rect 17040 8916 17092 8925
rect 17776 8959 17828 8968
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 18144 8959 18196 8968
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 19340 8984 19392 9036
rect 19708 8984 19760 9036
rect 20076 9027 20128 9036
rect 20076 8993 20085 9027
rect 20085 8993 20119 9027
rect 20119 8993 20128 9027
rect 20076 8984 20128 8993
rect 20260 9027 20312 9036
rect 20260 8993 20269 9027
rect 20269 8993 20303 9027
rect 20303 8993 20312 9027
rect 20260 8984 20312 8993
rect 18236 8848 18288 8900
rect 18788 8959 18840 8968
rect 18788 8925 18797 8959
rect 18797 8925 18831 8959
rect 18831 8925 18840 8959
rect 18788 8916 18840 8925
rect 18972 8959 19024 8968
rect 18972 8925 18981 8959
rect 18981 8925 19015 8959
rect 19015 8925 19024 8959
rect 18972 8916 19024 8925
rect 23112 8984 23164 9036
rect 25044 9052 25096 9104
rect 28356 9052 28408 9104
rect 27804 8984 27856 9036
rect 29368 9120 29420 9172
rect 30748 9163 30800 9172
rect 30748 9129 30757 9163
rect 30757 9129 30791 9163
rect 30791 9129 30800 9163
rect 30748 9120 30800 9129
rect 31484 9120 31536 9172
rect 32680 9120 32732 9172
rect 29092 9052 29144 9104
rect 30472 9052 30524 9104
rect 31944 9052 31996 9104
rect 36360 9120 36412 9172
rect 19248 8848 19300 8900
rect 20352 8848 20404 8900
rect 20536 8916 20588 8968
rect 23296 8916 23348 8968
rect 23388 8959 23440 8968
rect 23388 8925 23397 8959
rect 23397 8925 23431 8959
rect 23431 8925 23440 8959
rect 23388 8916 23440 8925
rect 23664 8959 23716 8968
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 18328 8780 18380 8832
rect 18512 8780 18564 8832
rect 19064 8780 19116 8832
rect 23112 8780 23164 8832
rect 23296 8780 23348 8832
rect 23572 8848 23624 8900
rect 26700 8891 26752 8900
rect 26700 8857 26709 8891
rect 26709 8857 26743 8891
rect 26743 8857 26752 8891
rect 26700 8848 26752 8857
rect 27068 8916 27120 8968
rect 27344 8916 27396 8968
rect 27620 8848 27672 8900
rect 25320 8780 25372 8832
rect 29092 8916 29144 8968
rect 29368 8959 29420 8968
rect 29368 8925 29377 8959
rect 29377 8925 29411 8959
rect 29411 8925 29420 8959
rect 29368 8916 29420 8925
rect 29828 8848 29880 8900
rect 31944 8916 31996 8968
rect 32404 8916 32456 8968
rect 33968 8984 34020 9036
rect 34244 9095 34296 9104
rect 34244 9061 34253 9095
rect 34253 9061 34287 9095
rect 34287 9061 34296 9095
rect 34244 9052 34296 9061
rect 34428 9052 34480 9104
rect 35716 9052 35768 9104
rect 34612 8984 34664 9036
rect 35072 8984 35124 9036
rect 32036 8848 32088 8900
rect 34152 8848 34204 8900
rect 34244 8848 34296 8900
rect 35164 8916 35216 8968
rect 35440 8916 35492 8968
rect 35624 8848 35676 8900
rect 29092 8823 29144 8832
rect 29092 8789 29101 8823
rect 29101 8789 29135 8823
rect 29135 8789 29144 8823
rect 29092 8780 29144 8789
rect 29460 8780 29512 8832
rect 29920 8780 29972 8832
rect 30104 8780 30156 8832
rect 33232 8780 33284 8832
rect 34336 8780 34388 8832
rect 34888 8780 34940 8832
rect 35532 8780 35584 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 4344 8576 4396 8628
rect 4620 8576 4672 8628
rect 5264 8576 5316 8628
rect 5356 8576 5408 8628
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 4896 8551 4948 8560
rect 4896 8517 4905 8551
rect 4905 8517 4939 8551
rect 4939 8517 4948 8551
rect 4896 8508 4948 8517
rect 1400 8440 1452 8492
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 4436 8440 4488 8492
rect 4528 8440 4580 8492
rect 5080 8440 5132 8492
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 4896 8372 4948 8424
rect 5448 8440 5500 8492
rect 6276 8508 6328 8560
rect 6552 8440 6604 8492
rect 6736 8440 6788 8492
rect 8024 8576 8076 8628
rect 8668 8576 8720 8628
rect 9220 8576 9272 8628
rect 10048 8576 10100 8628
rect 10416 8576 10468 8628
rect 11336 8576 11388 8628
rect 7748 8551 7800 8560
rect 7748 8517 7757 8551
rect 7757 8517 7791 8551
rect 7791 8517 7800 8551
rect 7748 8508 7800 8517
rect 8484 8551 8536 8560
rect 8484 8517 8493 8551
rect 8493 8517 8527 8551
rect 8527 8517 8536 8551
rect 8484 8508 8536 8517
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 7472 8440 7524 8492
rect 6092 8372 6144 8424
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 9312 8440 9364 8492
rect 5448 8304 5500 8356
rect 3884 8236 3936 8288
rect 5080 8236 5132 8288
rect 5908 8236 5960 8288
rect 7012 8304 7064 8356
rect 8944 8415 8996 8424
rect 8944 8381 8953 8415
rect 8953 8381 8987 8415
rect 8987 8381 8996 8415
rect 8944 8372 8996 8381
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10968 8508 11020 8560
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 10876 8440 10928 8492
rect 12164 8576 12216 8628
rect 12624 8576 12676 8628
rect 16120 8576 16172 8628
rect 10232 8304 10284 8356
rect 11612 8440 11664 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 13176 8508 13228 8560
rect 18144 8508 18196 8560
rect 14464 8440 14516 8492
rect 12808 8304 12860 8356
rect 13176 8304 13228 8356
rect 16672 8372 16724 8424
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 17316 8440 17368 8492
rect 17408 8440 17460 8492
rect 17592 8440 17644 8492
rect 17960 8440 18012 8492
rect 18788 8576 18840 8628
rect 19800 8576 19852 8628
rect 21548 8576 21600 8628
rect 23480 8576 23532 8628
rect 23756 8576 23808 8628
rect 24768 8576 24820 8628
rect 25412 8576 25464 8628
rect 26608 8576 26660 8628
rect 33048 8576 33100 8628
rect 33508 8576 33560 8628
rect 36084 8576 36136 8628
rect 18328 8551 18380 8560
rect 18328 8517 18337 8551
rect 18337 8517 18371 8551
rect 18371 8517 18380 8551
rect 18328 8508 18380 8517
rect 18512 8508 18564 8560
rect 29092 8508 29144 8560
rect 19064 8440 19116 8492
rect 20260 8440 20312 8492
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 17040 8372 17092 8424
rect 7196 8279 7248 8288
rect 7196 8245 7205 8279
rect 7205 8245 7239 8279
rect 7239 8245 7248 8279
rect 7196 8236 7248 8245
rect 8852 8236 8904 8288
rect 10784 8279 10836 8288
rect 10784 8245 10793 8279
rect 10793 8245 10827 8279
rect 10827 8245 10836 8279
rect 10784 8236 10836 8245
rect 11428 8236 11480 8288
rect 11612 8236 11664 8288
rect 11888 8236 11940 8288
rect 14280 8236 14332 8288
rect 16764 8304 16816 8356
rect 15936 8236 15988 8288
rect 18972 8372 19024 8424
rect 20720 8372 20772 8424
rect 21548 8372 21600 8424
rect 23296 8440 23348 8492
rect 20352 8236 20404 8288
rect 23204 8372 23256 8424
rect 23112 8304 23164 8356
rect 25412 8440 25464 8492
rect 23572 8415 23624 8424
rect 23572 8381 23581 8415
rect 23581 8381 23615 8415
rect 23615 8381 23624 8415
rect 23572 8372 23624 8381
rect 23756 8372 23808 8424
rect 23848 8372 23900 8424
rect 26148 8483 26200 8492
rect 26148 8449 26157 8483
rect 26157 8449 26191 8483
rect 26191 8449 26200 8483
rect 26148 8440 26200 8449
rect 26700 8440 26752 8492
rect 30104 8508 30156 8560
rect 30932 8508 30984 8560
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 29828 8483 29880 8492
rect 29828 8449 29837 8483
rect 29837 8449 29871 8483
rect 29871 8449 29880 8483
rect 29828 8440 29880 8449
rect 30380 8483 30432 8492
rect 30380 8449 30389 8483
rect 30389 8449 30423 8483
rect 30423 8449 30432 8483
rect 30380 8440 30432 8449
rect 25688 8372 25740 8424
rect 26056 8372 26108 8424
rect 30288 8372 30340 8424
rect 31852 8440 31904 8492
rect 32864 8483 32916 8492
rect 32864 8449 32873 8483
rect 32873 8449 32907 8483
rect 32907 8449 32916 8483
rect 32864 8440 32916 8449
rect 32772 8372 32824 8424
rect 32956 8372 33008 8424
rect 33968 8440 34020 8492
rect 34152 8483 34204 8492
rect 34152 8449 34161 8483
rect 34161 8449 34195 8483
rect 34195 8449 34204 8483
rect 34152 8440 34204 8449
rect 34428 8440 34480 8492
rect 34520 8372 34572 8424
rect 35072 8372 35124 8424
rect 23296 8236 23348 8288
rect 25688 8279 25740 8288
rect 25688 8245 25697 8279
rect 25697 8245 25731 8279
rect 25731 8245 25740 8279
rect 25688 8236 25740 8245
rect 25780 8236 25832 8288
rect 30104 8236 30156 8288
rect 34612 8236 34664 8288
rect 35164 8236 35216 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3516 8032 3568 8084
rect 4620 7964 4672 8016
rect 5448 8032 5500 8084
rect 7656 8032 7708 8084
rect 9036 8032 9088 8084
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 10784 8032 10836 8084
rect 13268 8032 13320 8084
rect 14372 8032 14424 8084
rect 15384 8032 15436 8084
rect 22100 8032 22152 8084
rect 23112 8075 23164 8084
rect 23112 8041 23121 8075
rect 23121 8041 23155 8075
rect 23155 8041 23164 8075
rect 23112 8032 23164 8041
rect 23296 8075 23348 8084
rect 23296 8041 23305 8075
rect 23305 8041 23339 8075
rect 23339 8041 23348 8075
rect 23296 8032 23348 8041
rect 23572 8032 23624 8084
rect 24400 8032 24452 8084
rect 6552 7964 6604 8016
rect 5908 7896 5960 7948
rect 6644 7896 6696 7948
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 4896 7760 4948 7812
rect 6276 7828 6328 7880
rect 6736 7828 6788 7880
rect 13820 7964 13872 8016
rect 8668 7896 8720 7948
rect 8760 7896 8812 7948
rect 9404 7896 9456 7948
rect 9496 7896 9548 7948
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 12716 7896 12768 7948
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 7748 7828 7800 7880
rect 10140 7828 10192 7880
rect 10232 7828 10284 7880
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 14740 7896 14792 7948
rect 14188 7828 14240 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 24308 7964 24360 8016
rect 17040 7896 17092 7948
rect 17316 7896 17368 7948
rect 20260 7896 20312 7948
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 4804 7692 4856 7744
rect 5080 7692 5132 7744
rect 5540 7692 5592 7744
rect 7012 7803 7064 7812
rect 7012 7769 7021 7803
rect 7021 7769 7055 7803
rect 7055 7769 7064 7803
rect 7012 7760 7064 7769
rect 7932 7760 7984 7812
rect 8392 7803 8444 7812
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 8668 7760 8720 7812
rect 10784 7760 10836 7812
rect 11152 7760 11204 7812
rect 6276 7692 6328 7744
rect 7288 7692 7340 7744
rect 8116 7692 8168 7744
rect 10324 7692 10376 7744
rect 13820 7760 13872 7812
rect 15108 7871 15160 7880
rect 15108 7837 15117 7871
rect 15117 7837 15151 7871
rect 15151 7837 15160 7871
rect 15108 7828 15160 7837
rect 15384 7828 15436 7880
rect 15936 7828 15988 7880
rect 19064 7828 19116 7880
rect 19340 7828 19392 7880
rect 20628 7828 20680 7880
rect 21916 7896 21968 7948
rect 22100 7896 22152 7948
rect 21088 7871 21140 7880
rect 21088 7837 21097 7871
rect 21097 7837 21131 7871
rect 21131 7837 21140 7871
rect 21088 7828 21140 7837
rect 21180 7828 21232 7880
rect 22928 7828 22980 7880
rect 23756 7896 23808 7948
rect 24584 7939 24636 7948
rect 24584 7905 24593 7939
rect 24593 7905 24627 7939
rect 24627 7905 24636 7939
rect 24584 7896 24636 7905
rect 25688 8032 25740 8084
rect 26976 8075 27028 8084
rect 26976 8041 26985 8075
rect 26985 8041 27019 8075
rect 27019 8041 27028 8075
rect 26976 8032 27028 8041
rect 27252 8032 27304 8084
rect 29828 8075 29880 8084
rect 29828 8041 29837 8075
rect 29837 8041 29871 8075
rect 29871 8041 29880 8075
rect 29828 8032 29880 8041
rect 30104 8075 30156 8084
rect 30104 8041 30113 8075
rect 30113 8041 30147 8075
rect 30147 8041 30156 8075
rect 30104 8032 30156 8041
rect 33876 8032 33928 8084
rect 35348 8075 35400 8084
rect 35348 8041 35357 8075
rect 35357 8041 35391 8075
rect 35391 8041 35400 8075
rect 35348 8032 35400 8041
rect 26148 7964 26200 8016
rect 23480 7871 23532 7880
rect 23480 7837 23489 7871
rect 23489 7837 23523 7871
rect 23523 7837 23532 7871
rect 23480 7828 23532 7837
rect 12900 7692 12952 7744
rect 13360 7692 13412 7744
rect 15568 7803 15620 7812
rect 15568 7769 15577 7803
rect 15577 7769 15611 7803
rect 15611 7769 15620 7803
rect 15568 7760 15620 7769
rect 15752 7803 15804 7812
rect 15752 7769 15761 7803
rect 15761 7769 15795 7803
rect 15795 7769 15804 7803
rect 15752 7760 15804 7769
rect 16948 7760 17000 7812
rect 18696 7760 18748 7812
rect 19248 7760 19300 7812
rect 19708 7760 19760 7812
rect 20536 7692 20588 7744
rect 20720 7692 20772 7744
rect 22468 7692 22520 7744
rect 23020 7692 23072 7744
rect 24676 7871 24728 7880
rect 24676 7837 24685 7871
rect 24685 7837 24719 7871
rect 24719 7837 24728 7871
rect 24676 7828 24728 7837
rect 25320 7871 25372 7880
rect 25320 7837 25329 7871
rect 25329 7837 25363 7871
rect 25363 7837 25372 7871
rect 25320 7828 25372 7837
rect 25504 7871 25556 7880
rect 25504 7837 25513 7871
rect 25513 7837 25547 7871
rect 25547 7837 25556 7871
rect 25504 7828 25556 7837
rect 25688 7871 25740 7880
rect 25688 7837 25697 7871
rect 25697 7837 25731 7871
rect 25731 7837 25740 7871
rect 25688 7828 25740 7837
rect 25780 7871 25832 7880
rect 25780 7837 25789 7871
rect 25789 7837 25823 7871
rect 25823 7837 25832 7871
rect 25780 7828 25832 7837
rect 26976 7896 27028 7948
rect 27804 7939 27856 7948
rect 27804 7905 27813 7939
rect 27813 7905 27847 7939
rect 27847 7905 27856 7939
rect 27804 7896 27856 7905
rect 26056 7871 26108 7880
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 25228 7760 25280 7812
rect 25412 7803 25464 7812
rect 25412 7769 25421 7803
rect 25421 7769 25455 7803
rect 25455 7769 25464 7803
rect 25412 7760 25464 7769
rect 24860 7692 24912 7744
rect 24952 7735 25004 7744
rect 24952 7701 24961 7735
rect 24961 7701 24995 7735
rect 24995 7701 25004 7735
rect 24952 7692 25004 7701
rect 25044 7692 25096 7744
rect 26516 7828 26568 7880
rect 27252 7828 27304 7880
rect 26608 7760 26660 7812
rect 27896 7871 27948 7880
rect 27896 7837 27905 7871
rect 27905 7837 27939 7871
rect 27939 7837 27948 7871
rect 27896 7828 27948 7837
rect 26792 7692 26844 7744
rect 28540 7939 28592 7948
rect 28540 7905 28549 7939
rect 28549 7905 28583 7939
rect 28583 7905 28592 7939
rect 28540 7896 28592 7905
rect 30288 7964 30340 8016
rect 30380 7964 30432 8016
rect 32220 7964 32272 8016
rect 34796 7964 34848 8016
rect 30840 7896 30892 7948
rect 35440 7896 35492 7948
rect 28724 7871 28776 7880
rect 28724 7837 28733 7871
rect 28733 7837 28767 7871
rect 28767 7837 28776 7871
rect 28724 7828 28776 7837
rect 29828 7760 29880 7812
rect 30932 7871 30984 7880
rect 30932 7837 30941 7871
rect 30941 7837 30975 7871
rect 30975 7837 30984 7871
rect 30932 7828 30984 7837
rect 32864 7828 32916 7880
rect 33416 7828 33468 7880
rect 31024 7760 31076 7812
rect 31852 7760 31904 7812
rect 29276 7692 29328 7744
rect 30656 7735 30708 7744
rect 30656 7701 30665 7735
rect 30665 7701 30699 7735
rect 30699 7701 30708 7735
rect 30656 7692 30708 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 4344 7488 4396 7540
rect 4620 7488 4672 7540
rect 5264 7488 5316 7540
rect 5816 7488 5868 7540
rect 6736 7488 6788 7540
rect 7472 7488 7524 7540
rect 8944 7488 8996 7540
rect 2964 7420 3016 7472
rect 7012 7420 7064 7472
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 5264 7352 5316 7404
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 4804 7284 4856 7336
rect 5172 7284 5224 7336
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 8392 7420 8444 7472
rect 8760 7463 8812 7472
rect 8760 7429 8769 7463
rect 8769 7429 8803 7463
rect 8803 7429 8812 7463
rect 8760 7420 8812 7429
rect 8852 7463 8904 7472
rect 8852 7429 8861 7463
rect 8861 7429 8895 7463
rect 8895 7429 8904 7463
rect 8852 7420 8904 7429
rect 9404 7420 9456 7472
rect 10508 7488 10560 7540
rect 10876 7488 10928 7540
rect 9772 7420 9824 7472
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 6000 7284 6052 7336
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 6000 7148 6052 7200
rect 7932 7284 7984 7336
rect 9588 7352 9640 7404
rect 10048 7352 10100 7404
rect 10324 7420 10376 7472
rect 12716 7488 12768 7540
rect 6644 7259 6696 7268
rect 6644 7225 6653 7259
rect 6653 7225 6687 7259
rect 6687 7225 6696 7259
rect 6644 7216 6696 7225
rect 8576 7216 8628 7268
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 12624 7420 12676 7472
rect 12900 7420 12952 7472
rect 13452 7488 13504 7540
rect 14188 7488 14240 7540
rect 15752 7488 15804 7540
rect 16672 7531 16724 7540
rect 16672 7497 16681 7531
rect 16681 7497 16715 7531
rect 16715 7497 16724 7531
rect 16672 7488 16724 7497
rect 18144 7531 18196 7540
rect 18144 7497 18153 7531
rect 18153 7497 18187 7531
rect 18187 7497 18196 7531
rect 18144 7488 18196 7497
rect 18604 7488 18656 7540
rect 18880 7488 18932 7540
rect 14556 7420 14608 7472
rect 14740 7463 14792 7472
rect 14740 7429 14749 7463
rect 14749 7429 14783 7463
rect 14783 7429 14792 7463
rect 14740 7420 14792 7429
rect 15200 7420 15252 7472
rect 11428 7352 11480 7404
rect 11612 7395 11664 7404
rect 11612 7361 11621 7395
rect 11621 7361 11655 7395
rect 11655 7361 11664 7395
rect 11612 7352 11664 7361
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 12256 7352 12308 7404
rect 14280 7352 14332 7404
rect 11796 7284 11848 7336
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 8208 7148 8260 7200
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 10232 7148 10284 7200
rect 10324 7148 10376 7200
rect 11704 7148 11756 7200
rect 12072 7148 12124 7200
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 12716 7284 12768 7336
rect 14648 7284 14700 7336
rect 16488 7352 16540 7404
rect 17316 7420 17368 7472
rect 18052 7420 18104 7472
rect 17132 7395 17184 7404
rect 17132 7361 17141 7395
rect 17141 7361 17175 7395
rect 17175 7361 17184 7395
rect 17132 7352 17184 7361
rect 18236 7352 18288 7404
rect 19524 7488 19576 7540
rect 19432 7420 19484 7472
rect 19708 7463 19760 7472
rect 19708 7429 19717 7463
rect 19717 7429 19751 7463
rect 19751 7429 19760 7463
rect 19708 7420 19760 7429
rect 20444 7488 20496 7540
rect 20536 7488 20588 7540
rect 19156 7352 19208 7404
rect 19248 7352 19300 7404
rect 21088 7420 21140 7472
rect 21916 7420 21968 7472
rect 17224 7284 17276 7336
rect 20628 7352 20680 7404
rect 20720 7352 20772 7404
rect 21640 7395 21692 7404
rect 21640 7361 21649 7395
rect 21649 7361 21683 7395
rect 21683 7361 21692 7395
rect 21640 7352 21692 7361
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 22376 7352 22428 7404
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 19156 7216 19208 7268
rect 12256 7191 12308 7200
rect 12256 7157 12265 7191
rect 12265 7157 12299 7191
rect 12299 7157 12308 7191
rect 12256 7148 12308 7157
rect 15384 7148 15436 7200
rect 16580 7148 16632 7200
rect 20720 7216 20772 7268
rect 19892 7191 19944 7200
rect 19892 7157 19901 7191
rect 19901 7157 19935 7191
rect 19935 7157 19944 7191
rect 19892 7148 19944 7157
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 22100 7259 22152 7268
rect 22100 7225 22109 7259
rect 22109 7225 22143 7259
rect 22143 7225 22152 7259
rect 22100 7216 22152 7225
rect 22836 7395 22888 7404
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 24952 7488 25004 7540
rect 26240 7488 26292 7540
rect 27436 7488 27488 7540
rect 27896 7488 27948 7540
rect 30932 7488 30984 7540
rect 31300 7488 31352 7540
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 25044 7420 25096 7472
rect 25688 7420 25740 7472
rect 25228 7352 25280 7404
rect 25596 7352 25648 7404
rect 26148 7352 26200 7404
rect 28080 7420 28132 7472
rect 27896 7395 27948 7404
rect 27896 7361 27905 7395
rect 27905 7361 27939 7395
rect 27939 7361 27948 7395
rect 27896 7352 27948 7361
rect 30840 7352 30892 7404
rect 23664 7216 23716 7268
rect 24952 7259 25004 7268
rect 24952 7225 24961 7259
rect 24961 7225 24995 7259
rect 24995 7225 25004 7259
rect 24952 7216 25004 7225
rect 25412 7284 25464 7336
rect 25688 7327 25740 7336
rect 25688 7293 25697 7327
rect 25697 7293 25731 7327
rect 25731 7293 25740 7327
rect 25688 7284 25740 7293
rect 26976 7284 27028 7336
rect 22652 7191 22704 7200
rect 22652 7157 22661 7191
rect 22661 7157 22695 7191
rect 22695 7157 22704 7191
rect 22652 7148 22704 7157
rect 23480 7148 23532 7200
rect 30656 7216 30708 7268
rect 25504 7148 25556 7200
rect 26516 7148 26568 7200
rect 27068 7148 27120 7200
rect 27528 7148 27580 7200
rect 30840 7148 30892 7200
rect 31392 7395 31444 7404
rect 31392 7361 31401 7395
rect 31401 7361 31435 7395
rect 31435 7361 31444 7395
rect 31392 7352 31444 7361
rect 33048 7463 33100 7472
rect 33048 7429 33057 7463
rect 33057 7429 33091 7463
rect 33091 7429 33100 7463
rect 33048 7420 33100 7429
rect 31852 7395 31904 7404
rect 31852 7361 31861 7395
rect 31861 7361 31895 7395
rect 31895 7361 31904 7395
rect 31852 7352 31904 7361
rect 32864 7395 32916 7404
rect 32864 7361 32873 7395
rect 32873 7361 32907 7395
rect 32907 7361 32916 7395
rect 32864 7352 32916 7361
rect 31668 7216 31720 7268
rect 31484 7148 31536 7200
rect 32496 7148 32548 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2964 6944 3016 6996
rect 3976 6944 4028 6996
rect 4620 6944 4672 6996
rect 4804 6944 4856 6996
rect 5172 6944 5224 6996
rect 4712 6876 4764 6928
rect 5908 6944 5960 6996
rect 3516 6740 3568 6792
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 4436 6740 4488 6792
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 4252 6672 4304 6724
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 6736 6876 6788 6928
rect 8576 6987 8628 6996
rect 8576 6953 8585 6987
rect 8585 6953 8619 6987
rect 8619 6953 8628 6987
rect 8576 6944 8628 6953
rect 9956 6944 10008 6996
rect 10416 6944 10468 6996
rect 8208 6876 8260 6928
rect 11060 6944 11112 6996
rect 12624 6944 12676 6996
rect 13360 6987 13412 6996
rect 13360 6953 13369 6987
rect 13369 6953 13403 6987
rect 13403 6953 13412 6987
rect 13360 6944 13412 6953
rect 13820 6944 13872 6996
rect 17224 6944 17276 6996
rect 17868 6944 17920 6996
rect 19892 6944 19944 6996
rect 20720 6944 20772 6996
rect 21640 6944 21692 6996
rect 22100 6944 22152 6996
rect 25320 6944 25372 6996
rect 25872 6944 25924 6996
rect 26424 6944 26476 6996
rect 5448 6672 5500 6724
rect 5908 6715 5960 6724
rect 5908 6681 5917 6715
rect 5917 6681 5951 6715
rect 5951 6681 5960 6715
rect 5908 6672 5960 6681
rect 6276 6740 6328 6792
rect 6552 6740 6604 6792
rect 7472 6740 7524 6792
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 8392 6808 8444 6860
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 13544 6876 13596 6928
rect 10324 6808 10376 6860
rect 10416 6808 10468 6860
rect 10968 6808 11020 6860
rect 11520 6851 11572 6860
rect 11520 6817 11529 6851
rect 11529 6817 11563 6851
rect 11563 6817 11572 6851
rect 11520 6808 11572 6817
rect 8852 6740 8904 6792
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 11060 6740 11112 6792
rect 6552 6604 6604 6656
rect 7196 6604 7248 6656
rect 7472 6604 7524 6656
rect 8484 6604 8536 6656
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 9956 6604 10008 6656
rect 10232 6672 10284 6724
rect 11244 6672 11296 6724
rect 11888 6672 11940 6724
rect 12164 6740 12216 6792
rect 13820 6808 13872 6860
rect 12992 6740 13044 6792
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 17132 6808 17184 6860
rect 17316 6808 17368 6860
rect 17868 6808 17920 6860
rect 20076 6876 20128 6928
rect 24216 6876 24268 6928
rect 25780 6876 25832 6928
rect 27528 6987 27580 6996
rect 27528 6953 27537 6987
rect 27537 6953 27571 6987
rect 27571 6953 27580 6987
rect 27528 6944 27580 6953
rect 32864 6944 32916 6996
rect 28816 6876 28868 6928
rect 18604 6851 18656 6860
rect 18604 6817 18613 6851
rect 18613 6817 18647 6851
rect 18647 6817 18656 6851
rect 18604 6808 18656 6817
rect 12440 6672 12492 6724
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 18880 6808 18932 6860
rect 22008 6808 22060 6860
rect 24124 6808 24176 6860
rect 25872 6808 25924 6860
rect 26332 6808 26384 6860
rect 17224 6672 17276 6724
rect 10416 6604 10468 6656
rect 11152 6604 11204 6656
rect 13360 6604 13412 6656
rect 13912 6604 13964 6656
rect 14648 6604 14700 6656
rect 18052 6672 18104 6724
rect 18236 6672 18288 6724
rect 18880 6672 18932 6724
rect 19708 6783 19760 6792
rect 19708 6749 19717 6783
rect 19717 6749 19751 6783
rect 19751 6749 19760 6783
rect 19708 6740 19760 6749
rect 20444 6740 20496 6792
rect 20536 6740 20588 6792
rect 18696 6604 18748 6656
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 21456 6672 21508 6724
rect 22928 6672 22980 6724
rect 26884 6715 26936 6724
rect 26884 6681 26893 6715
rect 26893 6681 26927 6715
rect 26927 6681 26936 6715
rect 26884 6672 26936 6681
rect 19616 6604 19668 6656
rect 20812 6604 20864 6656
rect 21548 6604 21600 6656
rect 25412 6604 25464 6656
rect 26240 6604 26292 6656
rect 27068 6647 27120 6656
rect 27068 6613 27098 6647
rect 27098 6613 27120 6647
rect 27068 6604 27120 6613
rect 27252 6647 27304 6656
rect 27252 6613 27261 6647
rect 27261 6613 27295 6647
rect 27295 6613 27304 6647
rect 27252 6604 27304 6613
rect 27344 6647 27396 6656
rect 27344 6613 27353 6647
rect 27353 6613 27387 6647
rect 27387 6613 27396 6647
rect 27344 6604 27396 6613
rect 29920 6851 29972 6860
rect 29920 6817 29929 6851
rect 29929 6817 29963 6851
rect 29963 6817 29972 6851
rect 29920 6808 29972 6817
rect 32496 6808 32548 6860
rect 33876 6808 33928 6860
rect 29828 6783 29880 6792
rect 29828 6749 29837 6783
rect 29837 6749 29871 6783
rect 29871 6749 29880 6783
rect 29828 6740 29880 6749
rect 32864 6740 32916 6792
rect 27620 6672 27672 6724
rect 31392 6672 31444 6724
rect 33416 6740 33468 6792
rect 34796 6876 34848 6928
rect 29092 6604 29144 6656
rect 30564 6604 30616 6656
rect 31668 6604 31720 6656
rect 33876 6604 33928 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 4344 6443 4396 6452
rect 4344 6409 4353 6443
rect 4353 6409 4387 6443
rect 4387 6409 4396 6443
rect 4344 6400 4396 6409
rect 5264 6400 5316 6452
rect 5356 6443 5408 6452
rect 5356 6409 5365 6443
rect 5365 6409 5399 6443
rect 5399 6409 5408 6443
rect 5356 6400 5408 6409
rect 5540 6400 5592 6452
rect 5908 6400 5960 6452
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 6184 6400 6236 6452
rect 6828 6400 6880 6452
rect 7656 6400 7708 6452
rect 8760 6443 8812 6452
rect 8760 6409 8769 6443
rect 8769 6409 8803 6443
rect 8803 6409 8812 6443
rect 8760 6400 8812 6409
rect 9956 6400 10008 6452
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 4344 6264 4396 6316
rect 4620 6264 4672 6316
rect 4896 6264 4948 6316
rect 7196 6332 7248 6384
rect 7748 6332 7800 6384
rect 9772 6332 9824 6384
rect 11520 6400 11572 6452
rect 13176 6400 13228 6452
rect 13544 6443 13596 6452
rect 13544 6409 13553 6443
rect 13553 6409 13587 6443
rect 13587 6409 13596 6443
rect 13544 6400 13596 6409
rect 13636 6400 13688 6452
rect 14096 6443 14148 6452
rect 14096 6409 14105 6443
rect 14105 6409 14139 6443
rect 14139 6409 14148 6443
rect 14096 6400 14148 6409
rect 12072 6332 12124 6384
rect 17316 6400 17368 6452
rect 17408 6400 17460 6452
rect 17684 6400 17736 6452
rect 5264 6196 5316 6248
rect 5632 6239 5684 6248
rect 5632 6205 5641 6239
rect 5641 6205 5675 6239
rect 5675 6205 5684 6239
rect 5632 6196 5684 6205
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 6276 6264 6328 6316
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 8668 6196 8720 6248
rect 9496 6264 9548 6316
rect 11612 6264 11664 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 10876 6196 10928 6248
rect 12440 6264 12492 6316
rect 9588 6128 9640 6180
rect 10968 6128 11020 6180
rect 4896 6060 4948 6112
rect 5448 6060 5500 6112
rect 7380 6060 7432 6112
rect 9404 6060 9456 6112
rect 10048 6060 10100 6112
rect 11520 6060 11572 6112
rect 12716 6196 12768 6248
rect 12900 6196 12952 6248
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 15108 6332 15160 6384
rect 13728 6196 13780 6248
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 16212 6332 16264 6384
rect 16948 6332 17000 6384
rect 18328 6400 18380 6452
rect 19616 6400 19668 6452
rect 20536 6400 20588 6452
rect 21456 6400 21508 6452
rect 21640 6400 21692 6452
rect 23756 6400 23808 6452
rect 24676 6400 24728 6452
rect 25872 6443 25924 6452
rect 25872 6409 25881 6443
rect 25881 6409 25915 6443
rect 25915 6409 25924 6443
rect 25872 6400 25924 6409
rect 15660 6264 15712 6316
rect 17868 6264 17920 6316
rect 16304 6196 16356 6248
rect 17132 6196 17184 6248
rect 18236 6196 18288 6248
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 19340 6332 19392 6384
rect 21088 6332 21140 6384
rect 21548 6332 21600 6384
rect 21824 6332 21876 6384
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 19708 6264 19760 6316
rect 20904 6264 20956 6316
rect 23112 6264 23164 6316
rect 24032 6375 24084 6384
rect 24032 6341 24041 6375
rect 24041 6341 24075 6375
rect 24075 6341 24084 6375
rect 24032 6332 24084 6341
rect 24124 6264 24176 6316
rect 25044 6332 25096 6384
rect 26056 6375 26108 6384
rect 26056 6341 26065 6375
rect 26065 6341 26099 6375
rect 26099 6341 26108 6375
rect 26056 6332 26108 6341
rect 27252 6332 27304 6384
rect 24676 6307 24728 6316
rect 24676 6273 24691 6307
rect 24691 6273 24725 6307
rect 24725 6273 24728 6307
rect 24676 6264 24728 6273
rect 12348 6128 12400 6180
rect 13912 6128 13964 6180
rect 15752 6128 15804 6180
rect 15844 6128 15896 6180
rect 22744 6196 22796 6248
rect 25504 6307 25556 6316
rect 25504 6273 25513 6307
rect 25513 6273 25547 6307
rect 25547 6273 25556 6307
rect 25504 6264 25556 6273
rect 25596 6264 25648 6316
rect 27344 6307 27396 6316
rect 27344 6273 27353 6307
rect 27353 6273 27387 6307
rect 27387 6273 27396 6307
rect 27344 6264 27396 6273
rect 28816 6400 28868 6452
rect 30932 6400 30984 6452
rect 33324 6443 33376 6452
rect 33324 6409 33333 6443
rect 33333 6409 33367 6443
rect 33367 6409 33376 6443
rect 33324 6400 33376 6409
rect 33876 6400 33928 6452
rect 30104 6332 30156 6384
rect 31668 6332 31720 6384
rect 32312 6375 32364 6384
rect 32312 6341 32321 6375
rect 32321 6341 32355 6375
rect 32355 6341 32364 6375
rect 32312 6332 32364 6341
rect 25412 6196 25464 6248
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 15292 6060 15344 6112
rect 15384 6103 15436 6112
rect 15384 6069 15393 6103
rect 15393 6069 15427 6103
rect 15427 6069 15436 6103
rect 15384 6060 15436 6069
rect 15476 6060 15528 6112
rect 18972 6060 19024 6112
rect 20720 6060 20772 6112
rect 21640 6060 21692 6112
rect 22376 6060 22428 6112
rect 24584 6060 24636 6112
rect 24676 6060 24728 6112
rect 26148 6128 26200 6180
rect 26792 6128 26844 6180
rect 28632 6264 28684 6316
rect 28908 6196 28960 6248
rect 29736 6264 29788 6316
rect 30288 6264 30340 6316
rect 30564 6307 30616 6316
rect 30564 6273 30573 6307
rect 30573 6273 30607 6307
rect 30607 6273 30616 6307
rect 30564 6264 30616 6273
rect 30840 6307 30892 6316
rect 30840 6273 30849 6307
rect 30849 6273 30883 6307
rect 30883 6273 30892 6307
rect 30840 6264 30892 6273
rect 30932 6264 30984 6316
rect 31392 6264 31444 6316
rect 29920 6196 29972 6248
rect 30748 6196 30800 6248
rect 32220 6196 32272 6248
rect 32864 6264 32916 6316
rect 33416 6264 33468 6316
rect 34612 6264 34664 6316
rect 29644 6128 29696 6180
rect 31484 6128 31536 6180
rect 34244 6128 34296 6180
rect 25688 6060 25740 6112
rect 26240 6103 26292 6112
rect 26240 6069 26249 6103
rect 26249 6069 26283 6103
rect 26283 6069 26292 6103
rect 26240 6060 26292 6069
rect 26516 6060 26568 6112
rect 28356 6060 28408 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5264 5899 5316 5908
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 5264 5856 5316 5865
rect 7288 5856 7340 5908
rect 10784 5856 10836 5908
rect 12440 5856 12492 5908
rect 16212 5899 16264 5908
rect 16212 5865 16221 5899
rect 16221 5865 16255 5899
rect 16255 5865 16264 5899
rect 16212 5856 16264 5865
rect 16304 5856 16356 5908
rect 20720 5856 20772 5908
rect 20904 5856 20956 5908
rect 21272 5856 21324 5908
rect 8116 5788 8168 5840
rect 5632 5720 5684 5772
rect 7104 5720 7156 5772
rect 5356 5695 5408 5704
rect 5356 5661 5365 5695
rect 5365 5661 5399 5695
rect 5399 5661 5408 5695
rect 5356 5652 5408 5661
rect 6368 5652 6420 5704
rect 9588 5763 9640 5772
rect 9588 5729 9597 5763
rect 9597 5729 9631 5763
rect 9631 5729 9640 5763
rect 9588 5720 9640 5729
rect 9956 5788 10008 5840
rect 13912 5788 13964 5840
rect 22560 5788 22612 5840
rect 22744 5856 22796 5908
rect 24584 5856 24636 5908
rect 25504 5856 25556 5908
rect 26792 5788 26844 5840
rect 30380 5856 30432 5908
rect 30564 5856 30616 5908
rect 31944 5899 31996 5908
rect 31944 5865 31953 5899
rect 31953 5865 31987 5899
rect 31987 5865 31996 5899
rect 31944 5856 31996 5865
rect 11796 5763 11848 5772
rect 11796 5729 11805 5763
rect 11805 5729 11839 5763
rect 11839 5729 11848 5763
rect 11796 5720 11848 5729
rect 12716 5720 12768 5772
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 10048 5584 10100 5636
rect 10876 5584 10928 5636
rect 11336 5584 11388 5636
rect 11612 5584 11664 5636
rect 12532 5584 12584 5636
rect 19248 5720 19300 5772
rect 14004 5652 14056 5704
rect 14740 5652 14792 5704
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 15660 5652 15712 5704
rect 16396 5652 16448 5704
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 8392 5516 8444 5568
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 9312 5516 9364 5568
rect 10784 5516 10836 5568
rect 15844 5584 15896 5636
rect 19432 5652 19484 5704
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 14556 5516 14608 5568
rect 15568 5516 15620 5568
rect 17408 5584 17460 5636
rect 17960 5584 18012 5636
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 19708 5695 19760 5704
rect 19708 5661 19717 5695
rect 19717 5661 19751 5695
rect 19751 5661 19760 5695
rect 19708 5652 19760 5661
rect 19984 5652 20036 5704
rect 20260 5652 20312 5704
rect 24676 5763 24728 5772
rect 24676 5729 24685 5763
rect 24685 5729 24719 5763
rect 24719 5729 24728 5763
rect 24676 5720 24728 5729
rect 18052 5516 18104 5568
rect 19340 5516 19392 5568
rect 19524 5516 19576 5568
rect 20720 5584 20772 5636
rect 21548 5695 21600 5704
rect 21548 5661 21557 5695
rect 21557 5661 21591 5695
rect 21591 5661 21600 5695
rect 21548 5652 21600 5661
rect 21640 5695 21692 5704
rect 21640 5661 21649 5695
rect 21649 5661 21683 5695
rect 21683 5661 21692 5695
rect 21640 5652 21692 5661
rect 21824 5695 21876 5704
rect 21824 5661 21833 5695
rect 21833 5661 21867 5695
rect 21867 5661 21876 5695
rect 21824 5652 21876 5661
rect 22836 5695 22888 5704
rect 22836 5661 22845 5695
rect 22845 5661 22879 5695
rect 22879 5661 22888 5695
rect 22836 5652 22888 5661
rect 23572 5652 23624 5704
rect 23756 5695 23808 5704
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 24584 5652 24636 5704
rect 25044 5720 25096 5772
rect 27252 5788 27304 5840
rect 27988 5788 28040 5840
rect 26148 5652 26200 5704
rect 23940 5516 23992 5568
rect 26332 5516 26384 5568
rect 26976 5695 27028 5704
rect 26976 5661 26985 5695
rect 26985 5661 27019 5695
rect 27019 5661 27028 5695
rect 26976 5652 27028 5661
rect 28908 5720 28960 5772
rect 27988 5695 28040 5704
rect 27988 5661 27997 5695
rect 27997 5661 28031 5695
rect 28031 5661 28040 5695
rect 27988 5652 28040 5661
rect 28356 5627 28408 5636
rect 28356 5593 28374 5627
rect 28374 5593 28408 5627
rect 28356 5584 28408 5593
rect 29736 5720 29788 5772
rect 30196 5788 30248 5840
rect 30656 5831 30708 5840
rect 30656 5797 30665 5831
rect 30665 5797 30699 5831
rect 30699 5797 30708 5831
rect 30656 5788 30708 5797
rect 30840 5788 30892 5840
rect 29644 5695 29696 5704
rect 29644 5661 29653 5695
rect 29653 5661 29687 5695
rect 29687 5661 29696 5695
rect 29644 5652 29696 5661
rect 30932 5763 30984 5772
rect 30932 5729 30941 5763
rect 30941 5729 30975 5763
rect 30975 5729 30984 5763
rect 30932 5720 30984 5729
rect 31484 5831 31536 5840
rect 31484 5797 31493 5831
rect 31493 5797 31527 5831
rect 31527 5797 31536 5831
rect 31484 5788 31536 5797
rect 30564 5652 30616 5704
rect 30104 5584 30156 5636
rect 27344 5516 27396 5568
rect 28172 5559 28224 5568
rect 28172 5525 28181 5559
rect 28181 5525 28215 5559
rect 28215 5525 28224 5559
rect 28172 5516 28224 5525
rect 29552 5516 29604 5568
rect 32128 5720 32180 5772
rect 32220 5695 32272 5704
rect 32220 5661 32229 5695
rect 32229 5661 32263 5695
rect 32263 5661 32272 5695
rect 32220 5652 32272 5661
rect 32864 5695 32916 5704
rect 32864 5661 32873 5695
rect 32873 5661 32907 5695
rect 32907 5661 32916 5695
rect 32864 5652 32916 5661
rect 33876 5652 33928 5704
rect 33416 5584 33468 5636
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 8116 5355 8168 5364
rect 8116 5321 8125 5355
rect 8125 5321 8159 5355
rect 8159 5321 8168 5355
rect 8116 5312 8168 5321
rect 7748 5244 7800 5296
rect 9312 5244 9364 5296
rect 11704 5312 11756 5364
rect 11796 5312 11848 5364
rect 11060 5287 11112 5296
rect 11060 5253 11069 5287
rect 11069 5253 11103 5287
rect 11103 5253 11112 5287
rect 11060 5244 11112 5253
rect 11244 5244 11296 5296
rect 10140 5176 10192 5228
rect 10232 5108 10284 5160
rect 9864 5040 9916 5092
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 11428 5176 11480 5228
rect 11888 5244 11940 5296
rect 12808 5244 12860 5296
rect 13084 5244 13136 5296
rect 14188 5244 14240 5296
rect 19156 5312 19208 5364
rect 22008 5312 22060 5364
rect 14372 5244 14424 5296
rect 15660 5244 15712 5296
rect 19248 5244 19300 5296
rect 18512 5176 18564 5228
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 11244 5108 11296 5160
rect 11888 5108 11940 5160
rect 13820 5108 13872 5160
rect 15016 5151 15068 5160
rect 15016 5117 15025 5151
rect 15025 5117 15059 5151
rect 15059 5117 15068 5151
rect 15016 5108 15068 5117
rect 15292 5108 15344 5160
rect 21732 5244 21784 5296
rect 24308 5312 24360 5364
rect 21180 5176 21232 5228
rect 22192 5219 22244 5228
rect 22192 5185 22201 5219
rect 22201 5185 22235 5219
rect 22235 5185 22244 5219
rect 22192 5176 22244 5185
rect 22468 5176 22520 5228
rect 24032 5176 24084 5228
rect 26884 5176 26936 5228
rect 27436 5176 27488 5228
rect 29828 5176 29880 5228
rect 30656 5176 30708 5228
rect 10784 4972 10836 5024
rect 11796 4972 11848 5024
rect 11888 4972 11940 5024
rect 13912 5040 13964 5092
rect 20168 5040 20220 5092
rect 21088 5040 21140 5092
rect 21640 5040 21692 5092
rect 30380 5083 30432 5092
rect 30380 5049 30389 5083
rect 30389 5049 30423 5083
rect 30423 5049 30432 5083
rect 30380 5040 30432 5049
rect 12992 4972 13044 5024
rect 13544 4972 13596 5024
rect 14372 5015 14424 5024
rect 14372 4981 14381 5015
rect 14381 4981 14415 5015
rect 14415 4981 14424 5015
rect 14372 4972 14424 4981
rect 19340 4972 19392 5024
rect 19708 5015 19760 5024
rect 19708 4981 19717 5015
rect 19717 4981 19751 5015
rect 19751 4981 19760 5015
rect 19708 4972 19760 4981
rect 22560 4972 22612 5024
rect 26976 5015 27028 5024
rect 26976 4981 26985 5015
rect 26985 4981 27019 5015
rect 27019 4981 27028 5015
rect 26976 4972 27028 4981
rect 27344 5015 27396 5024
rect 27344 4981 27353 5015
rect 27353 4981 27387 5015
rect 27387 4981 27396 5015
rect 27344 4972 27396 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 11244 4768 11296 4820
rect 11612 4768 11664 4820
rect 9956 4632 10008 4684
rect 11336 4700 11388 4752
rect 11888 4700 11940 4752
rect 11152 4632 11204 4684
rect 11244 4632 11296 4684
rect 12164 4632 12216 4684
rect 12348 4632 12400 4684
rect 8024 4564 8076 4616
rect 11704 4564 11756 4616
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 12072 4564 12124 4616
rect 15292 4768 15344 4820
rect 15660 4768 15712 4820
rect 17408 4768 17460 4820
rect 14372 4700 14424 4752
rect 15936 4700 15988 4752
rect 17500 4743 17552 4752
rect 13360 4675 13412 4684
rect 13360 4641 13369 4675
rect 13369 4641 13403 4675
rect 13403 4641 13412 4675
rect 13360 4632 13412 4641
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 15752 4632 15804 4684
rect 9864 4496 9916 4548
rect 10140 4496 10192 4548
rect 10968 4496 11020 4548
rect 11796 4428 11848 4480
rect 11980 4428 12032 4480
rect 12348 4471 12400 4480
rect 12348 4437 12357 4471
rect 12357 4437 12391 4471
rect 12391 4437 12400 4471
rect 12348 4428 12400 4437
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 15844 4564 15896 4616
rect 16028 4607 16080 4616
rect 16028 4573 16037 4607
rect 16037 4573 16071 4607
rect 16071 4573 16080 4607
rect 16028 4564 16080 4573
rect 17500 4709 17509 4743
rect 17509 4709 17543 4743
rect 17543 4709 17552 4743
rect 17500 4700 17552 4709
rect 18236 4700 18288 4752
rect 18512 4811 18564 4820
rect 18512 4777 18521 4811
rect 18521 4777 18555 4811
rect 18555 4777 18564 4811
rect 18512 4768 18564 4777
rect 20720 4768 20772 4820
rect 21088 4768 21140 4820
rect 22192 4768 22244 4820
rect 23112 4768 23164 4820
rect 24400 4768 24452 4820
rect 25412 4768 25464 4820
rect 34520 4768 34572 4820
rect 21272 4700 21324 4752
rect 21364 4700 21416 4752
rect 21732 4700 21784 4752
rect 17040 4632 17092 4684
rect 16120 4496 16172 4548
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 22652 4675 22704 4684
rect 22652 4641 22661 4675
rect 22661 4641 22695 4675
rect 22695 4641 22704 4675
rect 22652 4632 22704 4641
rect 18420 4564 18472 4616
rect 21640 4607 21692 4616
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 21824 4607 21876 4616
rect 21824 4573 21833 4607
rect 21833 4573 21867 4607
rect 21867 4573 21876 4607
rect 21824 4564 21876 4573
rect 22284 4607 22336 4616
rect 22284 4573 22293 4607
rect 22293 4573 22327 4607
rect 22327 4573 22336 4607
rect 22284 4564 22336 4573
rect 23940 4564 23992 4616
rect 16856 4496 16908 4548
rect 16212 4428 16264 4480
rect 17408 4496 17460 4548
rect 17684 4471 17736 4480
rect 17684 4437 17693 4471
rect 17693 4437 17727 4471
rect 17727 4437 17736 4471
rect 17684 4428 17736 4437
rect 18052 4496 18104 4548
rect 21364 4496 21416 4548
rect 23848 4539 23900 4548
rect 23848 4505 23857 4539
rect 23857 4505 23891 4539
rect 23891 4505 23900 4539
rect 23848 4496 23900 4505
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 9772 4224 9824 4276
rect 10784 4224 10836 4276
rect 13636 4224 13688 4276
rect 16028 4224 16080 4276
rect 18420 4267 18472 4276
rect 18420 4233 18429 4267
rect 18429 4233 18463 4267
rect 18463 4233 18472 4267
rect 18420 4224 18472 4233
rect 9680 4156 9732 4208
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 8852 4063 8904 4072
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 9220 4020 9272 4072
rect 9588 4020 9640 4072
rect 11060 4088 11112 4140
rect 11244 4020 11296 4072
rect 12164 4156 12216 4208
rect 12716 4156 12768 4208
rect 13452 4156 13504 4208
rect 14372 4156 14424 4208
rect 11704 4088 11756 4140
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 15844 4131 15896 4140
rect 15844 4097 15853 4131
rect 15853 4097 15887 4131
rect 15887 4097 15896 4131
rect 15844 4088 15896 4097
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16212 4088 16264 4140
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 12808 4020 12860 4072
rect 14464 4020 14516 4072
rect 15384 4020 15436 4072
rect 15660 4020 15712 4072
rect 16396 4020 16448 4072
rect 16488 4020 16540 4072
rect 17132 4020 17184 4072
rect 17684 4020 17736 4072
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 20996 4088 21048 4140
rect 21088 4131 21140 4140
rect 21088 4097 21097 4131
rect 21097 4097 21131 4131
rect 21131 4097 21140 4131
rect 21088 4088 21140 4097
rect 21364 4131 21416 4140
rect 21364 4097 21373 4131
rect 21373 4097 21407 4131
rect 21407 4097 21416 4131
rect 21364 4088 21416 4097
rect 21456 4131 21508 4140
rect 21456 4097 21465 4131
rect 21465 4097 21499 4131
rect 21499 4097 21508 4131
rect 21456 4088 21508 4097
rect 24308 4199 24360 4208
rect 24308 4165 24317 4199
rect 24317 4165 24351 4199
rect 24351 4165 24360 4199
rect 24308 4156 24360 4165
rect 24400 4199 24452 4208
rect 24400 4165 24409 4199
rect 24409 4165 24443 4199
rect 24443 4165 24452 4199
rect 24400 4156 24452 4165
rect 18604 3952 18656 4004
rect 21548 4020 21600 4072
rect 23572 4088 23624 4140
rect 24124 4131 24176 4140
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 24124 4088 24176 4097
rect 21456 3952 21508 4004
rect 22192 4063 22244 4072
rect 22192 4029 22201 4063
rect 22201 4029 22235 4063
rect 22235 4029 22244 4063
rect 22192 4020 22244 4029
rect 25320 4131 25372 4140
rect 25320 4097 25329 4131
rect 25329 4097 25363 4131
rect 25363 4097 25372 4131
rect 25320 4088 25372 4097
rect 26056 4088 26108 4140
rect 28632 4131 28684 4140
rect 28632 4097 28641 4131
rect 28641 4097 28675 4131
rect 28675 4097 28684 4131
rect 28632 4088 28684 4097
rect 29092 4088 29144 4140
rect 8300 3884 8352 3936
rect 10140 3884 10192 3936
rect 10876 3884 10928 3936
rect 13452 3884 13504 3936
rect 14832 3884 14884 3936
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 15752 3884 15804 3936
rect 16212 3884 16264 3936
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 17408 3884 17460 3936
rect 18788 3927 18840 3936
rect 18788 3893 18797 3927
rect 18797 3893 18831 3927
rect 18831 3893 18840 3927
rect 18788 3884 18840 3893
rect 21272 3884 21324 3936
rect 21916 3884 21968 3936
rect 22468 3884 22520 3936
rect 23940 3927 23992 3936
rect 23940 3893 23949 3927
rect 23949 3893 23983 3927
rect 23983 3893 23992 3927
rect 23940 3884 23992 3893
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 27436 3952 27488 4004
rect 26884 3884 26936 3936
rect 27068 3884 27120 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 8852 3680 8904 3732
rect 9128 3680 9180 3732
rect 9772 3612 9824 3664
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 8484 3544 8536 3596
rect 10784 3544 10836 3596
rect 10876 3587 10928 3596
rect 10876 3553 10885 3587
rect 10885 3553 10919 3587
rect 10919 3553 10928 3587
rect 10876 3544 10928 3553
rect 11704 3680 11756 3732
rect 11796 3680 11848 3732
rect 12900 3680 12952 3732
rect 14464 3680 14516 3732
rect 15292 3723 15344 3732
rect 15292 3689 15301 3723
rect 15301 3689 15335 3723
rect 15335 3689 15344 3723
rect 15292 3680 15344 3689
rect 16120 3680 16172 3732
rect 19524 3680 19576 3732
rect 20628 3680 20680 3732
rect 14004 3612 14056 3664
rect 14188 3612 14240 3664
rect 11244 3544 11296 3596
rect 11428 3587 11480 3596
rect 11428 3553 11437 3587
rect 11437 3553 11471 3587
rect 11471 3553 11480 3587
rect 11428 3544 11480 3553
rect 8116 3408 8168 3460
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 9220 3476 9272 3528
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 12716 3476 12768 3528
rect 13360 3544 13412 3596
rect 13728 3544 13780 3596
rect 17592 3612 17644 3664
rect 21088 3612 21140 3664
rect 22192 3612 22244 3664
rect 24032 3723 24084 3732
rect 24032 3689 24041 3723
rect 24041 3689 24075 3723
rect 24075 3689 24084 3723
rect 24032 3680 24084 3689
rect 27436 3723 27488 3732
rect 27436 3689 27445 3723
rect 27445 3689 27479 3723
rect 27479 3689 27488 3723
rect 27436 3680 27488 3689
rect 35992 3680 36044 3732
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 15016 3544 15068 3596
rect 12992 3476 13044 3528
rect 13452 3476 13504 3528
rect 15384 3476 15436 3528
rect 15844 3544 15896 3596
rect 16028 3544 16080 3596
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 18236 3587 18288 3596
rect 18236 3553 18245 3587
rect 18245 3553 18279 3587
rect 18279 3553 18288 3587
rect 18236 3544 18288 3553
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 21180 3544 21232 3596
rect 21456 3544 21508 3596
rect 26976 3612 27028 3664
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 9864 3408 9916 3460
rect 11612 3340 11664 3392
rect 14188 3408 14240 3460
rect 13268 3340 13320 3392
rect 15108 3340 15160 3392
rect 18604 3408 18656 3460
rect 19524 3408 19576 3460
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 21088 3519 21140 3528
rect 21088 3485 21097 3519
rect 21097 3485 21131 3519
rect 21131 3485 21140 3519
rect 21088 3476 21140 3485
rect 21272 3519 21324 3528
rect 21272 3485 21281 3519
rect 21281 3485 21315 3519
rect 21315 3485 21324 3519
rect 21272 3476 21324 3485
rect 21824 3519 21876 3528
rect 21824 3485 21833 3519
rect 21833 3485 21867 3519
rect 21867 3485 21876 3519
rect 21824 3476 21876 3485
rect 22560 3587 22612 3596
rect 22560 3553 22569 3587
rect 22569 3553 22603 3587
rect 22603 3553 22612 3587
rect 22560 3544 22612 3553
rect 23848 3544 23900 3596
rect 24676 3544 24728 3596
rect 28264 3544 28316 3596
rect 17500 3340 17552 3392
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 23572 3476 23624 3528
rect 22284 3408 22336 3460
rect 22100 3340 22152 3392
rect 22652 3340 22704 3392
rect 26148 3519 26200 3528
rect 26148 3485 26157 3519
rect 26157 3485 26191 3519
rect 26191 3485 26200 3519
rect 26148 3476 26200 3485
rect 26884 3476 26936 3528
rect 27528 3519 27580 3528
rect 27528 3485 27537 3519
rect 27537 3485 27571 3519
rect 27571 3485 27580 3519
rect 27528 3476 27580 3485
rect 29000 3476 29052 3528
rect 36084 3519 36136 3528
rect 36084 3485 36093 3519
rect 36093 3485 36127 3519
rect 36127 3485 36136 3519
rect 36084 3476 36136 3485
rect 25412 3408 25464 3460
rect 27068 3340 27120 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 8760 3136 8812 3188
rect 9036 3111 9088 3120
rect 9036 3077 9045 3111
rect 9045 3077 9079 3111
rect 9079 3077 9088 3111
rect 9036 3068 9088 3077
rect 12992 3136 13044 3188
rect 12348 3068 12400 3120
rect 13268 3068 13320 3120
rect 13820 3068 13872 3120
rect 8300 3000 8352 3052
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 9864 3000 9916 3052
rect 11244 3043 11296 3052
rect 11244 3009 11253 3043
rect 11253 3009 11287 3043
rect 11287 3009 11296 3043
rect 11244 3000 11296 3009
rect 12440 3000 12492 3052
rect 15108 3068 15160 3120
rect 15660 3068 15712 3120
rect 16028 3136 16080 3188
rect 16396 3179 16448 3188
rect 16396 3145 16405 3179
rect 16405 3145 16439 3179
rect 16439 3145 16448 3179
rect 16396 3136 16448 3145
rect 18420 3136 18472 3188
rect 18788 3136 18840 3188
rect 16672 3068 16724 3120
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 16212 3043 16264 3052
rect 16212 3009 16221 3043
rect 16221 3009 16255 3043
rect 16255 3009 16264 3043
rect 16212 3000 16264 3009
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 16396 3000 16448 3052
rect 17592 3068 17644 3120
rect 20444 3111 20496 3120
rect 20444 3077 20453 3111
rect 20453 3077 20487 3111
rect 20487 3077 20496 3111
rect 20444 3068 20496 3077
rect 22100 3136 22152 3188
rect 8484 2932 8536 2984
rect 9220 2932 9272 2984
rect 9312 2932 9364 2984
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 14280 2932 14332 2984
rect 18604 3000 18656 3052
rect 8668 2864 8720 2916
rect 16488 2864 16540 2916
rect 17132 2907 17184 2916
rect 17132 2873 17141 2907
rect 17141 2873 17175 2907
rect 17175 2873 17184 2907
rect 17132 2864 17184 2873
rect 8392 2796 8444 2848
rect 8944 2796 8996 2848
rect 9220 2796 9272 2848
rect 12256 2796 12308 2848
rect 14556 2796 14608 2848
rect 17500 2975 17552 2984
rect 17500 2941 17509 2975
rect 17509 2941 17543 2975
rect 17543 2941 17552 2975
rect 17500 2932 17552 2941
rect 17868 2932 17920 2984
rect 19984 3000 20036 3052
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 22192 3068 22244 3120
rect 23572 3068 23624 3120
rect 34060 3068 34112 3120
rect 26148 3000 26200 3052
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 21824 2864 21876 2916
rect 17684 2796 17736 2848
rect 19064 2839 19116 2848
rect 19064 2805 19073 2839
rect 19073 2805 19107 2839
rect 19107 2805 19116 2839
rect 19064 2796 19116 2805
rect 20720 2796 20772 2848
rect 21272 2839 21324 2848
rect 21272 2805 21281 2839
rect 21281 2805 21315 2839
rect 21315 2805 21324 2839
rect 21272 2796 21324 2805
rect 22560 2796 22612 2848
rect 23572 2839 23624 2848
rect 23572 2805 23581 2839
rect 23581 2805 23615 2839
rect 23615 2805 23624 2839
rect 23572 2796 23624 2805
rect 23664 2839 23716 2848
rect 23664 2805 23673 2839
rect 23673 2805 23707 2839
rect 23707 2805 23716 2839
rect 23664 2796 23716 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 10324 2592 10376 2644
rect 10784 2592 10836 2644
rect 12440 2592 12492 2644
rect 13728 2592 13780 2644
rect 14832 2592 14884 2644
rect 16304 2524 16356 2576
rect 8300 2456 8352 2508
rect 11244 2456 11296 2508
rect 11888 2456 11940 2508
rect 13820 2456 13872 2508
rect 8024 2431 8076 2440
rect 8024 2397 8033 2431
rect 8033 2397 8067 2431
rect 8067 2397 8076 2431
rect 8024 2388 8076 2397
rect 8576 2388 8628 2440
rect 10232 2388 10284 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 13544 2431 13596 2440
rect 13544 2397 13553 2431
rect 13553 2397 13587 2431
rect 13587 2397 13596 2431
rect 13544 2388 13596 2397
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 14004 2388 14056 2440
rect 18972 2592 19024 2644
rect 25136 2592 25188 2644
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 19064 2456 19116 2508
rect 22100 2456 22152 2508
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 21916 2388 21968 2440
rect 22652 2388 22704 2440
rect 23572 2456 23624 2508
rect 23664 2456 23716 2508
rect 9128 2320 9180 2372
rect 9220 2363 9272 2372
rect 9220 2329 9229 2363
rect 9229 2329 9263 2363
rect 9263 2329 9272 2363
rect 9220 2320 9272 2329
rect 9864 2320 9916 2372
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 12532 2320 12584 2372
rect 14372 2320 14424 2372
rect 15200 2320 15252 2372
rect 12164 2252 12216 2304
rect 14188 2252 14240 2304
rect 15476 2252 15528 2304
rect 15568 2252 15620 2304
rect 17408 2320 17460 2372
rect 16488 2252 16540 2304
rect 17868 2252 17920 2304
rect 20628 2252 20680 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 8208 2048 8260 2100
rect 11612 2048 11664 2100
<< metal2 >>
rect 22558 38926 22614 39726
rect 23202 38926 23258 39726
rect 23846 38926 23902 39726
rect 24490 38926 24546 39726
rect 25134 38926 25190 39726
rect 25778 38926 25834 39726
rect 26422 38926 26478 39726
rect 27066 38926 27122 39726
rect 28998 38926 29054 39726
rect 29642 38926 29698 39726
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 16948 37256 17000 37262
rect 16948 37198 17000 37204
rect 17040 37256 17092 37262
rect 17040 37198 17092 37204
rect 16580 37188 16632 37194
rect 16580 37130 16632 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 16120 36916 16172 36922
rect 16120 36858 16172 36864
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 8944 36304 8996 36310
rect 8944 36246 8996 36252
rect 8300 36236 8352 36242
rect 8300 36178 8352 36184
rect 6000 36168 6052 36174
rect 6000 36110 6052 36116
rect 7840 36168 7892 36174
rect 7840 36110 7892 36116
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 3698 35456 3754 35465
rect 3698 35391 3754 35400
rect 3332 32904 3384 32910
rect 3332 32846 3384 32852
rect 2964 32836 3016 32842
rect 2964 32778 3016 32784
rect 1306 32736 1362 32745
rect 1306 32671 1362 32680
rect 1320 32502 1348 32671
rect 1308 32496 1360 32502
rect 1308 32438 1360 32444
rect 1320 31890 1348 32438
rect 2504 32360 2556 32366
rect 2504 32302 2556 32308
rect 2410 32056 2466 32065
rect 2516 32026 2544 32302
rect 2596 32224 2648 32230
rect 2596 32166 2648 32172
rect 2410 31991 2466 32000
rect 2504 32020 2556 32026
rect 2424 31958 2452 31991
rect 2504 31962 2556 31968
rect 2412 31952 2464 31958
rect 2412 31894 2464 31900
rect 1308 31884 1360 31890
rect 1308 31826 1360 31832
rect 2424 31414 2452 31894
rect 2608 31822 2636 32166
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 1308 31408 1360 31414
rect 1306 31376 1308 31385
rect 2412 31408 2464 31414
rect 1360 31376 1362 31385
rect 2412 31350 2464 31356
rect 1306 31311 1362 31320
rect 1320 30598 1348 31311
rect 2792 31278 2820 31758
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2976 31210 3004 32778
rect 3344 31822 3372 32846
rect 3332 31816 3384 31822
rect 3332 31758 3384 31764
rect 3712 31754 3740 35391
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 6012 35290 6040 36110
rect 7104 36032 7156 36038
rect 7104 35974 7156 35980
rect 6736 35624 6788 35630
rect 6736 35566 6788 35572
rect 6748 35290 6776 35566
rect 6828 35488 6880 35494
rect 6828 35430 6880 35436
rect 6000 35284 6052 35290
rect 6000 35226 6052 35232
rect 6736 35284 6788 35290
rect 6736 35226 6788 35232
rect 6840 35154 6868 35430
rect 6828 35148 6880 35154
rect 6828 35090 6880 35096
rect 7116 35086 7144 35974
rect 7656 35556 7708 35562
rect 7656 35498 7708 35504
rect 7380 35216 7432 35222
rect 7380 35158 7432 35164
rect 6092 35080 6144 35086
rect 6092 35022 6144 35028
rect 6276 35080 6328 35086
rect 6276 35022 6328 35028
rect 6368 35080 6420 35086
rect 6368 35022 6420 35028
rect 6460 35080 6512 35086
rect 6460 35022 6512 35028
rect 7104 35080 7156 35086
rect 7104 35022 7156 35028
rect 7288 35080 7340 35086
rect 7288 35022 7340 35028
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 6104 34746 6132 35022
rect 6288 34746 6316 35022
rect 6092 34740 6144 34746
rect 6092 34682 6144 34688
rect 6276 34740 6328 34746
rect 6276 34682 6328 34688
rect 6184 34604 6236 34610
rect 6184 34546 6236 34552
rect 5448 34536 5500 34542
rect 5448 34478 5500 34484
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 5356 34060 5408 34066
rect 5356 34002 5408 34008
rect 4712 33992 4764 33998
rect 4712 33934 4764 33940
rect 4620 33856 4672 33862
rect 4620 33798 4672 33804
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4436 33040 4488 33046
rect 4436 32982 4488 32988
rect 4342 32872 4398 32881
rect 4342 32807 4344 32816
rect 4396 32807 4398 32816
rect 4344 32778 4396 32784
rect 4448 32502 4476 32982
rect 4632 32570 4660 33798
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 4436 32496 4488 32502
rect 4632 32450 4660 32506
rect 4436 32438 4488 32444
rect 4540 32422 4660 32450
rect 4724 32434 4752 33934
rect 5264 33924 5316 33930
rect 5264 33866 5316 33872
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 5276 33658 5304 33866
rect 5264 33652 5316 33658
rect 5264 33594 5316 33600
rect 5368 33522 5396 34002
rect 5356 33516 5408 33522
rect 5356 33458 5408 33464
rect 5264 33380 5316 33386
rect 5264 33322 5316 33328
rect 5276 33114 5304 33322
rect 5080 33108 5132 33114
rect 5080 33050 5132 33056
rect 5264 33108 5316 33114
rect 5264 33050 5316 33056
rect 4802 33008 4858 33017
rect 4802 32943 4804 32952
rect 4856 32943 4858 32952
rect 4804 32914 4856 32920
rect 5092 32910 5120 33050
rect 5172 33040 5224 33046
rect 5170 33008 5172 33017
rect 5224 33008 5226 33017
rect 5170 32943 5226 32952
rect 5460 32910 5488 34478
rect 5540 34196 5592 34202
rect 5540 34138 5592 34144
rect 6000 34196 6052 34202
rect 6000 34138 6052 34144
rect 5552 33590 5580 34138
rect 5540 33584 5592 33590
rect 5540 33526 5592 33532
rect 5540 33448 5592 33454
rect 5540 33390 5592 33396
rect 5552 33114 5580 33390
rect 5540 33108 5592 33114
rect 5540 33050 5592 33056
rect 5080 32904 5132 32910
rect 5080 32846 5132 32852
rect 5264 32904 5316 32910
rect 5264 32846 5316 32852
rect 5448 32904 5500 32910
rect 5448 32846 5500 32852
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 5092 32774 5120 32846
rect 4804 32768 4856 32774
rect 4804 32710 4856 32716
rect 5080 32768 5132 32774
rect 5080 32710 5132 32716
rect 4816 32434 4844 32710
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 5276 32570 5304 32846
rect 5264 32564 5316 32570
rect 5264 32506 5316 32512
rect 4986 32464 5042 32473
rect 4712 32428 4764 32434
rect 4540 32298 4568 32422
rect 4712 32370 4764 32376
rect 4804 32428 4856 32434
rect 4986 32399 5042 32408
rect 5264 32428 5316 32434
rect 4804 32370 4856 32376
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4528 32292 4580 32298
rect 4528 32234 4580 32240
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4160 32020 4212 32026
rect 4436 32020 4488 32026
rect 4160 31962 4212 31968
rect 4356 31980 4436 32008
rect 3712 31726 3832 31754
rect 3700 31680 3752 31686
rect 3700 31622 3752 31628
rect 2964 31204 3016 31210
rect 2964 31146 3016 31152
rect 1768 31136 1820 31142
rect 1768 31078 1820 31084
rect 1780 30666 1808 31078
rect 3148 30864 3200 30870
rect 3148 30806 3200 30812
rect 3160 30705 3188 30806
rect 3712 30802 3740 31622
rect 3700 30796 3752 30802
rect 3700 30738 3752 30744
rect 3240 30728 3292 30734
rect 3146 30696 3202 30705
rect 1768 30660 1820 30666
rect 1768 30602 1820 30608
rect 3056 30660 3108 30666
rect 3240 30670 3292 30676
rect 3146 30631 3202 30640
rect 3056 30602 3108 30608
rect 1308 30592 1360 30598
rect 1308 30534 1360 30540
rect 3068 30394 3096 30602
rect 3056 30388 3108 30394
rect 3056 30330 3108 30336
rect 1308 30184 1360 30190
rect 1308 30126 1360 30132
rect 1320 30025 1348 30126
rect 1306 30016 1362 30025
rect 1306 29951 1362 29960
rect 1320 29850 1348 29951
rect 1308 29844 1360 29850
rect 1308 29786 1360 29792
rect 3068 29510 3096 30330
rect 3160 29714 3188 30631
rect 3252 29714 3280 30670
rect 3712 30258 3740 30738
rect 3700 30252 3752 30258
rect 3700 30194 3752 30200
rect 3608 30116 3660 30122
rect 3608 30058 3660 30064
rect 3620 29850 3648 30058
rect 3608 29844 3660 29850
rect 3608 29786 3660 29792
rect 3712 29714 3740 30194
rect 3148 29708 3200 29714
rect 3148 29650 3200 29656
rect 3240 29708 3292 29714
rect 3700 29708 3752 29714
rect 3240 29650 3292 29656
rect 3620 29668 3700 29696
rect 3056 29504 3108 29510
rect 3056 29446 3108 29452
rect 1306 29336 1362 29345
rect 1306 29271 1362 29280
rect 1320 29238 1348 29271
rect 3068 29238 3096 29446
rect 3620 29238 3648 29668
rect 3700 29650 3752 29656
rect 1308 29232 1360 29238
rect 3056 29232 3108 29238
rect 1308 29174 1360 29180
rect 1950 29200 2006 29209
rect 3056 29174 3108 29180
rect 3608 29232 3660 29238
rect 3608 29174 3660 29180
rect 1950 29135 2006 29144
rect 1306 28656 1362 28665
rect 1306 28591 1308 28600
rect 1360 28591 1362 28600
rect 1308 28562 1360 28568
rect 1400 28008 1452 28014
rect 1398 27976 1400 27985
rect 1452 27976 1454 27985
rect 1398 27911 1454 27920
rect 1412 27402 1440 27911
rect 1400 27396 1452 27402
rect 1400 27338 1452 27344
rect 1676 25696 1728 25702
rect 1676 25638 1728 25644
rect 1688 25226 1716 25638
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 1676 24608 1728 24614
rect 1676 24550 1728 24556
rect 1688 24274 1716 24550
rect 1676 24268 1728 24274
rect 1676 24210 1728 24216
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 23662 1440 24142
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1412 23118 1440 23598
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 21486 1440 23054
rect 1676 23044 1728 23050
rect 1676 22986 1728 22992
rect 1688 22234 1716 22986
rect 1872 22778 1900 23598
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 19854 1440 21422
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 18766 1440 19790
rect 1676 19780 1728 19786
rect 1676 19722 1728 19728
rect 1688 19514 1716 19722
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 17134 1440 18702
rect 1676 18692 1728 18698
rect 1676 18634 1728 18640
rect 1688 18426 1716 18634
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1676 17128 1728 17134
rect 1676 17070 1728 17076
rect 1412 16114 1440 17070
rect 1688 16794 1716 17070
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15570 1440 16050
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1872 15026 1900 15506
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1872 14482 1900 14962
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1872 14074 1900 14418
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1964 13954 1992 29135
rect 2412 28960 2464 28966
rect 2412 28902 2464 28908
rect 2136 27668 2188 27674
rect 2136 27610 2188 27616
rect 2148 26042 2176 27610
rect 2424 27470 2452 28902
rect 3620 28626 3648 29174
rect 3608 28620 3660 28626
rect 3608 28562 3660 28568
rect 2780 28484 2832 28490
rect 2780 28426 2832 28432
rect 2792 28218 2820 28426
rect 2780 28212 2832 28218
rect 2780 28154 2832 28160
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 2504 27872 2556 27878
rect 2504 27814 2556 27820
rect 2412 27464 2464 27470
rect 2412 27406 2464 27412
rect 2136 26036 2188 26042
rect 2136 25978 2188 25984
rect 2148 25378 2176 25978
rect 2320 25832 2372 25838
rect 2320 25774 2372 25780
rect 2148 25350 2268 25378
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2056 14822 2084 23462
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 2148 21146 2176 21422
rect 2136 21140 2188 21146
rect 2136 21082 2188 21088
rect 2240 21010 2268 25350
rect 2332 25158 2360 25774
rect 2320 25152 2372 25158
rect 2320 25094 2372 25100
rect 2228 21004 2280 21010
rect 2228 20946 2280 20952
rect 2136 19508 2188 19514
rect 2136 19450 2188 19456
rect 2148 15366 2176 19450
rect 2240 16726 2268 20946
rect 2332 17678 2360 25094
rect 2516 24886 2544 27814
rect 2792 27062 2820 28154
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 3148 28008 3200 28014
rect 3148 27950 3200 27956
rect 3160 27606 3188 27950
rect 3148 27600 3200 27606
rect 3148 27542 3200 27548
rect 3436 27130 3464 28018
rect 2872 27124 2924 27130
rect 2872 27066 2924 27072
rect 3424 27124 3476 27130
rect 3424 27066 3476 27072
rect 2780 27056 2832 27062
rect 2780 26998 2832 27004
rect 2792 26382 2820 26998
rect 2884 26450 2912 27066
rect 2872 26444 2924 26450
rect 2872 26386 2924 26392
rect 2964 26444 3016 26450
rect 2964 26386 3016 26392
rect 2780 26376 2832 26382
rect 2780 26318 2832 26324
rect 2688 26240 2740 26246
rect 2688 26182 2740 26188
rect 2504 24880 2556 24886
rect 2504 24822 2556 24828
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2424 23186 2452 23598
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 2516 22642 2544 24822
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2516 18222 2544 22578
rect 2700 22250 2728 26182
rect 2792 25294 2820 26318
rect 2884 25702 2912 26386
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 2884 25362 2912 25638
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2780 25288 2832 25294
rect 2780 25230 2832 25236
rect 2792 24206 2820 25230
rect 2884 24818 2912 25298
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2976 24698 3004 26386
rect 3056 26036 3108 26042
rect 3056 25978 3108 25984
rect 3068 24750 3096 25978
rect 3424 25696 3476 25702
rect 3424 25638 3476 25644
rect 3148 25492 3200 25498
rect 3148 25434 3200 25440
rect 3160 25158 3188 25434
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 3148 24880 3200 24886
rect 3146 24848 3148 24857
rect 3200 24848 3202 24857
rect 3146 24783 3202 24792
rect 2884 24670 3004 24698
rect 3056 24744 3108 24750
rect 3056 24686 3108 24692
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2884 23712 2912 24670
rect 3160 24410 3188 24783
rect 3148 24404 3200 24410
rect 3148 24346 3200 24352
rect 2792 23684 2912 23712
rect 2964 23724 3016 23730
rect 2792 23338 2820 23684
rect 2964 23666 3016 23672
rect 2870 23624 2926 23633
rect 2870 23559 2926 23568
rect 2884 23526 2912 23559
rect 2872 23520 2924 23526
rect 2872 23462 2924 23468
rect 2792 23310 2912 23338
rect 2608 22222 2820 22250
rect 2608 19514 2636 22222
rect 2688 22160 2740 22166
rect 2688 22102 2740 22108
rect 2700 21010 2728 22102
rect 2792 22098 2820 22222
rect 2780 22092 2832 22098
rect 2780 22034 2832 22040
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2688 21004 2740 21010
rect 2688 20946 2740 20952
rect 2792 20942 2820 21286
rect 2884 21078 2912 23310
rect 2976 23050 3004 23666
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 2964 23044 3016 23050
rect 2964 22986 3016 22992
rect 2976 22642 3004 22986
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2976 21622 3004 22578
rect 3344 22574 3372 23122
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3344 22098 3372 22510
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3436 21622 3464 25638
rect 2964 21616 3016 21622
rect 2964 21558 3016 21564
rect 3424 21616 3476 21622
rect 3424 21558 3476 21564
rect 2872 21072 2924 21078
rect 2872 21014 2924 21020
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2976 20602 3004 21558
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 3068 20942 3096 21082
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2976 19786 3004 20538
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 3068 19334 3096 20878
rect 3240 20800 3292 20806
rect 3240 20742 3292 20748
rect 2596 19304 2648 19310
rect 3068 19306 3188 19334
rect 2596 19246 2648 19252
rect 2608 18222 2636 19246
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2332 16590 2360 16934
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2424 15910 2452 16594
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 2240 14618 2268 14894
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2424 14074 2452 14282
rect 2516 14278 2544 18158
rect 2608 16658 2636 18158
rect 2792 17202 2820 18702
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 3068 17338 3096 17546
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2608 16153 2636 16594
rect 2594 16144 2650 16153
rect 2792 16114 2820 17138
rect 2594 16079 2650 16088
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 1964 13926 2084 13954
rect 2056 13870 2084 13926
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1688 13530 1716 13806
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 2042 12880 2098 12889
rect 2792 12850 2820 13874
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2884 13394 2912 13738
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13394 3096 13670
rect 2872 13388 2924 13394
rect 3056 13388 3108 13394
rect 2872 13330 2924 13336
rect 2976 13348 3056 13376
rect 2042 12815 2098 12824
rect 2780 12844 2832 12850
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1412 10674 1440 12718
rect 1688 12442 1716 12718
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 2056 12238 2084 12815
rect 2780 12786 2832 12792
rect 2976 12374 3004 13348
rect 3056 13330 3108 13336
rect 3160 12986 3188 19306
rect 3252 17610 3280 20742
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3332 19440 3384 19446
rect 3332 19382 3384 19388
rect 3344 17882 3372 19382
rect 3436 19378 3464 19654
rect 3528 19514 3556 28154
rect 3620 28082 3648 28562
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3700 26920 3752 26926
rect 3700 26862 3752 26868
rect 3712 26586 3740 26862
rect 3700 26580 3752 26586
rect 3700 26522 3752 26528
rect 3608 24404 3660 24410
rect 3608 24346 3660 24352
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 3620 19378 3648 24346
rect 3700 22976 3752 22982
rect 3700 22918 3752 22924
rect 3712 22574 3740 22918
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3712 19854 3740 22510
rect 3700 19848 3752 19854
rect 3804 19825 3832 31726
rect 4172 31414 4200 31962
rect 4356 31754 4384 31980
rect 4436 31962 4488 31968
rect 4344 31748 4396 31754
rect 4344 31690 4396 31696
rect 4252 31680 4304 31686
rect 4252 31622 4304 31628
rect 4264 31482 4292 31622
rect 4252 31476 4304 31482
rect 4252 31418 4304 31424
rect 4632 31414 4660 32302
rect 4724 31890 4752 32370
rect 4712 31884 4764 31890
rect 4712 31826 4764 31832
rect 4160 31408 4212 31414
rect 4160 31350 4212 31356
rect 4620 31408 4672 31414
rect 4620 31350 4672 31356
rect 4724 31346 4752 31826
rect 4712 31340 4764 31346
rect 4712 31282 4764 31288
rect 4068 31272 4120 31278
rect 4068 31214 4120 31220
rect 4620 31272 4672 31278
rect 4620 31214 4672 31220
rect 4080 30938 4108 31214
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30938 4660 31214
rect 4068 30932 4120 30938
rect 4068 30874 4120 30880
rect 4620 30932 4672 30938
rect 4620 30874 4672 30880
rect 3976 30184 4028 30190
rect 3976 30126 4028 30132
rect 3988 29850 4016 30126
rect 3976 29844 4028 29850
rect 3976 29786 4028 29792
rect 4080 29646 4108 30874
rect 4434 30832 4490 30841
rect 4434 30767 4436 30776
rect 4488 30767 4490 30776
rect 4436 30738 4488 30744
rect 4816 30734 4844 32370
rect 4896 32292 4948 32298
rect 4896 32234 4948 32240
rect 4908 31754 4936 32234
rect 5000 32230 5028 32399
rect 5264 32370 5316 32376
rect 5448 32428 5500 32434
rect 5448 32370 5500 32376
rect 5276 32337 5304 32370
rect 5078 32328 5134 32337
rect 5078 32263 5134 32272
rect 5262 32328 5318 32337
rect 5262 32263 5318 32272
rect 5092 32230 5120 32263
rect 5460 32230 5488 32370
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 5080 32224 5132 32230
rect 5080 32166 5132 32172
rect 5448 32224 5500 32230
rect 5448 32166 5500 32172
rect 5092 31890 5120 32166
rect 5080 31884 5132 31890
rect 5080 31826 5132 31832
rect 5460 31822 5488 32166
rect 5644 31890 5672 32846
rect 5828 32774 5856 32846
rect 5816 32768 5868 32774
rect 5816 32710 5868 32716
rect 5828 32586 5856 32710
rect 5736 32558 5856 32586
rect 5736 32366 5764 32558
rect 5724 32360 5776 32366
rect 5724 32302 5776 32308
rect 5632 31884 5684 31890
rect 5632 31826 5684 31832
rect 5448 31816 5500 31822
rect 5736 31793 5764 32302
rect 5816 31816 5868 31822
rect 5448 31758 5500 31764
rect 5722 31784 5778 31793
rect 4908 31748 5304 31754
rect 4908 31726 5080 31748
rect 4908 31686 4936 31726
rect 5132 31726 5304 31748
rect 5080 31690 5132 31696
rect 4896 31680 4948 31686
rect 4896 31622 4948 31628
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 4896 31136 4948 31142
rect 4896 31078 4948 31084
rect 4908 30938 4936 31078
rect 4896 30932 4948 30938
rect 4896 30874 4948 30880
rect 4988 30932 5040 30938
rect 4988 30874 5040 30880
rect 5000 30784 5028 30874
rect 5184 30802 5212 31282
rect 4908 30756 5028 30784
rect 5172 30796 5224 30802
rect 4804 30728 4856 30734
rect 4526 30696 4582 30705
rect 4804 30670 4856 30676
rect 4526 30631 4582 30640
rect 4540 30598 4568 30631
rect 4528 30592 4580 30598
rect 4908 30580 4936 30756
rect 5172 30738 5224 30744
rect 4986 30696 5042 30705
rect 4986 30631 4988 30640
rect 5040 30631 5042 30640
rect 4988 30602 5040 30608
rect 4528 30534 4580 30540
rect 4816 30552 4936 30580
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4068 29640 4120 29646
rect 4068 29582 4120 29588
rect 4080 29102 4108 29582
rect 4712 29504 4764 29510
rect 4712 29446 4764 29452
rect 4068 29096 4120 29102
rect 4068 29038 4120 29044
rect 4080 28490 4108 29038
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28484 4120 28490
rect 4068 28426 4120 28432
rect 4080 27470 4108 28426
rect 4620 27872 4672 27878
rect 4620 27814 4672 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4528 27532 4580 27538
rect 4528 27474 4580 27480
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 4540 26926 4568 27474
rect 4632 27470 4660 27814
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 4528 26920 4580 26926
rect 4528 26862 4580 26868
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 4080 26450 4108 26794
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4436 26512 4488 26518
rect 4436 26454 4488 26460
rect 3884 26444 3936 26450
rect 3884 26386 3936 26392
rect 4068 26444 4120 26450
rect 4068 26386 4120 26392
rect 4344 26444 4396 26450
rect 4344 26386 4396 26392
rect 3896 25770 3924 26386
rect 4356 26042 4384 26386
rect 4448 26042 4476 26454
rect 4632 26382 4660 27066
rect 4620 26376 4672 26382
rect 4724 26364 4752 29446
rect 4816 29238 4844 30552
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5276 30326 5304 31726
rect 5816 31758 5868 31764
rect 5722 31719 5778 31728
rect 5540 31680 5592 31686
rect 5446 31648 5502 31657
rect 5540 31622 5592 31628
rect 5724 31680 5776 31686
rect 5724 31622 5776 31628
rect 5446 31583 5502 31592
rect 5356 30592 5408 30598
rect 5356 30534 5408 30540
rect 5264 30320 5316 30326
rect 5264 30262 5316 30268
rect 5264 30184 5316 30190
rect 5264 30126 5316 30132
rect 5172 30048 5224 30054
rect 5172 29990 5224 29996
rect 5184 29510 5212 29990
rect 5172 29504 5224 29510
rect 5172 29446 5224 29452
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 5276 28966 5304 30126
rect 5368 29889 5396 30534
rect 5354 29880 5410 29889
rect 5354 29815 5410 29824
rect 5368 29578 5396 29815
rect 5356 29572 5408 29578
rect 5356 29514 5408 29520
rect 5460 28994 5488 31583
rect 5552 31414 5580 31622
rect 5736 31482 5764 31622
rect 5724 31476 5776 31482
rect 5724 31418 5776 31424
rect 5540 31408 5592 31414
rect 5540 31350 5592 31356
rect 5540 31272 5592 31278
rect 5828 31260 5856 31758
rect 5920 31362 5948 32846
rect 6012 31498 6040 34138
rect 6092 34128 6144 34134
rect 6092 34070 6144 34076
rect 6104 33504 6132 34070
rect 6196 33658 6224 34546
rect 6380 34202 6408 35022
rect 6368 34196 6420 34202
rect 6368 34138 6420 34144
rect 6276 33992 6328 33998
rect 6276 33934 6328 33940
rect 6184 33652 6236 33658
rect 6184 33594 6236 33600
rect 6184 33516 6236 33522
rect 6104 33476 6184 33504
rect 6184 33458 6236 33464
rect 6184 33312 6236 33318
rect 6184 33254 6236 33260
rect 6196 33114 6224 33254
rect 6184 33108 6236 33114
rect 6184 33050 6236 33056
rect 6092 32904 6144 32910
rect 6092 32846 6144 32852
rect 6184 32904 6236 32910
rect 6288 32881 6316 33934
rect 6472 33538 6500 35022
rect 7012 34944 7064 34950
rect 7012 34886 7064 34892
rect 7024 34610 7052 34886
rect 7116 34678 7144 35022
rect 7104 34672 7156 34678
rect 7104 34614 7156 34620
rect 7300 34610 7328 35022
rect 7392 34610 7420 35158
rect 7668 35086 7696 35498
rect 7852 35290 7880 36110
rect 8312 35834 8340 36178
rect 8300 35828 8352 35834
rect 8300 35770 8352 35776
rect 7932 35760 7984 35766
rect 7932 35702 7984 35708
rect 7840 35284 7892 35290
rect 7840 35226 7892 35232
rect 7944 35086 7972 35702
rect 8208 35284 8260 35290
rect 8208 35226 8260 35232
rect 7656 35080 7708 35086
rect 7656 35022 7708 35028
rect 7932 35080 7984 35086
rect 7932 35022 7984 35028
rect 7668 34610 7696 35022
rect 7012 34604 7064 34610
rect 7012 34546 7064 34552
rect 7288 34604 7340 34610
rect 7288 34546 7340 34552
rect 7380 34604 7432 34610
rect 7380 34546 7432 34552
rect 7472 34604 7524 34610
rect 7472 34546 7524 34552
rect 7656 34604 7708 34610
rect 7656 34546 7708 34552
rect 7104 34536 7156 34542
rect 7104 34478 7156 34484
rect 7116 34134 7144 34478
rect 7196 34400 7248 34406
rect 7196 34342 7248 34348
rect 7012 34128 7064 34134
rect 7012 34070 7064 34076
rect 7104 34128 7156 34134
rect 7104 34070 7156 34076
rect 6828 33992 6880 33998
rect 6828 33934 6880 33940
rect 6920 33992 6972 33998
rect 6920 33934 6972 33940
rect 6552 33856 6604 33862
rect 6550 33824 6552 33833
rect 6644 33856 6696 33862
rect 6604 33824 6606 33833
rect 6644 33798 6696 33804
rect 6550 33759 6606 33768
rect 6656 33590 6684 33798
rect 6380 33510 6500 33538
rect 6644 33584 6696 33590
rect 6644 33526 6696 33532
rect 6736 33516 6788 33522
rect 6184 32846 6236 32852
rect 6274 32872 6330 32881
rect 6104 32774 6132 32846
rect 6092 32768 6144 32774
rect 6092 32710 6144 32716
rect 6104 32570 6132 32710
rect 6092 32564 6144 32570
rect 6092 32506 6144 32512
rect 6196 32366 6224 32846
rect 6274 32807 6330 32816
rect 6184 32360 6236 32366
rect 6182 32328 6184 32337
rect 6236 32328 6238 32337
rect 6092 32292 6144 32298
rect 6182 32263 6238 32272
rect 6092 32234 6144 32240
rect 6104 31822 6132 32234
rect 6092 31816 6144 31822
rect 6092 31758 6144 31764
rect 6104 31686 6132 31758
rect 6092 31680 6144 31686
rect 6288 31657 6316 32807
rect 6092 31622 6144 31628
rect 6274 31648 6330 31657
rect 6274 31583 6330 31592
rect 6012 31470 6316 31498
rect 5920 31334 6224 31362
rect 6288 31346 6316 31470
rect 5540 31214 5592 31220
rect 5722 31240 5778 31249
rect 5552 30734 5580 31214
rect 5828 31232 5948 31260
rect 5722 31175 5724 31184
rect 5776 31175 5778 31184
rect 5724 31146 5776 31152
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5816 31136 5868 31142
rect 5816 31078 5868 31084
rect 5540 30728 5592 30734
rect 5540 30670 5592 30676
rect 5540 30592 5592 30598
rect 5540 30534 5592 30540
rect 5552 29646 5580 30534
rect 5644 29646 5672 31078
rect 5722 30968 5778 30977
rect 5722 30903 5724 30912
rect 5776 30903 5778 30912
rect 5724 30874 5776 30880
rect 5724 30660 5776 30666
rect 5724 30602 5776 30608
rect 5736 30394 5764 30602
rect 5724 30388 5776 30394
rect 5724 30330 5776 30336
rect 5724 30252 5776 30258
rect 5724 30194 5776 30200
rect 5540 29640 5592 29646
rect 5540 29582 5592 29588
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5736 29510 5764 30194
rect 5828 30190 5856 31078
rect 5920 30938 5948 31232
rect 6092 31136 6144 31142
rect 6092 31078 6144 31084
rect 5908 30932 5960 30938
rect 5908 30874 5960 30880
rect 6104 30666 6132 31078
rect 6092 30660 6144 30666
rect 6092 30602 6144 30608
rect 6000 30592 6052 30598
rect 6000 30534 6052 30540
rect 6012 30394 6040 30534
rect 6000 30388 6052 30394
rect 6000 30330 6052 30336
rect 5816 30184 5868 30190
rect 5816 30126 5868 30132
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5724 29504 5776 29510
rect 5724 29446 5776 29452
rect 5736 29209 5764 29446
rect 5722 29200 5778 29209
rect 5722 29135 5778 29144
rect 5460 28966 5672 28994
rect 5264 28960 5316 28966
rect 5264 28902 5316 28908
rect 5356 28960 5408 28966
rect 5356 28902 5408 28908
rect 5368 28626 5396 28902
rect 5356 28620 5408 28626
rect 5356 28562 5408 28568
rect 5262 28520 5318 28529
rect 5262 28455 5264 28464
rect 5316 28455 5318 28464
rect 5264 28426 5316 28432
rect 4804 28416 4856 28422
rect 4804 28358 4856 28364
rect 4816 27402 4844 28358
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5276 28082 5304 28426
rect 5264 28076 5316 28082
rect 5264 28018 5316 28024
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 5000 27674 5028 27950
rect 5264 27940 5316 27946
rect 5264 27882 5316 27888
rect 5276 27674 5304 27882
rect 4988 27668 5040 27674
rect 4988 27610 5040 27616
rect 5264 27668 5316 27674
rect 5264 27610 5316 27616
rect 5368 27538 5396 28562
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 4804 27396 4856 27402
rect 4804 27338 4856 27344
rect 4816 26518 4844 27338
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5368 27062 5396 27270
rect 5356 27056 5408 27062
rect 5356 26998 5408 27004
rect 4988 26920 5040 26926
rect 4988 26862 5040 26868
rect 4804 26512 4856 26518
rect 4804 26454 4856 26460
rect 5000 26382 5028 26862
rect 5264 26852 5316 26858
rect 5264 26794 5316 26800
rect 4988 26376 5040 26382
rect 4724 26336 4844 26364
rect 4620 26318 4672 26324
rect 4712 26240 4764 26246
rect 4712 26182 4764 26188
rect 4724 26042 4752 26182
rect 4344 26036 4396 26042
rect 4344 25978 4396 25984
rect 4436 26036 4488 26042
rect 4436 25978 4488 25984
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4356 25906 4384 25978
rect 4620 25968 4672 25974
rect 4620 25910 4672 25916
rect 3976 25900 4028 25906
rect 3976 25842 4028 25848
rect 4344 25900 4396 25906
rect 4344 25842 4396 25848
rect 3884 25764 3936 25770
rect 3884 25706 3936 25712
rect 3988 25294 4016 25842
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25498 4660 25910
rect 4712 25832 4764 25838
rect 4712 25774 4764 25780
rect 4724 25498 4752 25774
rect 4620 25492 4672 25498
rect 4620 25434 4672 25440
rect 4712 25492 4764 25498
rect 4712 25434 4764 25440
rect 3976 25288 4028 25294
rect 3976 25230 4028 25236
rect 3988 24954 4016 25230
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 3976 24948 4028 24954
rect 3976 24890 4028 24896
rect 3976 24744 4028 24750
rect 3976 24686 4028 24692
rect 3988 24410 4016 24686
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 4080 24177 4108 25162
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4066 24168 4122 24177
rect 4066 24103 4122 24112
rect 4080 23798 4108 24103
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4252 23316 4304 23322
rect 4632 23304 4660 25094
rect 4816 24274 4844 26336
rect 4988 26318 5040 26324
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5276 26042 5304 26794
rect 5368 26586 5396 26998
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5264 26036 5316 26042
rect 5264 25978 5316 25984
rect 5368 25922 5396 26182
rect 5000 25894 5396 25922
rect 5000 25838 5028 25894
rect 4988 25832 5040 25838
rect 4988 25774 5040 25780
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 5356 25696 5408 25702
rect 5356 25638 5408 25644
rect 5276 25362 5304 25638
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5276 24274 5304 24550
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 5264 24268 5316 24274
rect 5264 24210 5316 24216
rect 4816 23730 4844 24210
rect 5368 24138 5396 25638
rect 5460 25158 5488 26726
rect 5540 25832 5592 25838
rect 5540 25774 5592 25780
rect 5552 25362 5580 25774
rect 5540 25356 5592 25362
rect 5540 25298 5592 25304
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 5552 24970 5580 25298
rect 5460 24942 5580 24970
rect 5460 24313 5488 24942
rect 5446 24304 5502 24313
rect 5446 24239 5448 24248
rect 5500 24239 5502 24248
rect 5448 24210 5500 24216
rect 5356 24132 5408 24138
rect 5356 24074 5408 24080
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5356 23792 5408 23798
rect 5354 23760 5356 23769
rect 5408 23760 5410 23769
rect 4804 23724 4856 23730
rect 5354 23695 5410 23704
rect 4804 23666 4856 23672
rect 5356 23588 5408 23594
rect 5356 23530 5408 23536
rect 4712 23520 4764 23526
rect 5264 23520 5316 23526
rect 4712 23462 4764 23468
rect 5078 23488 5134 23497
rect 4252 23258 4304 23264
rect 4356 23276 4660 23304
rect 3884 23248 3936 23254
rect 3884 23190 3936 23196
rect 3700 19790 3752 19796
rect 3790 19816 3846 19825
rect 3790 19751 3846 19760
rect 3896 19700 3924 23190
rect 4264 23186 4292 23258
rect 4252 23180 4304 23186
rect 4252 23122 4304 23128
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3804 19672 3924 19700
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3528 18290 3556 18906
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3804 17678 3832 19672
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3896 18970 3924 19314
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 3882 18864 3938 18873
rect 3882 18799 3938 18808
rect 3424 17672 3476 17678
rect 3792 17672 3844 17678
rect 3424 17614 3476 17620
rect 3698 17640 3754 17649
rect 3240 17604 3292 17610
rect 3240 17546 3292 17552
rect 3332 16584 3384 16590
rect 3330 16552 3332 16561
rect 3384 16552 3386 16561
rect 3330 16487 3386 16496
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3252 15094 3280 15438
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3252 14414 3280 15030
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 13938 3280 14350
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3252 12986 3280 13194
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 8498 1440 10610
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10062 1716 10406
rect 1676 10056 1728 10062
rect 2240 10033 2268 12174
rect 2424 11898 2452 12242
rect 3068 12238 3096 12650
rect 3160 12374 3188 12922
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 1676 9998 1728 10004
rect 2226 10024 2282 10033
rect 2226 9959 2282 9968
rect 2332 9654 2360 10406
rect 2424 10062 2452 11222
rect 2516 11082 2544 11698
rect 2792 11234 2820 11698
rect 2884 11354 2912 12106
rect 3068 11626 3096 12174
rect 3160 11898 3188 12174
rect 3344 11898 3372 12174
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 3344 11286 3372 11834
rect 3332 11280 3384 11286
rect 2792 11206 2912 11234
rect 3332 11222 3384 11228
rect 2884 11150 2912 11206
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 3148 11144 3200 11150
rect 3200 11104 3372 11132
rect 3148 11086 3200 11092
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2424 9926 2452 9998
rect 2516 9994 2544 11018
rect 2608 10266 2636 11086
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2424 9586 2452 9862
rect 2700 9654 2728 11086
rect 2884 10198 2912 11086
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2516 8498 2544 9046
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2976 7478 3004 10678
rect 3068 9518 3096 10950
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3160 9994 3188 10746
rect 3344 10713 3372 11104
rect 3436 10810 3464 17614
rect 3608 17604 3660 17610
rect 3792 17614 3844 17620
rect 3698 17575 3754 17584
rect 3608 17546 3660 17552
rect 3620 17270 3648 17546
rect 3608 17264 3660 17270
rect 3608 17206 3660 17212
rect 3712 16794 3740 17575
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3620 16250 3648 16390
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3712 14890 3740 16458
rect 3896 16250 3924 18799
rect 3988 17202 4016 23054
rect 4068 22976 4120 22982
rect 4252 22976 4304 22982
rect 4068 22918 4120 22924
rect 4250 22944 4252 22953
rect 4356 22964 4384 23276
rect 4528 23112 4580 23118
rect 4304 22944 4384 22964
rect 4306 22936 4384 22944
rect 4448 23072 4528 23100
rect 4080 22710 4108 22918
rect 4250 22879 4306 22888
rect 4448 22817 4476 23072
rect 4528 23054 4580 23060
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4434 22808 4490 22817
rect 4434 22743 4490 22752
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 4160 22704 4212 22710
rect 4160 22646 4212 22652
rect 4172 22556 4200 22646
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 4080 22528 4200 22556
rect 4080 22438 4108 22528
rect 4356 22506 4384 22578
rect 4344 22500 4396 22506
rect 4344 22442 4396 22448
rect 4068 22432 4120 22438
rect 4068 22374 4120 22380
rect 4080 22098 4108 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22234 4660 22986
rect 4724 22778 4752 23462
rect 5264 23462 5316 23468
rect 5078 23423 5134 23432
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4080 21554 4108 22034
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 20942 4660 21966
rect 4724 21962 4752 22374
rect 4816 21962 4844 22986
rect 5092 22982 5120 23423
rect 5170 23352 5226 23361
rect 5170 23287 5226 23296
rect 5184 23118 5212 23287
rect 5276 23225 5304 23462
rect 5262 23216 5318 23225
rect 5262 23151 5318 23160
rect 5172 23112 5224 23118
rect 5172 23054 5224 23060
rect 5080 22976 5132 22982
rect 5080 22918 5132 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4896 22772 4948 22778
rect 4896 22714 4948 22720
rect 4908 22681 4936 22714
rect 4894 22672 4950 22681
rect 5276 22642 5304 23151
rect 5368 22794 5396 23530
rect 5368 22766 5488 22794
rect 4894 22607 4950 22616
rect 5264 22636 5316 22642
rect 5264 22578 5316 22584
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5170 22536 5226 22545
rect 5092 22166 5120 22510
rect 5170 22471 5226 22480
rect 5080 22160 5132 22166
rect 5080 22102 5132 22108
rect 5184 22098 5212 22471
rect 5276 22438 5304 22578
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5276 22030 5304 22374
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 4712 21956 4764 21962
rect 4712 21898 4764 21904
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4724 21010 4752 21490
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4620 20936 4672 20942
rect 4618 20904 4620 20913
rect 4672 20904 4674 20913
rect 4618 20839 4674 20848
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4540 20466 4568 20742
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4436 19916 4488 19922
rect 4436 19858 4488 19864
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3884 16244 3936 16250
rect 3804 16204 3884 16232
rect 3700 14884 3752 14890
rect 3700 14826 3752 14832
rect 3712 14414 3740 14826
rect 3804 14482 3832 16204
rect 3884 16186 3936 16192
rect 3882 16144 3938 16153
rect 3882 16079 3938 16088
rect 3896 16046 3924 16079
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3712 14074 3740 14214
rect 3700 14068 3752 14074
rect 3752 14028 3924 14056
rect 3700 14010 3752 14016
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3620 12442 3648 12786
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3712 12306 3740 12718
rect 3804 12306 3832 13126
rect 3896 12753 3924 14028
rect 3988 13802 4016 17138
rect 4080 17066 4108 19450
rect 4264 19378 4292 19790
rect 4344 19780 4396 19786
rect 4344 19722 4396 19728
rect 4356 19514 4384 19722
rect 4448 19514 4476 19858
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4632 19292 4660 20334
rect 4724 19446 4752 20946
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4632 19264 4752 19292
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18902 4660 19110
rect 4620 18896 4672 18902
rect 4620 18838 4672 18844
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4448 18193 4476 18702
rect 4434 18184 4490 18193
rect 4434 18119 4490 18128
rect 4618 18048 4674 18057
rect 4214 17980 4522 17989
rect 4618 17983 4674 17992
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 17983
rect 4724 17921 4752 19264
rect 4816 18034 4844 21286
rect 5000 20942 5028 21626
rect 5276 21486 5304 21830
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 5276 21010 5304 21422
rect 5368 21010 5396 21490
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5356 21004 5408 21010
rect 5356 20946 5408 20952
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5078 20496 5134 20505
rect 4896 20460 4948 20466
rect 5078 20431 5134 20440
rect 4896 20402 4948 20408
rect 4908 20058 4936 20402
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 5092 19922 5120 20431
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4908 18766 4936 19450
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 5000 18834 5028 19314
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4816 18006 4936 18034
rect 4710 17912 4766 17921
rect 4620 17876 4672 17882
rect 4710 17847 4766 17856
rect 4620 17818 4672 17824
rect 4908 17796 4936 18006
rect 4342 17776 4398 17785
rect 4342 17711 4344 17720
rect 4396 17711 4398 17720
rect 4816 17768 4936 17796
rect 4344 17682 4396 17688
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 4172 16998 4200 17546
rect 4250 17368 4306 17377
rect 4250 17303 4252 17312
rect 4304 17303 4306 17312
rect 4252 17274 4304 17280
rect 4356 17202 4384 17682
rect 4816 17678 4844 17768
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4804 17672 4856 17678
rect 4896 17672 4948 17678
rect 4804 17614 4856 17620
rect 4894 17640 4896 17649
rect 4948 17640 4950 17649
rect 4540 17202 4568 17614
rect 4724 17377 4752 17614
rect 4894 17575 4950 17584
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4710 17368 4766 17377
rect 4710 17303 4766 17312
rect 4816 17270 4844 17478
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 5276 17134 5304 20742
rect 5460 20380 5488 22766
rect 5552 22545 5580 24074
rect 5644 23662 5672 28966
rect 5828 28762 5856 29582
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5724 28552 5776 28558
rect 5724 28494 5776 28500
rect 5736 28218 5764 28494
rect 5724 28212 5776 28218
rect 5724 28154 5776 28160
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 5736 26994 5764 27270
rect 5724 26988 5776 26994
rect 5724 26930 5776 26936
rect 5724 26444 5776 26450
rect 5724 26386 5776 26392
rect 5736 25265 5764 26386
rect 5722 25256 5778 25265
rect 5722 25191 5778 25200
rect 5724 25152 5776 25158
rect 5724 25094 5776 25100
rect 5736 24886 5764 25094
rect 5724 24880 5776 24886
rect 5724 24822 5776 24828
rect 5828 24410 5856 28698
rect 6000 28144 6052 28150
rect 6000 28086 6052 28092
rect 5908 28076 5960 28082
rect 5908 28018 5960 28024
rect 5920 27334 5948 28018
rect 6012 27470 6040 28086
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 6092 27396 6144 27402
rect 6092 27338 6144 27344
rect 5908 27328 5960 27334
rect 5906 27296 5908 27305
rect 5960 27296 5962 27305
rect 5906 27231 5962 27240
rect 6000 26580 6052 26586
rect 6000 26522 6052 26528
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5920 24954 5948 25230
rect 6012 25208 6040 26522
rect 6104 26314 6132 27338
rect 6092 26308 6144 26314
rect 6092 26250 6144 26256
rect 6104 26042 6132 26250
rect 6092 26036 6144 26042
rect 6092 25978 6144 25984
rect 6092 25220 6144 25226
rect 6012 25180 6092 25208
rect 6092 25162 6144 25168
rect 6104 25129 6132 25162
rect 6090 25120 6146 25129
rect 6090 25055 6146 25064
rect 6090 24984 6146 24993
rect 5908 24948 5960 24954
rect 6090 24919 6146 24928
rect 5908 24890 5960 24896
rect 6104 24886 6132 24919
rect 6092 24880 6144 24886
rect 6092 24822 6144 24828
rect 6196 24426 6224 31334
rect 6276 31340 6328 31346
rect 6276 31282 6328 31288
rect 6288 30394 6316 31282
rect 6276 30388 6328 30394
rect 6276 30330 6328 30336
rect 6288 29714 6316 30330
rect 6276 29708 6328 29714
rect 6276 29650 6328 29656
rect 6274 28792 6330 28801
rect 6274 28727 6330 28736
rect 6288 28694 6316 28727
rect 6276 28688 6328 28694
rect 6276 28630 6328 28636
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 5816 24404 5868 24410
rect 5816 24346 5868 24352
rect 6104 24398 6224 24426
rect 5816 24132 5868 24138
rect 5816 24074 5868 24080
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 5828 23730 5856 24074
rect 5816 23724 5868 23730
rect 5816 23666 5868 23672
rect 5632 23656 5684 23662
rect 5632 23598 5684 23604
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5644 23120 5672 23462
rect 5632 23114 5684 23120
rect 5632 23056 5684 23062
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5644 22681 5672 22918
rect 5630 22672 5686 22681
rect 5630 22607 5686 22616
rect 5538 22536 5594 22545
rect 5538 22471 5594 22480
rect 5736 22234 5764 23598
rect 5828 22817 5856 23666
rect 5906 23624 5962 23633
rect 5906 23559 5962 23568
rect 5920 23526 5948 23559
rect 5908 23520 5960 23526
rect 5908 23462 5960 23468
rect 6012 23322 6040 24074
rect 6104 23866 6132 24398
rect 6184 24336 6236 24342
rect 6288 24324 6316 26318
rect 6236 24296 6316 24324
rect 6184 24278 6236 24284
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 6090 23624 6146 23633
rect 6090 23559 6146 23568
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 6000 23316 6052 23322
rect 6000 23258 6052 23264
rect 5814 22808 5870 22817
rect 5814 22743 5870 22752
rect 5814 22672 5870 22681
rect 5814 22607 5816 22616
rect 5868 22607 5870 22616
rect 5816 22578 5868 22584
rect 5816 22500 5868 22506
rect 5816 22442 5868 22448
rect 5724 22228 5776 22234
rect 5724 22170 5776 22176
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5552 21486 5580 22102
rect 5828 21690 5856 22442
rect 5920 22098 5948 23258
rect 6000 23044 6052 23050
rect 6104 23032 6132 23559
rect 6052 23004 6132 23032
rect 6000 22986 6052 22992
rect 6090 22808 6146 22817
rect 6090 22743 6146 22752
rect 5998 22672 6054 22681
rect 6104 22642 6132 22743
rect 5998 22607 6000 22616
rect 6052 22607 6054 22616
rect 6092 22636 6144 22642
rect 6000 22578 6052 22584
rect 6092 22578 6144 22584
rect 6092 22432 6144 22438
rect 6092 22374 6144 22380
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5630 20904 5686 20913
rect 5630 20839 5686 20848
rect 5644 20398 5672 20839
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5368 20352 5488 20380
rect 5632 20392 5684 20398
rect 5368 18698 5396 20352
rect 5632 20334 5684 20340
rect 5538 19952 5594 19961
rect 5538 19887 5594 19896
rect 5552 19718 5580 19887
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5460 18970 5488 19314
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5356 18692 5408 18698
rect 5356 18634 5408 18640
rect 5460 18426 5488 18770
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5460 17785 5488 18362
rect 5446 17776 5502 17785
rect 5446 17711 5502 17720
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5368 17270 5396 17614
rect 5552 17610 5580 19654
rect 5828 19446 5856 20402
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5736 18222 5764 19246
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 5644 17338 5672 17546
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5552 17218 5580 17274
rect 4804 17128 4856 17134
rect 5264 17128 5316 17134
rect 4856 17076 4936 17082
rect 4804 17070 4936 17076
rect 5264 17070 5316 17076
rect 4816 17054 4936 17070
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4356 16182 4384 16594
rect 4448 16590 4476 16730
rect 4526 16688 4582 16697
rect 4526 16623 4582 16632
rect 4436 16584 4488 16590
rect 4434 16552 4436 16561
rect 4488 16552 4490 16561
rect 4540 16522 4568 16623
rect 4816 16538 4844 16934
rect 4908 16658 4936 17054
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4434 16487 4490 16496
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4724 16510 4844 16538
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 15094 4108 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15201 4660 16458
rect 4618 15192 4674 15201
rect 4618 15127 4674 15136
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4264 13938 4292 14418
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4448 13870 4476 14418
rect 4436 13864 4488 13870
rect 4632 13841 4660 15127
rect 4724 14550 4752 16510
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 15706 4844 16390
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5368 16114 5396 17206
rect 5552 17190 5672 17218
rect 5736 17202 5764 18158
rect 5828 17882 5856 19382
rect 6104 18204 6132 22374
rect 6196 19854 6224 24278
rect 6380 24206 6408 33510
rect 6736 33458 6788 33464
rect 6460 33448 6512 33454
rect 6460 33390 6512 33396
rect 6472 33114 6500 33390
rect 6460 33108 6512 33114
rect 6460 33050 6512 33056
rect 6552 33108 6604 33114
rect 6552 33050 6604 33056
rect 6644 33108 6696 33114
rect 6644 33050 6696 33056
rect 6458 33008 6514 33017
rect 6564 32978 6592 33050
rect 6656 32978 6684 33050
rect 6748 32978 6776 33458
rect 6458 32943 6514 32952
rect 6552 32972 6604 32978
rect 6472 32502 6500 32943
rect 6552 32914 6604 32920
rect 6644 32972 6696 32978
rect 6644 32914 6696 32920
rect 6736 32972 6788 32978
rect 6736 32914 6788 32920
rect 6840 32858 6868 33934
rect 6932 33318 6960 33934
rect 6920 33312 6972 33318
rect 6920 33254 6972 33260
rect 6656 32842 6868 32858
rect 6644 32836 6868 32842
rect 6696 32830 6868 32836
rect 6644 32778 6696 32784
rect 6736 32768 6788 32774
rect 6736 32710 6788 32716
rect 6828 32768 6880 32774
rect 6828 32710 6880 32716
rect 6748 32570 6776 32710
rect 6736 32564 6788 32570
rect 6736 32506 6788 32512
rect 6460 32496 6512 32502
rect 6840 32473 6868 32710
rect 6932 32570 6960 33254
rect 6920 32564 6972 32570
rect 6920 32506 6972 32512
rect 6460 32438 6512 32444
rect 6826 32464 6882 32473
rect 6826 32399 6882 32408
rect 6552 32360 6604 32366
rect 6552 32302 6604 32308
rect 6564 31958 6592 32302
rect 7024 32026 7052 34070
rect 7208 33998 7236 34342
rect 7196 33992 7248 33998
rect 7196 33934 7248 33940
rect 7288 33992 7340 33998
rect 7288 33934 7340 33940
rect 7104 33856 7156 33862
rect 7104 33798 7156 33804
rect 7116 32910 7144 33798
rect 7208 33658 7236 33934
rect 7196 33652 7248 33658
rect 7196 33594 7248 33600
rect 7300 33640 7328 33934
rect 7392 33862 7420 34546
rect 7484 34066 7512 34546
rect 7472 34060 7524 34066
rect 7472 34002 7524 34008
rect 7380 33856 7432 33862
rect 7380 33798 7432 33804
rect 7300 33612 7512 33640
rect 7196 33516 7248 33522
rect 7300 33504 7328 33612
rect 7248 33476 7328 33504
rect 7380 33516 7432 33522
rect 7196 33458 7248 33464
rect 7380 33458 7432 33464
rect 7288 33380 7340 33386
rect 7288 33322 7340 33328
rect 7196 33312 7248 33318
rect 7196 33254 7248 33260
rect 7208 33114 7236 33254
rect 7300 33114 7328 33322
rect 7196 33108 7248 33114
rect 7196 33050 7248 33056
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 7392 33046 7420 33458
rect 7380 33040 7432 33046
rect 7378 33008 7380 33017
rect 7432 33008 7434 33017
rect 7378 32943 7434 32952
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7484 32434 7512 33612
rect 7104 32428 7156 32434
rect 7472 32428 7524 32434
rect 7156 32388 7472 32416
rect 7104 32370 7156 32376
rect 7012 32020 7064 32026
rect 7012 31962 7064 31968
rect 6552 31952 6604 31958
rect 6552 31894 6604 31900
rect 6920 31952 6972 31958
rect 6920 31894 6972 31900
rect 6460 31680 6512 31686
rect 6460 31622 6512 31628
rect 6472 30666 6500 31622
rect 6564 31346 6592 31894
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6642 31648 6698 31657
rect 6642 31583 6698 31592
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 6460 30660 6512 30666
rect 6460 30602 6512 30608
rect 6472 30433 6500 30602
rect 6552 30592 6604 30598
rect 6552 30534 6604 30540
rect 6458 30424 6514 30433
rect 6458 30359 6514 30368
rect 6564 29646 6592 30534
rect 6552 29640 6604 29646
rect 6552 29582 6604 29588
rect 6460 29232 6512 29238
rect 6460 29174 6512 29180
rect 6472 28558 6500 29174
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 6472 27554 6500 28494
rect 6472 27526 6592 27554
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6472 27062 6500 27406
rect 6460 27056 6512 27062
rect 6460 26998 6512 27004
rect 6460 26580 6512 26586
rect 6460 26522 6512 26528
rect 6472 24614 6500 26522
rect 6564 26314 6592 27526
rect 6552 26308 6604 26314
rect 6552 26250 6604 26256
rect 6564 25906 6592 26250
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6460 24608 6512 24614
rect 6460 24550 6512 24556
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 6276 24132 6328 24138
rect 6276 24074 6328 24080
rect 6288 23526 6316 24074
rect 6380 23712 6408 24142
rect 6472 23848 6500 24550
rect 6656 24154 6684 31583
rect 6840 31482 6868 31758
rect 6932 31482 6960 31894
rect 6828 31476 6880 31482
rect 6828 31418 6880 31424
rect 6920 31476 6972 31482
rect 6920 31418 6972 31424
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 6736 30728 6788 30734
rect 6736 30670 6788 30676
rect 6748 30258 6776 30670
rect 6736 30252 6788 30258
rect 6736 30194 6788 30200
rect 6736 28416 6788 28422
rect 6736 28358 6788 28364
rect 6748 28082 6776 28358
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 6736 25832 6788 25838
rect 6736 25774 6788 25780
rect 6748 24818 6776 25774
rect 6840 25226 6868 31282
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 6932 30734 6960 31214
rect 7208 30734 7236 32388
rect 7472 32370 7524 32376
rect 7564 32428 7616 32434
rect 7564 32370 7616 32376
rect 7300 32298 7512 32314
rect 7300 32292 7524 32298
rect 7300 32286 7472 32292
rect 7300 30870 7328 32286
rect 7472 32234 7524 32240
rect 7380 32224 7432 32230
rect 7380 32166 7432 32172
rect 7392 31346 7420 32166
rect 7576 32026 7604 32370
rect 7668 32348 7696 34546
rect 7840 34536 7892 34542
rect 7840 34478 7892 34484
rect 7852 34202 7880 34478
rect 7944 34474 7972 35022
rect 8220 34610 8248 35226
rect 8208 34604 8260 34610
rect 8208 34546 8260 34552
rect 7932 34468 7984 34474
rect 7932 34410 7984 34416
rect 7840 34196 7892 34202
rect 7840 34138 7892 34144
rect 7748 33992 7800 33998
rect 7748 33934 7800 33940
rect 7760 32842 7788 33934
rect 7944 32910 7972 34410
rect 8208 34060 8260 34066
rect 8208 34002 8260 34008
rect 8116 33992 8168 33998
rect 8116 33934 8168 33940
rect 8128 33658 8156 33934
rect 8116 33652 8168 33658
rect 8116 33594 8168 33600
rect 8116 33448 8168 33454
rect 8116 33390 8168 33396
rect 8128 33114 8156 33390
rect 8116 33108 8168 33114
rect 8116 33050 8168 33056
rect 7932 32904 7984 32910
rect 7932 32846 7984 32852
rect 8024 32904 8076 32910
rect 8076 32864 8156 32892
rect 8024 32846 8076 32852
rect 7748 32836 7800 32842
rect 7748 32778 7800 32784
rect 7668 32320 7788 32348
rect 7656 32224 7708 32230
rect 7656 32166 7708 32172
rect 7564 32020 7616 32026
rect 7564 31962 7616 31968
rect 7472 31884 7524 31890
rect 7472 31826 7524 31832
rect 7484 31414 7512 31826
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7472 31408 7524 31414
rect 7472 31350 7524 31356
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7484 31210 7512 31350
rect 7576 31278 7604 31758
rect 7668 31754 7696 32166
rect 7656 31748 7708 31754
rect 7656 31690 7708 31696
rect 7668 31482 7696 31690
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7564 31272 7616 31278
rect 7564 31214 7616 31220
rect 7472 31204 7524 31210
rect 7472 31146 7524 31152
rect 7576 30938 7604 31214
rect 7564 30932 7616 30938
rect 7564 30874 7616 30880
rect 7760 30870 7788 32320
rect 7944 32298 7972 32846
rect 7932 32292 7984 32298
rect 7932 32234 7984 32240
rect 8022 32056 8078 32065
rect 8022 31991 8024 32000
rect 8076 31991 8078 32000
rect 8024 31962 8076 31968
rect 8128 31958 8156 32864
rect 8116 31952 8168 31958
rect 8116 31894 8168 31900
rect 7840 31816 7892 31822
rect 7840 31758 7892 31764
rect 7852 31346 7880 31758
rect 7932 31476 7984 31482
rect 7932 31418 7984 31424
rect 7840 31340 7892 31346
rect 7840 31282 7892 31288
rect 7852 30938 7880 31282
rect 7840 30932 7892 30938
rect 7840 30874 7892 30880
rect 7288 30864 7340 30870
rect 7748 30864 7800 30870
rect 7288 30806 7340 30812
rect 7576 30812 7748 30818
rect 7944 30818 7972 31418
rect 7576 30806 7800 30812
rect 7576 30790 7788 30806
rect 7852 30790 7972 30818
rect 7576 30734 7604 30790
rect 6920 30728 6972 30734
rect 6920 30670 6972 30676
rect 7104 30728 7156 30734
rect 7104 30670 7156 30676
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 7564 30728 7616 30734
rect 7564 30670 7616 30676
rect 6932 30122 6960 30670
rect 7012 30184 7064 30190
rect 7012 30126 7064 30132
rect 6920 30116 6972 30122
rect 6920 30058 6972 30064
rect 7024 29034 7052 30126
rect 7116 30054 7144 30670
rect 7288 30252 7340 30258
rect 7288 30194 7340 30200
rect 7104 30048 7156 30054
rect 7104 29990 7156 29996
rect 7300 29753 7328 30194
rect 7656 30184 7708 30190
rect 7656 30126 7708 30132
rect 7286 29744 7342 29753
rect 7104 29708 7156 29714
rect 7286 29679 7342 29688
rect 7104 29650 7156 29656
rect 7116 29238 7144 29650
rect 7104 29232 7156 29238
rect 7104 29174 7156 29180
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7012 29028 7064 29034
rect 7012 28970 7064 28976
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 6932 28150 6960 28698
rect 7024 28558 7052 28970
rect 7104 28688 7156 28694
rect 7104 28630 7156 28636
rect 7012 28552 7064 28558
rect 7012 28494 7064 28500
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 7012 28144 7064 28150
rect 7012 28086 7064 28092
rect 6920 25356 6972 25362
rect 6920 25298 6972 25304
rect 6932 25226 6960 25298
rect 6828 25220 6880 25226
rect 6828 25162 6880 25168
rect 6920 25220 6972 25226
rect 6920 25162 6972 25168
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6564 24138 6684 24154
rect 6552 24132 6684 24138
rect 6604 24126 6684 24132
rect 6552 24074 6604 24080
rect 6472 23820 6684 23848
rect 6550 23760 6606 23769
rect 6460 23724 6512 23730
rect 6380 23684 6460 23712
rect 6550 23695 6606 23704
rect 6460 23666 6512 23672
rect 6460 23588 6512 23594
rect 6460 23530 6512 23536
rect 6276 23520 6328 23526
rect 6276 23462 6328 23468
rect 6368 23316 6420 23322
rect 6288 23276 6368 23304
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6012 18176 6132 18204
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5920 17202 5948 17478
rect 5644 16522 5672 17190
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5736 16794 5764 17138
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4908 15586 4936 16050
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4816 15558 4936 15586
rect 5092 15570 5120 15982
rect 5368 15570 5396 16050
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15706 5488 15846
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5080 15564 5132 15570
rect 4816 15434 4844 15558
rect 5080 15506 5132 15512
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5092 15450 5120 15506
rect 4804 15428 4856 15434
rect 5092 15422 5396 15450
rect 4804 15370 4856 15376
rect 4816 15094 4844 15370
rect 5264 15360 5316 15366
rect 5262 15328 5264 15337
rect 5316 15328 5318 15337
rect 4874 15260 5182 15269
rect 5262 15263 5318 15272
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4724 13938 4752 14486
rect 5368 14482 5396 15422
rect 5552 15162 5580 15982
rect 5644 15706 5672 16458
rect 5828 16046 5856 17138
rect 5920 16726 5948 17138
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5736 15026 5764 15914
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4908 13938 5028 13954
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4896 13932 5028 13938
rect 4948 13926 5028 13932
rect 4896 13874 4948 13880
rect 4436 13806 4488 13812
rect 4618 13832 4674 13841
rect 3976 13796 4028 13802
rect 4618 13767 4674 13776
rect 4804 13796 4856 13802
rect 3976 13738 4028 13744
rect 4804 13738 4856 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4066 12880 4122 12889
rect 4066 12815 4068 12824
rect 4120 12815 4122 12824
rect 4068 12786 4120 12792
rect 3882 12744 3938 12753
rect 4172 12730 4200 13194
rect 4448 12918 4476 13466
rect 4724 13190 4752 13466
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 3882 12679 3938 12688
rect 4080 12702 4200 12730
rect 4540 12714 4568 13126
rect 4816 12968 4844 13738
rect 5000 13394 5028 13926
rect 5368 13530 5396 14214
rect 5552 13938 5580 14894
rect 6012 14414 6040 18176
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6104 15570 6132 16730
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6288 15094 6316 23276
rect 6368 23258 6420 23264
rect 6366 22944 6422 22953
rect 6366 22879 6422 22888
rect 6380 22438 6408 22879
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6472 22080 6500 23530
rect 6564 22710 6592 23695
rect 6656 23594 6684 23820
rect 6644 23588 6696 23594
rect 6644 23530 6696 23536
rect 6642 23352 6698 23361
rect 6642 23287 6698 23296
rect 6656 23186 6684 23287
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6552 22704 6604 22710
rect 6656 22681 6684 22986
rect 6552 22646 6604 22652
rect 6642 22672 6698 22681
rect 6564 22234 6592 22646
rect 6642 22607 6698 22616
rect 6552 22228 6604 22234
rect 6552 22170 6604 22176
rect 6380 22052 6500 22080
rect 6380 21078 6408 22052
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6368 21072 6420 21078
rect 6368 21014 6420 21020
rect 6380 20058 6408 21014
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6380 19922 6408 19994
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6472 17134 6500 21898
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21622 6592 21830
rect 6552 21616 6604 21622
rect 6552 21558 6604 21564
rect 6748 21434 6776 24754
rect 6840 22778 6868 25162
rect 7024 24818 7052 28086
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7012 24676 7064 24682
rect 7012 24618 7064 24624
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6932 24070 6960 24346
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6932 23254 6960 23666
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 6932 22778 6960 23054
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6828 22500 6880 22506
rect 6828 22442 6880 22448
rect 6656 21406 6776 21434
rect 6656 20058 6684 21406
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6748 20942 6776 21286
rect 6840 21146 6868 22442
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6920 21072 6972 21078
rect 6920 21014 6972 21020
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6932 20448 6960 21014
rect 7024 20942 7052 24618
rect 7116 22964 7144 28630
rect 7208 28218 7236 29106
rect 7300 28558 7328 29679
rect 7564 29640 7616 29646
rect 7564 29582 7616 29588
rect 7472 29096 7524 29102
rect 7472 29038 7524 29044
rect 7484 28694 7512 29038
rect 7472 28688 7524 28694
rect 7472 28630 7524 28636
rect 7576 28626 7604 29582
rect 7564 28620 7616 28626
rect 7564 28562 7616 28568
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7380 28552 7432 28558
rect 7380 28494 7432 28500
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 7196 28212 7248 28218
rect 7196 28154 7248 28160
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7208 27713 7236 27950
rect 7194 27704 7250 27713
rect 7194 27639 7250 27648
rect 7208 26994 7236 27639
rect 7300 26994 7328 28358
rect 7392 27538 7420 28494
rect 7472 27668 7524 27674
rect 7472 27610 7524 27616
rect 7380 27532 7432 27538
rect 7380 27474 7432 27480
rect 7484 27010 7512 27610
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 7288 26988 7340 26994
rect 7288 26930 7340 26936
rect 7392 26982 7512 27010
rect 7208 26450 7236 26930
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 7300 26586 7328 26726
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7196 26444 7248 26450
rect 7196 26386 7248 26392
rect 7208 25906 7236 26386
rect 7392 25974 7420 26982
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7484 26586 7512 26862
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7380 25968 7432 25974
rect 7380 25910 7432 25916
rect 7196 25900 7248 25906
rect 7196 25842 7248 25848
rect 7380 25424 7432 25430
rect 7380 25366 7432 25372
rect 7576 25378 7604 28562
rect 7668 26994 7696 30126
rect 7748 29300 7800 29306
rect 7748 29242 7800 29248
rect 7760 29170 7788 29242
rect 7748 29164 7800 29170
rect 7748 29106 7800 29112
rect 7760 28694 7788 29106
rect 7748 28688 7800 28694
rect 7748 28630 7800 28636
rect 7748 28144 7800 28150
rect 7748 28086 7800 28092
rect 7760 27713 7788 28086
rect 7852 27878 7880 30790
rect 7932 30728 7984 30734
rect 7932 30670 7984 30676
rect 8116 30728 8168 30734
rect 8116 30670 8168 30676
rect 7944 30054 7972 30670
rect 8128 30598 8156 30670
rect 8116 30592 8168 30598
rect 8116 30534 8168 30540
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 8116 30048 8168 30054
rect 8116 29990 8168 29996
rect 8128 29646 8156 29990
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 8116 29028 8168 29034
rect 8116 28970 8168 28976
rect 7932 28620 7984 28626
rect 7932 28562 7984 28568
rect 7944 28490 7972 28562
rect 7932 28484 7984 28490
rect 7932 28426 7984 28432
rect 8128 28082 8156 28970
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7746 27704 7802 27713
rect 7746 27639 7748 27648
rect 7800 27639 7802 27648
rect 7748 27610 7800 27616
rect 8036 27402 8064 27950
rect 8128 27878 8156 28018
rect 8116 27872 8168 27878
rect 8116 27814 8168 27820
rect 8024 27396 8076 27402
rect 8024 27338 8076 27344
rect 8116 27396 8168 27402
rect 8116 27338 8168 27344
rect 8036 27305 8064 27338
rect 8022 27296 8078 27305
rect 8022 27231 8078 27240
rect 8128 27130 8156 27338
rect 7932 27124 7984 27130
rect 7932 27066 7984 27072
rect 8116 27124 8168 27130
rect 8116 27066 8168 27072
rect 7656 26988 7708 26994
rect 7656 26930 7708 26936
rect 7668 26586 7696 26930
rect 7656 26580 7708 26586
rect 7656 26522 7708 26528
rect 7840 25968 7892 25974
rect 7840 25910 7892 25916
rect 7852 25702 7880 25910
rect 7840 25696 7892 25702
rect 7838 25664 7840 25673
rect 7892 25664 7894 25673
rect 7838 25599 7894 25608
rect 7392 25294 7420 25366
rect 7576 25350 7788 25378
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7656 25288 7708 25294
rect 7656 25230 7708 25236
rect 7208 24206 7236 25230
rect 7288 24812 7340 24818
rect 7288 24754 7340 24760
rect 7300 24342 7328 24754
rect 7288 24336 7340 24342
rect 7288 24278 7340 24284
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 7208 23662 7236 24142
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7208 23322 7236 23462
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7196 23112 7248 23118
rect 7194 23080 7196 23089
rect 7248 23080 7250 23089
rect 7194 23015 7250 23024
rect 7116 22936 7236 22964
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 7116 22030 7144 22510
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7116 20602 7144 21558
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7012 20460 7064 20466
rect 6932 20420 7012 20448
rect 7012 20402 7064 20408
rect 7024 20369 7052 20402
rect 7010 20360 7066 20369
rect 6920 20324 6972 20330
rect 7010 20295 7066 20304
rect 6920 20266 6972 20272
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6472 16658 6500 17070
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5276 12986 5304 13398
rect 5460 13297 5488 13738
rect 5446 13288 5502 13297
rect 5446 13223 5502 13232
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5264 12980 5316 12986
rect 4816 12940 5120 12968
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4528 12708 4580 12714
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3896 12442 3924 12582
rect 3884 12436 3936 12442
rect 4080 12434 4108 12702
rect 4580 12668 4660 12696
rect 4528 12650 4580 12656
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4252 12436 4304 12442
rect 4080 12406 4200 12434
rect 3884 12378 3936 12384
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3620 12102 3648 12174
rect 4172 12170 4200 12406
rect 4252 12378 4304 12384
rect 4264 12306 4292 12378
rect 4342 12336 4398 12345
rect 4252 12300 4304 12306
rect 4632 12306 4660 12668
rect 4724 12481 4752 12718
rect 4710 12472 4766 12481
rect 4710 12407 4766 12416
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4342 12271 4398 12280
rect 4620 12300 4672 12306
rect 4252 12242 4304 12248
rect 4356 12238 4384 12271
rect 4620 12242 4672 12248
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 4172 11898 4200 12106
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4356 11694 4384 12174
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4632 11898 4660 12106
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3330 10704 3386 10713
rect 3240 10668 3292 10674
rect 3330 10639 3386 10648
rect 3240 10610 3292 10616
rect 3252 10198 3280 10610
rect 3344 10470 3372 10639
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3436 9722 3464 9998
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3528 8090 3556 11562
rect 3620 10674 3648 11630
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4252 11144 4304 11150
rect 4724 11098 4752 12310
rect 4816 12209 4844 12786
rect 4894 12608 4950 12617
rect 4894 12543 4950 12552
rect 4908 12238 4936 12543
rect 4896 12232 4948 12238
rect 4802 12200 4858 12209
rect 5000 12209 5028 12786
rect 4896 12174 4948 12180
rect 4986 12200 5042 12209
rect 4802 12135 4858 12144
rect 4986 12135 5042 12144
rect 4804 12096 4856 12102
rect 5092 12084 5120 12940
rect 5264 12922 5316 12928
rect 5172 12844 5224 12850
rect 5276 12832 5304 12922
rect 5224 12804 5304 12832
rect 5172 12786 5224 12792
rect 5184 12617 5212 12786
rect 5170 12608 5226 12617
rect 5170 12543 5226 12552
rect 5092 12056 5304 12084
rect 4804 12038 4856 12044
rect 4816 11642 4844 12038
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11937 5304 12056
rect 5262 11928 5318 11937
rect 5262 11863 5318 11872
rect 4894 11792 4950 11801
rect 4894 11727 4896 11736
rect 4948 11727 4950 11736
rect 5264 11756 5316 11762
rect 4896 11698 4948 11704
rect 5264 11698 5316 11704
rect 5170 11656 5226 11665
rect 4816 11614 5028 11642
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4252 11086 4304 11092
rect 4264 11014 4292 11086
rect 4632 11070 4752 11098
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 3712 10742 3740 10950
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 4172 10674 4200 10950
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3620 10554 3648 10610
rect 3792 10600 3844 10606
rect 3620 10526 3740 10554
rect 3792 10542 3844 10548
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3620 10130 3648 10406
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3712 9081 3740 10526
rect 3804 10266 3832 10542
rect 3896 10266 3924 10610
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3896 10062 3924 10202
rect 3988 10062 4016 10406
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3976 10056 4028 10062
rect 4080 10044 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4160 10056 4212 10062
rect 4080 10016 4160 10044
rect 3976 9998 4028 10004
rect 4252 10056 4304 10062
rect 4160 9998 4212 10004
rect 4250 10024 4252 10033
rect 4304 10024 4306 10033
rect 4250 9959 4306 9968
rect 3976 9920 4028 9926
rect 3882 9888 3938 9897
rect 3976 9862 4028 9868
rect 3882 9823 3938 9832
rect 3698 9072 3754 9081
rect 3698 9007 3754 9016
rect 3896 8294 3924 9823
rect 3988 9450 4016 9862
rect 4632 9654 4660 11070
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4724 10606 4752 10950
rect 4816 10674 4844 11154
rect 4908 11150 4936 11494
rect 5000 11150 5028 11614
rect 5170 11591 5226 11600
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5184 10996 5212 11591
rect 5276 11286 5304 11698
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 5276 11150 5304 11222
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5184 10968 5304 10996
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 5276 10538 5304 10968
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10198 4936 10406
rect 4896 10192 4948 10198
rect 4710 10160 4766 10169
rect 4896 10134 4948 10140
rect 4710 10095 4766 10104
rect 4724 10062 4752 10095
rect 4908 10062 4936 10134
rect 5368 10130 5396 13126
rect 5460 12646 5488 13126
rect 5552 12832 5580 13874
rect 5644 13172 5672 13874
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5736 13326 5764 13738
rect 5828 13530 5856 13874
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5828 13172 5856 13330
rect 5644 13144 5856 13172
rect 5828 12986 5856 13144
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5816 12844 5868 12850
rect 5552 12804 5816 12832
rect 5816 12786 5868 12792
rect 5538 12744 5594 12753
rect 5538 12679 5594 12688
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5448 12368 5500 12374
rect 5552 12356 5580 12679
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5814 12608 5870 12617
rect 5500 12328 5580 12356
rect 5448 12310 5500 12316
rect 5460 12238 5488 12310
rect 5644 12288 5672 12582
rect 5814 12543 5870 12552
rect 5552 12260 5672 12288
rect 5724 12300 5776 12306
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 11762 5488 12174
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5446 11656 5502 11665
rect 5446 11591 5502 11600
rect 5460 11014 5488 11591
rect 5552 11286 5580 12260
rect 5724 12242 5776 12248
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5644 11762 5672 12106
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 11558 5672 11698
rect 5736 11626 5764 12242
rect 5828 11762 5856 12543
rect 5920 12442 5948 14214
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5920 11898 5948 12378
rect 6012 11898 6040 13194
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6104 11778 6132 14758
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 14074 6408 14214
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6196 12753 6224 13194
rect 6182 12744 6238 12753
rect 6182 12679 6238 12688
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 6012 11750 6132 11778
rect 6196 11762 6224 12582
rect 6288 12434 6316 13806
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6380 12782 6408 13262
rect 6472 12850 6500 16594
rect 6564 14906 6592 19654
rect 6656 18902 6684 19994
rect 6932 19922 6960 20266
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6748 18970 6776 19246
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6656 15366 6684 17614
rect 6736 16652 6788 16658
rect 6840 16640 6868 19722
rect 6932 19446 6960 19858
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6932 18902 6960 19382
rect 7024 18986 7052 20198
rect 7116 19718 7144 20538
rect 7208 20262 7236 22936
rect 7300 20534 7328 24278
rect 7380 24200 7432 24206
rect 7378 24168 7380 24177
rect 7432 24168 7434 24177
rect 7434 24126 7512 24154
rect 7378 24103 7434 24112
rect 7378 23760 7434 23769
rect 7378 23695 7380 23704
rect 7432 23695 7434 23704
rect 7380 23666 7432 23672
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7392 23497 7420 23530
rect 7378 23488 7434 23497
rect 7378 23423 7434 23432
rect 7380 23044 7432 23050
rect 7380 22986 7432 22992
rect 7392 22710 7420 22986
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 7484 22030 7512 24126
rect 7564 23520 7616 23526
rect 7564 23462 7616 23468
rect 7472 22024 7524 22030
rect 7470 21992 7472 22001
rect 7524 21992 7526 22001
rect 7470 21927 7526 21936
rect 7576 21570 7604 23462
rect 7668 22817 7696 25230
rect 7654 22808 7710 22817
rect 7654 22743 7710 22752
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7484 21542 7604 21570
rect 7484 21078 7512 21542
rect 7668 21350 7696 22510
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7472 21072 7524 21078
rect 7656 21072 7708 21078
rect 7472 21014 7524 21020
rect 7576 21020 7656 21026
rect 7576 21014 7708 21020
rect 7576 20998 7696 21014
rect 7576 20806 7604 20998
rect 7656 20936 7708 20942
rect 7760 20924 7788 25350
rect 7944 23848 7972 27066
rect 8116 26308 8168 26314
rect 8116 26250 8168 26256
rect 8024 25288 8076 25294
rect 8024 25230 8076 25236
rect 8036 24886 8064 25230
rect 8024 24880 8076 24886
rect 8024 24822 8076 24828
rect 7944 23820 8064 23848
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7852 22642 7880 22918
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7944 22166 7972 23666
rect 7932 22160 7984 22166
rect 7932 22102 7984 22108
rect 8036 22094 8064 23820
rect 8128 23526 8156 26250
rect 8220 25430 8248 34002
rect 8312 33658 8340 35770
rect 8956 35698 8984 36246
rect 9312 36168 9364 36174
rect 9312 36110 9364 36116
rect 9692 36156 9720 36790
rect 14832 36780 14884 36786
rect 14832 36722 14884 36728
rect 14924 36780 14976 36786
rect 14924 36722 14976 36728
rect 15292 36780 15344 36786
rect 15844 36780 15896 36786
rect 15344 36740 15844 36768
rect 15292 36722 15344 36728
rect 15844 36722 15896 36728
rect 10692 36712 10744 36718
rect 10692 36654 10744 36660
rect 11060 36712 11112 36718
rect 11060 36654 11112 36660
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 13268 36712 13320 36718
rect 13268 36654 13320 36660
rect 14096 36712 14148 36718
rect 14096 36654 14148 36660
rect 14740 36712 14792 36718
rect 14740 36654 14792 36660
rect 9772 36168 9824 36174
rect 9692 36128 9772 36156
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 8944 35692 8996 35698
rect 8996 35652 9076 35680
rect 8944 35634 8996 35640
rect 8576 35488 8628 35494
rect 8576 35430 8628 35436
rect 8588 35086 8616 35430
rect 8772 35290 8800 35634
rect 8944 35556 8996 35562
rect 8944 35498 8996 35504
rect 8760 35284 8812 35290
rect 8760 35226 8812 35232
rect 8956 35086 8984 35498
rect 9048 35154 9076 35652
rect 9324 35290 9352 36110
rect 9588 36100 9640 36106
rect 9588 36042 9640 36048
rect 9600 35630 9628 36042
rect 9692 35766 9720 36128
rect 9772 36110 9824 36116
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 9680 35760 9732 35766
rect 9680 35702 9732 35708
rect 9588 35624 9640 35630
rect 9588 35566 9640 35572
rect 9312 35284 9364 35290
rect 9312 35226 9364 35232
rect 9036 35148 9088 35154
rect 9036 35090 9088 35096
rect 8576 35080 8628 35086
rect 8576 35022 8628 35028
rect 8944 35080 8996 35086
rect 8944 35022 8996 35028
rect 8588 34610 8616 35022
rect 8852 35012 8904 35018
rect 8852 34954 8904 34960
rect 8760 34944 8812 34950
rect 8760 34886 8812 34892
rect 8576 34604 8628 34610
rect 8576 34546 8628 34552
rect 8392 34128 8444 34134
rect 8392 34070 8444 34076
rect 8300 33652 8352 33658
rect 8300 33594 8352 33600
rect 8312 32434 8340 33594
rect 8404 32910 8432 34070
rect 8484 34060 8536 34066
rect 8484 34002 8536 34008
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 8300 32428 8352 32434
rect 8300 32370 8352 32376
rect 8208 25424 8260 25430
rect 8208 25366 8260 25372
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8220 24682 8248 25230
rect 8208 24676 8260 24682
rect 8208 24618 8260 24624
rect 8312 24274 8340 32370
rect 8496 32366 8524 34002
rect 8576 33312 8628 33318
rect 8576 33254 8628 33260
rect 8484 32360 8536 32366
rect 8484 32302 8536 32308
rect 8392 32292 8444 32298
rect 8392 32234 8444 32240
rect 8404 31890 8432 32234
rect 8482 32056 8538 32065
rect 8482 31991 8538 32000
rect 8392 31884 8444 31890
rect 8392 31826 8444 31832
rect 8496 31346 8524 31991
rect 8484 31340 8536 31346
rect 8484 31282 8536 31288
rect 8588 31249 8616 33254
rect 8772 32978 8800 34886
rect 8864 34542 8892 34954
rect 8956 34610 8984 35022
rect 9048 34746 9076 35090
rect 9036 34740 9088 34746
rect 9036 34682 9088 34688
rect 9324 34678 9352 35226
rect 9600 35086 9628 35566
rect 9588 35080 9640 35086
rect 9588 35022 9640 35028
rect 9312 34672 9364 34678
rect 9312 34614 9364 34620
rect 9404 34672 9456 34678
rect 9404 34614 9456 34620
rect 8944 34604 8996 34610
rect 8944 34546 8996 34552
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8864 33425 8892 34478
rect 8956 34134 8984 34546
rect 8944 34128 8996 34134
rect 8944 34070 8996 34076
rect 9128 34128 9180 34134
rect 9128 34070 9180 34076
rect 8850 33416 8906 33425
rect 8850 33351 8906 33360
rect 8760 32972 8812 32978
rect 8760 32914 8812 32920
rect 8760 32836 8812 32842
rect 8864 32824 8892 33351
rect 8812 32796 8892 32824
rect 8760 32778 8812 32784
rect 8772 32042 8800 32778
rect 9036 32496 9088 32502
rect 9036 32438 9088 32444
rect 8852 32224 8904 32230
rect 8904 32184 8984 32212
rect 8852 32166 8904 32172
rect 8772 32014 8892 32042
rect 8864 31736 8892 32014
rect 8956 31890 8984 32184
rect 8944 31884 8996 31890
rect 8944 31826 8996 31832
rect 8772 31708 8892 31736
rect 8668 31680 8720 31686
rect 8668 31622 8720 31628
rect 8574 31240 8630 31249
rect 8574 31175 8576 31184
rect 8628 31175 8630 31184
rect 8576 31146 8628 31152
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 8496 30938 8524 31078
rect 8680 30938 8708 31622
rect 8484 30932 8536 30938
rect 8484 30874 8536 30880
rect 8668 30932 8720 30938
rect 8668 30874 8720 30880
rect 8668 30796 8720 30802
rect 8668 30738 8720 30744
rect 8576 30184 8628 30190
rect 8576 30126 8628 30132
rect 8392 30048 8444 30054
rect 8392 29990 8444 29996
rect 8404 29714 8432 29990
rect 8392 29708 8444 29714
rect 8392 29650 8444 29656
rect 8588 28762 8616 30126
rect 8680 29646 8708 30738
rect 8668 29640 8720 29646
rect 8668 29582 8720 29588
rect 8668 29164 8720 29170
rect 8668 29106 8720 29112
rect 8576 28756 8628 28762
rect 8576 28698 8628 28704
rect 8392 26512 8444 26518
rect 8392 26454 8444 26460
rect 8404 26353 8432 26454
rect 8390 26344 8446 26353
rect 8390 26279 8446 26288
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 8496 25430 8524 25842
rect 8484 25424 8536 25430
rect 8484 25366 8536 25372
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8496 24750 8524 25230
rect 8588 24834 8616 28698
rect 8680 28558 8708 29106
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 8588 24806 8708 24834
rect 8484 24744 8536 24750
rect 8484 24686 8536 24692
rect 8576 24676 8628 24682
rect 8576 24618 8628 24624
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8312 23730 8340 24210
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8114 23352 8170 23361
rect 8114 23287 8170 23296
rect 8128 22710 8156 23287
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 8220 22778 8248 23122
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8116 22704 8168 22710
rect 8116 22646 8168 22652
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8116 22568 8168 22574
rect 8116 22510 8168 22516
rect 8128 22409 8156 22510
rect 8220 22438 8248 22578
rect 8208 22432 8260 22438
rect 8114 22400 8170 22409
rect 8208 22374 8260 22380
rect 8114 22335 8170 22344
rect 8036 22066 8156 22094
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 7840 20936 7892 20942
rect 7760 20904 7840 20924
rect 7892 20904 7894 20913
rect 7760 20896 7838 20904
rect 7656 20878 7708 20884
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7208 19174 7236 20198
rect 7300 19922 7328 20334
rect 7484 20262 7512 20538
rect 7668 20398 7696 20878
rect 7838 20839 7894 20848
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7392 20058 7420 20198
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19514 7328 19654
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7024 18958 7328 18986
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6932 17270 6960 18838
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 7024 17134 7052 18770
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7116 17882 7144 18294
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17338 7236 17478
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6840 16612 6960 16640
rect 6736 16594 6788 16600
rect 6748 16182 6776 16594
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 6748 15638 6776 16118
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6564 14878 6776 14906
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6564 13938 6592 14758
rect 6656 14006 6684 14758
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6748 13802 6776 14878
rect 6840 14414 6868 14962
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6840 14074 6868 14350
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13530 6776 13738
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6564 13326 6592 13398
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6840 13258 6868 14010
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6932 12986 6960 16612
rect 7024 16153 7052 17070
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7010 16144 7066 16153
rect 7010 16079 7066 16088
rect 7116 15706 7144 16526
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7208 15706 7236 15982
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7300 14482 7328 18958
rect 7576 18426 7604 19450
rect 7760 18578 7788 20742
rect 7944 20398 7972 21966
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 8036 21418 8064 21898
rect 8024 21412 8076 21418
rect 8024 21354 8076 21360
rect 8128 20890 8156 22066
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8036 20862 8156 20890
rect 8036 20534 8064 20862
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 8128 20602 8156 20742
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 8114 20496 8170 20505
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7932 19440 7984 19446
rect 7838 19408 7894 19417
rect 7932 19382 7984 19388
rect 7838 19343 7894 19352
rect 7668 18550 7788 18578
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13938 7328 14214
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7392 13394 7420 18022
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7576 17270 7604 17478
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7576 15502 7604 16390
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7484 15026 7512 15370
rect 7668 15042 7696 18550
rect 7746 18456 7802 18465
rect 7852 18426 7880 19343
rect 7746 18391 7748 18400
rect 7800 18391 7802 18400
rect 7840 18420 7892 18426
rect 7748 18362 7800 18368
rect 7840 18362 7892 18368
rect 7760 17610 7788 18362
rect 7944 17678 7972 19382
rect 8036 18766 8064 20470
rect 8220 20466 8248 22034
rect 8312 22030 8340 23666
rect 8390 23216 8446 23225
rect 8390 23151 8446 23160
rect 8404 23118 8432 23151
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8312 21622 8340 21966
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8404 21554 8432 23054
rect 8484 23044 8536 23050
rect 8484 22986 8536 22992
rect 8496 22098 8524 22986
rect 8588 22982 8616 24618
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 8484 22092 8536 22098
rect 8484 22034 8536 22040
rect 8482 21992 8538 22001
rect 8588 21962 8616 22442
rect 8680 22137 8708 24806
rect 8772 24721 8800 31708
rect 8956 31346 8984 31826
rect 9048 31754 9076 32438
rect 9036 31748 9088 31754
rect 9036 31690 9088 31696
rect 9140 31686 9168 34070
rect 9416 34066 9444 34614
rect 9496 34196 9548 34202
rect 9496 34138 9548 34144
rect 9508 34066 9536 34138
rect 9404 34060 9456 34066
rect 9404 34002 9456 34008
rect 9496 34060 9548 34066
rect 9496 34002 9548 34008
rect 9496 33856 9548 33862
rect 9496 33798 9548 33804
rect 9404 33652 9456 33658
rect 9324 33612 9404 33640
rect 9220 31816 9272 31822
rect 9220 31758 9272 31764
rect 9128 31680 9180 31686
rect 9128 31622 9180 31628
rect 9140 31346 9168 31622
rect 9232 31482 9260 31758
rect 9220 31476 9272 31482
rect 9220 31418 9272 31424
rect 8944 31340 8996 31346
rect 9128 31340 9180 31346
rect 8996 31300 9076 31328
rect 8944 31282 8996 31288
rect 9048 31142 9076 31300
rect 9128 31282 9180 31288
rect 9220 31340 9272 31346
rect 9220 31282 9272 31288
rect 9140 31210 9168 31282
rect 9128 31204 9180 31210
rect 9128 31146 9180 31152
rect 9036 31136 9088 31142
rect 9036 31078 9088 31084
rect 8852 30252 8904 30258
rect 8852 30194 8904 30200
rect 8944 30252 8996 30258
rect 8944 30194 8996 30200
rect 8864 30054 8892 30194
rect 8852 30048 8904 30054
rect 8852 29990 8904 29996
rect 8956 29850 8984 30194
rect 8944 29844 8996 29850
rect 8944 29786 8996 29792
rect 9048 28994 9076 31078
rect 9126 30968 9182 30977
rect 9232 30938 9260 31282
rect 9126 30903 9182 30912
rect 9220 30932 9272 30938
rect 9140 30784 9168 30903
rect 9220 30874 9272 30880
rect 9324 30802 9352 33612
rect 9404 33594 9456 33600
rect 9404 33448 9456 33454
rect 9402 33416 9404 33425
rect 9456 33416 9458 33425
rect 9508 33386 9536 33798
rect 9692 33674 9720 35702
rect 9772 35692 9824 35698
rect 9772 35634 9824 35640
rect 9784 34746 9812 35634
rect 9876 35018 9904 36110
rect 10416 36100 10468 36106
rect 10416 36042 10468 36048
rect 10140 36032 10192 36038
rect 10140 35974 10192 35980
rect 10152 35698 10180 35974
rect 10428 35834 10456 36042
rect 10416 35828 10468 35834
rect 10416 35770 10468 35776
rect 10140 35692 10192 35698
rect 10140 35634 10192 35640
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 10244 35086 10272 35430
rect 10704 35086 10732 36654
rect 11072 35834 11100 36654
rect 12636 36310 12664 36654
rect 12716 36576 12768 36582
rect 12716 36518 12768 36524
rect 12624 36304 12676 36310
rect 12624 36246 12676 36252
rect 12624 36168 12676 36174
rect 12624 36110 12676 36116
rect 12164 36100 12216 36106
rect 12164 36042 12216 36048
rect 11060 35828 11112 35834
rect 11060 35770 11112 35776
rect 10876 35692 10928 35698
rect 10876 35634 10928 35640
rect 10784 35624 10836 35630
rect 10784 35566 10836 35572
rect 10232 35080 10284 35086
rect 10232 35022 10284 35028
rect 10692 35080 10744 35086
rect 10692 35022 10744 35028
rect 10796 35034 10824 35566
rect 10888 35290 10916 35634
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 11980 35624 12032 35630
rect 11980 35566 12032 35572
rect 10876 35284 10928 35290
rect 10876 35226 10928 35232
rect 10980 35222 11008 35566
rect 11060 35556 11112 35562
rect 11060 35498 11112 35504
rect 11428 35556 11480 35562
rect 11428 35498 11480 35504
rect 10968 35216 11020 35222
rect 10968 35158 11020 35164
rect 10968 35080 11020 35086
rect 10796 35028 10968 35034
rect 10796 35022 11020 35028
rect 9864 35012 9916 35018
rect 9864 34954 9916 34960
rect 10704 34746 10732 35022
rect 10796 35006 11008 35022
rect 9772 34740 9824 34746
rect 9772 34682 9824 34688
rect 10692 34740 10744 34746
rect 10692 34682 10744 34688
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 9876 34202 9904 34546
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 9956 34060 10008 34066
rect 9956 34002 10008 34008
rect 10692 34060 10744 34066
rect 10692 34002 10744 34008
rect 9600 33646 9904 33674
rect 9600 33590 9628 33646
rect 9588 33584 9640 33590
rect 9588 33526 9640 33532
rect 9680 33584 9732 33590
rect 9680 33526 9732 33532
rect 9402 33351 9458 33360
rect 9496 33380 9548 33386
rect 9496 33322 9548 33328
rect 9404 33312 9456 33318
rect 9404 33254 9456 33260
rect 9312 30796 9364 30802
rect 9140 30756 9260 30784
rect 9128 30320 9180 30326
rect 9126 30288 9128 30297
rect 9180 30288 9182 30297
rect 9126 30223 9182 30232
rect 9232 29850 9260 30756
rect 9312 30738 9364 30744
rect 9310 29880 9366 29889
rect 9220 29844 9272 29850
rect 9310 29815 9366 29824
rect 9220 29786 9272 29792
rect 9128 29776 9180 29782
rect 9126 29744 9128 29753
rect 9180 29744 9182 29753
rect 9126 29679 9182 29688
rect 9324 29646 9352 29815
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9220 29504 9272 29510
rect 9220 29446 9272 29452
rect 9232 29170 9260 29446
rect 9416 29238 9444 33254
rect 9508 32910 9536 33322
rect 9692 32978 9720 33526
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9496 32904 9548 32910
rect 9548 32852 9720 32858
rect 9496 32846 9720 32852
rect 9508 32830 9720 32846
rect 9692 32416 9720 32830
rect 9772 32836 9824 32842
rect 9772 32778 9824 32784
rect 9784 32609 9812 32778
rect 9770 32600 9826 32609
rect 9876 32570 9904 33646
rect 9968 33130 9996 34002
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 9968 33102 10180 33130
rect 10244 33114 10272 33934
rect 10416 33856 10468 33862
rect 10416 33798 10468 33804
rect 10598 33824 10654 33833
rect 10428 33522 10456 33798
rect 10598 33759 10654 33768
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10428 33386 10456 33458
rect 10416 33380 10468 33386
rect 10416 33322 10468 33328
rect 9968 32774 9996 33102
rect 10152 33046 10180 33102
rect 10232 33108 10284 33114
rect 10232 33050 10284 33056
rect 10048 33040 10100 33046
rect 10048 32982 10100 32988
rect 10140 33040 10192 33046
rect 10140 32982 10192 32988
rect 9956 32768 10008 32774
rect 9956 32710 10008 32716
rect 9770 32535 9826 32544
rect 9864 32564 9916 32570
rect 9864 32506 9916 32512
rect 9692 32388 9904 32416
rect 9496 32360 9548 32366
rect 9496 32302 9548 32308
rect 9588 32360 9640 32366
rect 9588 32302 9640 32308
rect 9770 32328 9826 32337
rect 9508 31770 9536 32302
rect 9600 32065 9628 32302
rect 9770 32263 9826 32272
rect 9586 32056 9642 32065
rect 9586 31991 9642 32000
rect 9600 31958 9628 31991
rect 9588 31952 9640 31958
rect 9588 31894 9640 31900
rect 9678 31920 9734 31929
rect 9678 31855 9680 31864
rect 9732 31855 9734 31864
rect 9680 31826 9732 31832
rect 9784 31822 9812 32263
rect 9588 31816 9640 31822
rect 9508 31764 9588 31770
rect 9508 31758 9640 31764
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9508 31742 9628 31758
rect 9508 31346 9536 31742
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9496 31340 9548 31346
rect 9496 31282 9548 31288
rect 9692 30870 9720 31418
rect 9784 31210 9812 31758
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9680 30864 9732 30870
rect 9494 30832 9550 30841
rect 9680 30806 9732 30812
rect 9494 30767 9550 30776
rect 9508 30666 9536 30767
rect 9588 30728 9640 30734
rect 9588 30670 9640 30676
rect 9496 30660 9548 30666
rect 9496 30602 9548 30608
rect 9600 30190 9628 30670
rect 9588 30184 9640 30190
rect 9586 30152 9588 30161
rect 9640 30152 9642 30161
rect 9586 30087 9642 30096
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 9496 29504 9548 29510
rect 9496 29446 9548 29452
rect 9404 29232 9456 29238
rect 9404 29174 9456 29180
rect 9220 29164 9272 29170
rect 9220 29106 9272 29112
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 8956 28966 9076 28994
rect 8852 28076 8904 28082
rect 8852 28018 8904 28024
rect 8864 25430 8892 28018
rect 8852 25424 8904 25430
rect 8852 25366 8904 25372
rect 8850 24848 8906 24857
rect 8850 24783 8906 24792
rect 8864 24750 8892 24783
rect 8852 24744 8904 24750
rect 8758 24712 8814 24721
rect 8852 24686 8904 24692
rect 8758 24647 8814 24656
rect 8772 23118 8800 24647
rect 8956 23866 8984 28966
rect 9220 28688 9272 28694
rect 9220 28630 9272 28636
rect 9232 28558 9260 28630
rect 9416 28558 9444 29038
rect 9220 28552 9272 28558
rect 9220 28494 9272 28500
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9048 27606 9076 28018
rect 9036 27600 9088 27606
rect 9036 27542 9088 27548
rect 9140 27470 9168 28358
rect 9324 28150 9352 28358
rect 9312 28144 9364 28150
rect 9312 28086 9364 28092
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 9232 27538 9260 28018
rect 9416 27577 9444 28494
rect 9402 27568 9458 27577
rect 9220 27532 9272 27538
rect 9402 27503 9458 27512
rect 9220 27474 9272 27480
rect 9508 27470 9536 29446
rect 9600 29170 9628 29990
rect 9772 29708 9824 29714
rect 9772 29650 9824 29656
rect 9588 29164 9640 29170
rect 9588 29106 9640 29112
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9600 28082 9628 28902
rect 9784 28694 9812 29650
rect 9772 28688 9824 28694
rect 9772 28630 9824 28636
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9692 28218 9720 28494
rect 9784 28218 9812 28494
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 9770 28112 9826 28121
rect 9588 28076 9640 28082
rect 9770 28047 9772 28056
rect 9588 28018 9640 28024
rect 9824 28047 9826 28056
rect 9772 28018 9824 28024
rect 9600 27878 9628 28018
rect 9680 28008 9732 28014
rect 9678 27976 9680 27985
rect 9732 27976 9734 27985
rect 9678 27911 9734 27920
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9496 27464 9548 27470
rect 9496 27406 9548 27412
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9508 27130 9536 27406
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9036 26784 9088 26790
rect 9036 26726 9088 26732
rect 9048 26450 9076 26726
rect 9036 26444 9088 26450
rect 9036 26386 9088 26392
rect 9036 25424 9088 25430
rect 9036 25366 9088 25372
rect 9048 25226 9076 25366
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 9048 24614 9076 24754
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 8944 23860 8996 23866
rect 8996 23820 9076 23848
rect 8944 23802 8996 23808
rect 9048 23202 9076 23820
rect 9140 23798 9168 26930
rect 9600 26858 9628 27406
rect 9588 26852 9640 26858
rect 9588 26794 9640 26800
rect 9600 26382 9628 26794
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9496 26240 9548 26246
rect 9416 26200 9496 26228
rect 9416 25974 9444 26200
rect 9496 26182 9548 26188
rect 9404 25968 9456 25974
rect 9404 25910 9456 25916
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 9508 25786 9536 25842
rect 9324 25758 9536 25786
rect 9588 25764 9640 25770
rect 9324 25702 9352 25758
rect 9588 25706 9640 25712
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 9496 25696 9548 25702
rect 9496 25638 9548 25644
rect 9220 24948 9272 24954
rect 9220 24890 9272 24896
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 8864 23174 9076 23202
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8772 22166 8800 22918
rect 8760 22160 8812 22166
rect 8666 22128 8722 22137
rect 8760 22102 8812 22108
rect 8666 22063 8722 22072
rect 8482 21927 8538 21936
rect 8576 21956 8628 21962
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8392 21004 8444 21010
rect 8392 20946 8444 20952
rect 8298 20632 8354 20641
rect 8298 20567 8354 20576
rect 8114 20431 8170 20440
rect 8208 20460 8260 20466
rect 8128 20398 8156 20431
rect 8208 20402 8260 20408
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8220 19990 8248 20402
rect 8208 19984 8260 19990
rect 8208 19926 8260 19932
rect 8312 19378 8340 20567
rect 8404 20058 8432 20946
rect 8496 20058 8524 21927
rect 8772 21944 8800 22102
rect 8576 21898 8628 21904
rect 8680 21916 8800 21944
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8588 20874 8616 21626
rect 8680 21554 8708 21916
rect 8864 21842 8892 23174
rect 9140 22710 9168 23258
rect 9128 22704 9180 22710
rect 9034 22672 9090 22681
rect 9128 22646 9180 22652
rect 9034 22607 9036 22616
rect 9088 22607 9090 22616
rect 9036 22578 9088 22584
rect 9126 22536 9182 22545
rect 9126 22471 9128 22480
rect 9180 22471 9182 22480
rect 9128 22442 9180 22448
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8772 21814 8892 21842
rect 8772 21554 8800 21814
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8956 21010 8984 22034
rect 9036 21072 9088 21078
rect 9036 21014 9088 21020
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8576 20868 8628 20874
rect 8760 20868 8812 20874
rect 8628 20828 8708 20856
rect 8576 20810 8628 20816
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8404 19938 8432 19994
rect 8404 19910 8616 19938
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7944 17338 7972 17614
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8036 15502 8064 18702
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8128 15094 8156 15846
rect 8220 15706 8248 19314
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8312 16454 8340 19178
rect 8404 18834 8432 19382
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 18290 8432 18566
rect 8496 18426 8524 19790
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8588 18290 8616 19910
rect 8680 19553 8708 20828
rect 8760 20810 8812 20816
rect 8666 19544 8722 19553
rect 8666 19479 8722 19488
rect 8772 19242 8800 20810
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8956 20534 8984 20742
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8942 19952 8998 19961
rect 8852 19916 8904 19922
rect 8942 19887 8998 19896
rect 8852 19858 8904 19864
rect 8864 19786 8892 19858
rect 8956 19854 8984 19887
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8852 19780 8904 19786
rect 8852 19722 8904 19728
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8758 19136 8814 19145
rect 8680 18290 8708 19110
rect 8758 19071 8814 19080
rect 8772 18970 8800 19071
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8772 18766 8800 18906
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8864 18630 8892 19722
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8956 19417 8984 19654
rect 8942 19408 8998 19417
rect 8942 19343 8998 19352
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8404 18086 8432 18226
rect 8864 18222 8892 18566
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8852 18216 8904 18222
rect 8482 18184 8538 18193
rect 8852 18158 8904 18164
rect 8482 18119 8538 18128
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8496 17746 8524 18119
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8404 15570 8432 16662
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8496 16250 8524 16526
rect 8588 16522 8616 17682
rect 8864 17202 8892 18158
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8956 16590 8984 18226
rect 9048 17814 9076 21014
rect 9128 20800 9180 20806
rect 9128 20742 9180 20748
rect 9140 20505 9168 20742
rect 9126 20496 9182 20505
rect 9126 20431 9182 20440
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9140 19854 9168 19994
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9232 19718 9260 24890
rect 9324 24886 9352 25638
rect 9416 25498 9444 25638
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 9508 25378 9536 25638
rect 9416 25350 9536 25378
rect 9416 25294 9444 25350
rect 9600 25294 9628 25706
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9588 25288 9640 25294
rect 9588 25230 9640 25236
rect 9312 24880 9364 24886
rect 9312 24822 9364 24828
rect 9416 24818 9444 25230
rect 9600 24818 9628 25230
rect 9404 24812 9456 24818
rect 9404 24754 9456 24760
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9692 24698 9720 27814
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9784 25702 9812 25910
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9784 25294 9812 25434
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9508 24670 9720 24698
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9324 19854 9352 23734
rect 9402 23352 9458 23361
rect 9402 23287 9458 23296
rect 9416 22982 9444 23287
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9416 22574 9444 22918
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9404 21004 9456 21010
rect 9508 20992 9536 24670
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9692 24138 9720 24550
rect 9770 24304 9826 24313
rect 9770 24239 9826 24248
rect 9784 24206 9812 24239
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9588 24132 9640 24138
rect 9588 24074 9640 24080
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 9600 23497 9628 24074
rect 9784 23633 9812 24142
rect 9770 23624 9826 23633
rect 9770 23559 9826 23568
rect 9586 23488 9642 23497
rect 9586 23423 9642 23432
rect 9586 23216 9642 23225
rect 9586 23151 9588 23160
rect 9640 23151 9642 23160
rect 9588 23122 9640 23128
rect 9600 22624 9628 23122
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9680 22636 9732 22642
rect 9600 22596 9680 22624
rect 9680 22578 9732 22584
rect 9784 22386 9812 22646
rect 9876 22386 9904 32388
rect 10060 31890 10088 32982
rect 10232 32972 10284 32978
rect 10232 32914 10284 32920
rect 10244 32858 10272 32914
rect 10152 32830 10272 32858
rect 10324 32904 10376 32910
rect 10324 32846 10376 32852
rect 10152 31958 10180 32830
rect 10232 32768 10284 32774
rect 10232 32710 10284 32716
rect 10244 32026 10272 32710
rect 10336 32366 10364 32846
rect 10428 32842 10456 33322
rect 10508 32904 10560 32910
rect 10508 32846 10560 32852
rect 10416 32836 10468 32842
rect 10416 32778 10468 32784
rect 10324 32360 10376 32366
rect 10324 32302 10376 32308
rect 10428 32212 10456 32778
rect 10336 32184 10456 32212
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10140 31952 10192 31958
rect 10140 31894 10192 31900
rect 10048 31884 10100 31890
rect 10048 31826 10100 31832
rect 9956 31680 10008 31686
rect 9956 31622 10008 31628
rect 9968 31346 9996 31622
rect 10060 31482 10088 31826
rect 10140 31680 10192 31686
rect 10140 31622 10192 31628
rect 10048 31476 10100 31482
rect 10048 31418 10100 31424
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 10152 31278 10180 31622
rect 10140 31272 10192 31278
rect 10140 31214 10192 31220
rect 10152 30394 10180 31214
rect 10232 30796 10284 30802
rect 10232 30738 10284 30744
rect 10140 30388 10192 30394
rect 10140 30330 10192 30336
rect 10244 30326 10272 30738
rect 10232 30320 10284 30326
rect 10232 30262 10284 30268
rect 10244 29510 10272 30262
rect 10232 29504 10284 29510
rect 10230 29472 10232 29481
rect 10284 29472 10286 29481
rect 10230 29407 10286 29416
rect 10336 29238 10364 32184
rect 10520 31278 10548 32846
rect 10612 32502 10640 33759
rect 10704 33658 10732 34002
rect 10874 33960 10930 33969
rect 10874 33895 10930 33904
rect 10692 33652 10744 33658
rect 10692 33594 10744 33600
rect 10600 32496 10652 32502
rect 10600 32438 10652 32444
rect 10600 32020 10652 32026
rect 10600 31962 10652 31968
rect 10612 31822 10640 31962
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10888 31414 10916 33895
rect 10980 33114 11008 35006
rect 11072 34950 11100 35498
rect 11336 35148 11388 35154
rect 11336 35090 11388 35096
rect 11060 34944 11112 34950
rect 11060 34886 11112 34892
rect 11348 34610 11376 35090
rect 11440 35086 11468 35498
rect 11612 35488 11664 35494
rect 11612 35430 11664 35436
rect 11624 35086 11652 35430
rect 11992 35290 12020 35566
rect 11980 35284 12032 35290
rect 11980 35226 12032 35232
rect 11428 35080 11480 35086
rect 11428 35022 11480 35028
rect 11520 35080 11572 35086
rect 11520 35022 11572 35028
rect 11612 35080 11664 35086
rect 11612 35022 11664 35028
rect 11336 34604 11388 34610
rect 11336 34546 11388 34552
rect 11532 34202 11560 35022
rect 12176 34950 12204 36042
rect 12440 35828 12492 35834
rect 12440 35770 12492 35776
rect 12164 34944 12216 34950
rect 12164 34886 12216 34892
rect 12452 34746 12480 35770
rect 12636 34746 12664 36110
rect 12440 34740 12492 34746
rect 12440 34682 12492 34688
rect 12624 34740 12676 34746
rect 12624 34682 12676 34688
rect 12728 34626 12756 36518
rect 13280 36378 13308 36654
rect 13636 36576 13688 36582
rect 13636 36518 13688 36524
rect 13648 36378 13676 36518
rect 13268 36372 13320 36378
rect 13268 36314 13320 36320
rect 13636 36372 13688 36378
rect 13636 36314 13688 36320
rect 13360 36236 13412 36242
rect 13360 36178 13412 36184
rect 13544 36236 13596 36242
rect 13544 36178 13596 36184
rect 12808 36168 12860 36174
rect 12808 36110 12860 36116
rect 12900 36168 12952 36174
rect 12900 36110 12952 36116
rect 12992 36168 13044 36174
rect 13176 36168 13228 36174
rect 13044 36128 13124 36156
rect 12992 36110 13044 36116
rect 12820 35834 12848 36110
rect 12912 35834 12940 36110
rect 12808 35828 12860 35834
rect 12808 35770 12860 35776
rect 12900 35828 12952 35834
rect 12900 35770 12952 35776
rect 12808 35692 12860 35698
rect 12808 35634 12860 35640
rect 12900 35692 12952 35698
rect 12900 35634 12952 35640
rect 12992 35692 13044 35698
rect 12992 35634 13044 35640
rect 12820 34746 12848 35634
rect 12912 35154 12940 35634
rect 12900 35148 12952 35154
rect 12900 35090 12952 35096
rect 12808 34740 12860 34746
rect 12808 34682 12860 34688
rect 12164 34604 12216 34610
rect 12164 34546 12216 34552
rect 12440 34604 12492 34610
rect 12440 34546 12492 34552
rect 12532 34604 12584 34610
rect 12532 34546 12584 34552
rect 12636 34598 12756 34626
rect 11980 34536 12032 34542
rect 11980 34478 12032 34484
rect 11520 34196 11572 34202
rect 11520 34138 11572 34144
rect 11428 34060 11480 34066
rect 11428 34002 11480 34008
rect 11060 33924 11112 33930
rect 11060 33866 11112 33872
rect 11072 33454 11100 33866
rect 11440 33658 11468 34002
rect 11428 33652 11480 33658
rect 11428 33594 11480 33600
rect 11060 33448 11112 33454
rect 11060 33390 11112 33396
rect 11520 33448 11572 33454
rect 11520 33390 11572 33396
rect 10968 33108 11020 33114
rect 10968 33050 11020 33056
rect 10980 32910 11008 33050
rect 11336 32972 11388 32978
rect 11336 32914 11388 32920
rect 10968 32904 11020 32910
rect 10968 32846 11020 32852
rect 10968 32768 11020 32774
rect 10968 32710 11020 32716
rect 10980 31929 11008 32710
rect 11244 32292 11296 32298
rect 11244 32234 11296 32240
rect 10966 31920 11022 31929
rect 10966 31855 11022 31864
rect 10980 31822 11008 31855
rect 11256 31822 11284 32234
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 11244 31816 11296 31822
rect 11244 31758 11296 31764
rect 11152 31748 11204 31754
rect 11152 31690 11204 31696
rect 10876 31408 10928 31414
rect 10876 31350 10928 31356
rect 10692 31340 10744 31346
rect 10692 31282 10744 31288
rect 10508 31272 10560 31278
rect 10508 31214 10560 31220
rect 10416 30728 10468 30734
rect 10416 30670 10468 30676
rect 10428 29850 10456 30670
rect 10508 30592 10560 30598
rect 10508 30534 10560 30540
rect 10520 29850 10548 30534
rect 10704 30394 10732 31282
rect 11164 30870 11192 31690
rect 11348 31346 11376 32914
rect 11428 32224 11480 32230
rect 11428 32166 11480 32172
rect 11440 31822 11468 32166
rect 11428 31816 11480 31822
rect 11428 31758 11480 31764
rect 11336 31340 11388 31346
rect 11336 31282 11388 31288
rect 11348 31142 11376 31282
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11244 30932 11296 30938
rect 11244 30874 11296 30880
rect 11152 30864 11204 30870
rect 11152 30806 11204 30812
rect 10876 30592 10928 30598
rect 10876 30534 10928 30540
rect 10888 30394 10916 30534
rect 10692 30388 10744 30394
rect 10692 30330 10744 30336
rect 10876 30388 10928 30394
rect 10876 30330 10928 30336
rect 10600 30320 10652 30326
rect 10600 30262 10652 30268
rect 10416 29844 10468 29850
rect 10416 29786 10468 29792
rect 10508 29844 10560 29850
rect 10508 29786 10560 29792
rect 10428 29646 10456 29786
rect 10612 29646 10640 30262
rect 10704 30138 10732 30330
rect 11256 30258 11284 30874
rect 11428 30796 11480 30802
rect 11428 30738 11480 30744
rect 11440 30394 11468 30738
rect 11428 30388 11480 30394
rect 11428 30330 11480 30336
rect 10968 30252 11020 30258
rect 10968 30194 11020 30200
rect 11244 30252 11296 30258
rect 11244 30194 11296 30200
rect 10704 30110 10824 30138
rect 10796 30054 10824 30110
rect 10784 30048 10836 30054
rect 10784 29990 10836 29996
rect 10796 29646 10824 29990
rect 10980 29850 11008 30194
rect 11060 30184 11112 30190
rect 11058 30152 11060 30161
rect 11112 30152 11114 30161
rect 11058 30087 11114 30096
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 10416 29640 10468 29646
rect 10600 29640 10652 29646
rect 10468 29600 10548 29628
rect 10416 29582 10468 29588
rect 10324 29232 10376 29238
rect 10324 29174 10376 29180
rect 9956 29164 10008 29170
rect 9956 29106 10008 29112
rect 9968 28762 9996 29106
rect 10048 29028 10100 29034
rect 10048 28970 10100 28976
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 10060 28642 10088 28970
rect 10140 28756 10192 28762
rect 10140 28698 10192 28704
rect 9968 28614 10088 28642
rect 9968 24750 9996 28614
rect 10048 27940 10100 27946
rect 10048 27882 10100 27888
rect 10060 27674 10088 27882
rect 10048 27668 10100 27674
rect 10048 27610 10100 27616
rect 10152 25974 10180 28698
rect 10232 28688 10284 28694
rect 10232 28630 10284 28636
rect 10324 28688 10376 28694
rect 10324 28630 10376 28636
rect 10244 28490 10272 28630
rect 10336 28558 10364 28630
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10232 28484 10284 28490
rect 10232 28426 10284 28432
rect 10336 28082 10364 28494
rect 10416 28212 10468 28218
rect 10416 28154 10468 28160
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 10324 28076 10376 28082
rect 10324 28018 10376 28024
rect 10244 27674 10272 28018
rect 10232 27668 10284 27674
rect 10232 27610 10284 27616
rect 10428 27470 10456 28154
rect 10416 27464 10468 27470
rect 10416 27406 10468 27412
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 10140 25968 10192 25974
rect 10140 25910 10192 25916
rect 10230 25528 10286 25537
rect 10140 25492 10192 25498
rect 10230 25463 10286 25472
rect 10140 25434 10192 25440
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9968 24206 9996 24550
rect 10060 24342 10088 25230
rect 10048 24336 10100 24342
rect 10048 24278 10100 24284
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 9784 22358 9904 22386
rect 9678 22264 9734 22273
rect 9678 22199 9680 22208
rect 9732 22199 9734 22208
rect 9680 22170 9732 22176
rect 9784 22094 9812 22358
rect 9968 22234 9996 22918
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 10060 22273 10088 22714
rect 10046 22264 10102 22273
rect 9956 22228 10008 22234
rect 10046 22199 10102 22208
rect 9956 22170 10008 22176
rect 9784 22066 9904 22094
rect 9772 21956 9824 21962
rect 9772 21898 9824 21904
rect 9784 21622 9812 21898
rect 9772 21616 9824 21622
rect 9456 20964 9536 20992
rect 9404 20946 9456 20952
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 9416 20602 9444 20810
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9402 20360 9458 20369
rect 9402 20295 9458 20304
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9416 19786 9444 20295
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9126 19544 9182 19553
rect 9126 19479 9182 19488
rect 9402 19544 9458 19553
rect 9402 19479 9458 19488
rect 9140 18306 9168 19479
rect 9310 19408 9366 19417
rect 9416 19378 9444 19479
rect 9310 19343 9366 19352
rect 9404 19372 9456 19378
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9232 18834 9260 19246
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9232 18426 9260 18634
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9140 18278 9260 18306
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9036 17808 9088 17814
rect 9036 17750 9088 17756
rect 9140 17678 9168 18090
rect 9232 18086 9260 18278
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8576 16516 8628 16522
rect 8576 16458 8628 16464
rect 8956 16454 8984 16526
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 9048 16250 9076 17546
rect 9232 17513 9260 18022
rect 9324 17542 9352 19343
rect 9404 19314 9456 19320
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9312 17536 9364 17542
rect 9218 17504 9274 17513
rect 9312 17478 9364 17484
rect 9218 17439 9274 17448
rect 9324 17338 9352 17478
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9324 16658 9352 17274
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8496 15502 8524 16186
rect 8574 15600 8630 15609
rect 8574 15535 8630 15544
rect 8588 15502 8616 15535
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8116 15088 8168 15094
rect 7472 15020 7524 15026
rect 7668 15014 7788 15042
rect 8116 15030 8168 15036
rect 7472 14962 7524 14968
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7484 14074 7512 14282
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6644 12912 6696 12918
rect 7024 12866 7052 13262
rect 6644 12854 6696 12860
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6288 12406 6408 12434
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6288 11830 6316 12038
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6184 11756 6236 11762
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10810 5580 10950
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 4080 8974 4108 9522
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4356 8634 4384 9114
rect 4632 8906 4660 9590
rect 4724 9042 4752 9862
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4986 9616 5042 9625
rect 4986 9551 4988 9560
rect 5040 9551 5042 9560
rect 5264 9580 5316 9586
rect 4988 9522 5040 9528
rect 5368 9568 5396 10066
rect 5460 9704 5488 10746
rect 5644 9994 5672 11018
rect 5736 9994 5764 11086
rect 5920 11082 5948 11630
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 5816 10736 5868 10742
rect 5814 10704 5816 10713
rect 5868 10704 5870 10713
rect 5814 10639 5870 10648
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5644 9722 5672 9930
rect 5632 9716 5684 9722
rect 5460 9676 5580 9704
rect 5316 9540 5396 9568
rect 5446 9616 5502 9625
rect 5446 9551 5448 9560
rect 5264 9522 5316 9528
rect 5500 9551 5502 9560
rect 5448 9522 5500 9528
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4816 8974 4844 9318
rect 4908 9217 4936 9386
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 4894 9208 4950 9217
rect 4894 9143 4950 9152
rect 4894 9072 4950 9081
rect 4894 9007 4896 9016
rect 4948 9007 4950 9016
rect 4896 8978 4948 8984
rect 5184 8974 5212 9318
rect 4804 8968 4856 8974
rect 4710 8936 4766 8945
rect 4620 8900 4672 8906
rect 4804 8910 4856 8916
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 4710 8871 4766 8880
rect 5356 8900 5408 8906
rect 4620 8842 4672 8848
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4540 8498 4568 8774
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4448 8401 4476 8434
rect 4434 8392 4490 8401
rect 4434 8327 4490 8336
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2976 7002 3004 7414
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 3528 6905 3556 8026
rect 4632 8022 4660 8570
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4724 7834 4752 8871
rect 5356 8842 5408 8848
rect 4988 8832 5040 8838
rect 4816 8792 4988 8820
rect 4816 7886 4844 8792
rect 4988 8774 5040 8780
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8634 5304 8774
rect 5368 8634 5396 8842
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4896 8560 4948 8566
rect 4894 8528 4896 8537
rect 4948 8528 4950 8537
rect 4894 8463 4950 8472
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5172 8492 5224 8498
rect 5224 8452 5304 8480
rect 5172 8434 5224 8440
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4632 7806 4752 7834
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4908 7818 4936 8366
rect 5092 8294 5120 8434
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4896 7812 4948 7818
rect 4160 7744 4212 7750
rect 4632 7732 4660 7806
rect 4896 7754 4948 7760
rect 5092 7750 5120 8230
rect 4160 7686 4212 7692
rect 4540 7704 4660 7732
rect 4712 7744 4764 7750
rect 4172 7290 4200 7686
rect 4344 7540 4396 7546
rect 4540 7528 4568 7704
rect 4712 7686 4764 7692
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4396 7500 4568 7528
rect 4344 7482 4396 7488
rect 4540 7410 4568 7500
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4080 7262 4200 7290
rect 3976 6996 4028 7002
rect 4080 6984 4108 7262
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 7002 4660 7482
rect 4620 6996 4672 7002
rect 4080 6956 4200 6984
rect 3976 6938 4028 6944
rect 3514 6896 3570 6905
rect 3514 6831 3570 6840
rect 3528 6798 3556 6831
rect 3516 6792 3568 6798
rect 3988 6769 4016 6938
rect 3516 6734 3568 6740
rect 3974 6760 4030 6769
rect 3974 6695 4030 6704
rect 4172 6712 4200 6956
rect 4620 6938 4672 6944
rect 4724 6934 4752 7686
rect 4816 7449 4844 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7546 5304 8452
rect 5368 7886 5396 8570
rect 5460 8498 5488 9522
rect 5552 8906 5580 9676
rect 5632 9658 5684 9664
rect 5630 9072 5686 9081
rect 5630 9007 5686 9016
rect 5644 8974 5672 9007
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5460 8362 5488 8434
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5460 8242 5488 8298
rect 5460 8214 5580 8242
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4802 7440 4858 7449
rect 5460 7410 5488 8026
rect 5552 7750 5580 8214
rect 5540 7744 5592 7750
rect 5828 7698 5856 10639
rect 5920 10266 5948 11018
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5920 10062 5948 10202
rect 6012 10198 6040 11750
rect 6184 11698 6236 11704
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6104 11150 6132 11630
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 6380 10130 6408 12406
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 6472 11354 6500 12106
rect 6564 11898 6592 12174
rect 6656 12102 6684 12854
rect 6932 12850 7052 12866
rect 6920 12844 7052 12850
rect 6972 12838 7052 12844
rect 6920 12786 6972 12792
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6932 12442 6960 12650
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6734 12336 6790 12345
rect 6734 12271 6790 12280
rect 6920 12300 6972 12306
rect 6748 12238 6776 12271
rect 6920 12242 6972 12248
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6748 11898 6776 12174
rect 6932 12073 6960 12242
rect 6918 12064 6974 12073
rect 6918 11999 6974 12008
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6472 11150 6500 11290
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6656 10538 6684 11698
rect 6748 11218 6776 11698
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6840 11014 6868 11698
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6932 10198 6960 11999
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7024 10810 7052 11086
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5920 9382 5948 9862
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 6288 9042 6316 9930
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6380 9178 6408 9522
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 7954 5948 8230
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5540 7686 5592 7692
rect 5736 7670 5856 7698
rect 4802 7375 4858 7384
rect 5264 7404 5316 7410
rect 4816 7342 4844 7375
rect 5264 7346 5316 7352
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5184 7002 5212 7278
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4816 6798 4844 6938
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4252 6724 4304 6730
rect 4172 6684 4252 6712
rect 4172 6322 4200 6684
rect 4252 6666 4304 6672
rect 4356 6458 4384 6734
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4344 6316 4396 6322
rect 4448 6304 4476 6734
rect 4396 6276 4476 6304
rect 4620 6316 4672 6322
rect 4344 6258 4396 6264
rect 4816 6304 4844 6734
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5276 6458 5304 7346
rect 5736 7290 5764 7670
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5460 7262 5764 7290
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 6458 5396 6734
rect 5460 6730 5488 7262
rect 5632 6860 5684 6866
rect 5828 6848 5856 7482
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 7002 5948 7346
rect 6012 7342 6040 8842
rect 6104 8430 6132 8978
rect 6380 8922 6408 9114
rect 6564 9042 6592 9862
rect 6932 9586 6960 10134
rect 7116 10112 7144 13330
rect 7484 13326 7512 14010
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12986 7236 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7196 12776 7248 12782
rect 7194 12744 7196 12753
rect 7248 12744 7250 12753
rect 7194 12679 7250 12688
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7208 11762 7236 12378
rect 7300 12306 7328 12786
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7300 10248 7328 11766
rect 7392 11762 7420 12582
rect 7668 12434 7696 14758
rect 7760 13462 7788 15014
rect 8680 14634 8708 16186
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8772 15638 8800 15846
rect 9324 15706 9352 16050
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 9036 15360 9088 15366
rect 8758 15328 8814 15337
rect 9036 15302 9088 15308
rect 8758 15263 8814 15272
rect 8588 14606 8708 14634
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7760 13258 7788 13398
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7484 12406 7696 12434
rect 7484 12186 7512 12406
rect 7564 12368 7616 12374
rect 7760 12322 7788 12718
rect 7616 12316 7788 12322
rect 7564 12310 7788 12316
rect 7576 12294 7788 12310
rect 7748 12232 7800 12238
rect 7484 12158 7696 12186
rect 7748 12174 7800 12180
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7484 11898 7512 12038
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 11218 7420 11562
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7300 10220 7420 10248
rect 7116 10084 7328 10112
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6736 9376 6788 9382
rect 7024 9353 7052 9454
rect 6736 9318 6788 9324
rect 7010 9344 7066 9353
rect 6552 9036 6604 9042
rect 6288 8894 6408 8922
rect 6472 8996 6552 9024
rect 6288 8566 6316 8894
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6380 8634 6408 8774
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6288 7886 6316 8502
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6000 7336 6052 7342
rect 5998 7304 6000 7313
rect 6052 7304 6054 7313
rect 5998 7239 6054 7248
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5684 6820 5856 6848
rect 5632 6802 5684 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 4672 6276 4844 6304
rect 4896 6316 4948 6322
rect 4620 6258 4672 6264
rect 4896 6258 4948 6264
rect 4908 6118 4936 6258
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 5276 5914 5304 6190
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5368 5710 5396 6394
rect 5460 6118 5488 6666
rect 5552 6458 5580 6734
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5552 6236 5580 6394
rect 5828 6322 5856 6820
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5920 6458 5948 6666
rect 6012 6458 6040 7142
rect 6196 6458 6224 7346
rect 6288 6798 6316 7686
rect 6368 7336 6420 7342
rect 6472 7324 6500 8996
rect 6552 8978 6604 8984
rect 6656 8974 6684 9318
rect 6748 8974 6776 9318
rect 7010 9279 7066 9288
rect 7116 8974 7144 9862
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6564 8498 6592 8774
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 7104 8492 7156 8498
rect 7208 8480 7236 9930
rect 7156 8452 7236 8480
rect 7104 8434 7156 8440
rect 6564 8022 6592 8434
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6420 7296 6500 7324
rect 6368 7278 6420 7284
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6288 6322 6316 6734
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 5632 6248 5684 6254
rect 5552 6208 5632 6236
rect 5632 6190 5684 6196
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5644 5778 5672 6190
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 6380 5710 6408 7278
rect 6656 7274 6684 7890
rect 6748 7886 6776 8434
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 7024 7818 7052 8298
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6550 6896 6606 6905
rect 6550 6831 6606 6840
rect 6564 6798 6592 6831
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6552 6656 6604 6662
rect 6656 6610 6684 7210
rect 6748 6934 6776 7482
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6748 6633 6776 6870
rect 6604 6604 6684 6610
rect 6552 6598 6684 6604
rect 6564 6582 6684 6598
rect 6734 6624 6790 6633
rect 6564 6322 6592 6582
rect 6734 6559 6790 6568
rect 6840 6458 6868 7142
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 7024 6322 7052 7414
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7116 5778 7144 8434
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7410 7236 8230
rect 7300 7970 7328 10084
rect 7392 9625 7420 10220
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9654 7512 9862
rect 7472 9648 7524 9654
rect 7378 9616 7434 9625
rect 7472 9590 7524 9596
rect 7378 9551 7380 9560
rect 7432 9551 7434 9560
rect 7380 9522 7432 9528
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 8974 7512 9454
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7472 8492 7524 8498
rect 7576 8480 7604 12038
rect 7668 10062 7696 12158
rect 7760 12073 7788 12174
rect 7746 12064 7802 12073
rect 7746 11999 7802 12008
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7668 9586 7696 9998
rect 7760 9654 7788 11018
rect 7852 10062 7880 14010
rect 8220 14006 8248 14418
rect 8496 14414 8524 14486
rect 8300 14408 8352 14414
rect 8484 14408 8536 14414
rect 8352 14368 8432 14396
rect 8300 14350 8352 14356
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8312 14074 8340 14214
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7944 12646 7972 13194
rect 8036 13190 8064 13874
rect 8298 13696 8354 13705
rect 8298 13631 8354 13640
rect 8312 13326 8340 13631
rect 8300 13320 8352 13326
rect 8404 13308 8432 14368
rect 8484 14350 8536 14356
rect 8496 13870 8524 14350
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8484 13320 8536 13326
rect 8404 13280 8484 13308
rect 8300 13262 8352 13268
rect 8484 13262 8536 13268
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8036 12918 8064 13126
rect 8220 12986 8248 13126
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8496 12918 8524 13262
rect 8588 13172 8616 14606
rect 8666 14512 8722 14521
rect 8666 14447 8668 14456
rect 8720 14447 8722 14456
rect 8668 14418 8720 14424
rect 8772 13938 8800 15263
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8864 13870 8892 14282
rect 9048 14074 9076 15302
rect 9140 14958 9168 15574
rect 9416 15502 9444 18906
rect 9508 18358 9536 20964
rect 9692 21576 9772 21604
rect 9692 20534 9720 21576
rect 9772 21558 9824 21564
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9784 21146 9812 21422
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9680 20528 9732 20534
rect 9732 20488 9812 20516
rect 9680 20470 9732 20476
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 9600 19961 9628 19994
rect 9586 19952 9642 19961
rect 9586 19887 9642 19896
rect 9692 19378 9720 20334
rect 9784 20262 9812 20488
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9784 19310 9812 20198
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9876 18970 9904 22066
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9496 18352 9548 18358
rect 9496 18294 9548 18300
rect 9508 17610 9536 18294
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9600 17241 9628 18770
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9692 17746 9720 18022
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9586 17232 9642 17241
rect 9586 17167 9642 17176
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9508 16658 9536 17070
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9692 16522 9720 17478
rect 9784 17338 9812 18634
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9876 18222 9904 18566
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9862 17912 9918 17921
rect 9862 17847 9918 17856
rect 9876 17678 9904 17847
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9968 17524 9996 19994
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19378 10088 19654
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10046 19136 10102 19145
rect 10046 19071 10102 19080
rect 10060 18358 10088 19071
rect 10152 18358 10180 25434
rect 10244 22778 10272 25463
rect 10336 23254 10364 26386
rect 10428 25498 10456 27406
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10520 24698 10548 29600
rect 10600 29582 10652 29588
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 10692 29232 10744 29238
rect 10692 29174 10744 29180
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 10612 28082 10640 28494
rect 10600 28076 10652 28082
rect 10600 28018 10652 28024
rect 10598 26344 10654 26353
rect 10598 26279 10654 26288
rect 10612 26246 10640 26279
rect 10704 26246 10732 29174
rect 11152 29096 11204 29102
rect 11152 29038 11204 29044
rect 11164 28762 11192 29038
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 10968 28552 11020 28558
rect 10888 28500 10968 28506
rect 11020 28500 11100 28506
rect 10888 28478 11100 28500
rect 10888 28422 10916 28478
rect 10876 28416 10928 28422
rect 10876 28358 10928 28364
rect 10968 28416 11020 28422
rect 10968 28358 11020 28364
rect 10980 28150 11008 28358
rect 10968 28144 11020 28150
rect 10782 28112 10838 28121
rect 10968 28086 11020 28092
rect 10782 28047 10784 28056
rect 10836 28047 10838 28056
rect 10784 28018 10836 28024
rect 11072 27946 11100 28478
rect 11244 28076 11296 28082
rect 11244 28018 11296 28024
rect 11060 27940 11112 27946
rect 11060 27882 11112 27888
rect 10784 27872 10836 27878
rect 10784 27814 10836 27820
rect 10796 27470 10824 27814
rect 11072 27674 11100 27882
rect 11060 27668 11112 27674
rect 11060 27610 11112 27616
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 10796 27334 10824 27406
rect 11256 27334 11284 28018
rect 11532 27946 11560 33390
rect 11992 33386 12020 34478
rect 12176 34134 12204 34546
rect 12452 34202 12480 34546
rect 12544 34513 12572 34546
rect 12530 34504 12586 34513
rect 12530 34439 12586 34448
rect 12440 34196 12492 34202
rect 12440 34138 12492 34144
rect 12164 34128 12216 34134
rect 12164 34070 12216 34076
rect 12346 34096 12402 34105
rect 12176 33833 12204 34070
rect 12346 34031 12348 34040
rect 12400 34031 12402 34040
rect 12348 34002 12400 34008
rect 12256 33992 12308 33998
rect 12256 33934 12308 33940
rect 12162 33824 12218 33833
rect 12162 33759 12218 33768
rect 12268 33658 12296 33934
rect 12256 33652 12308 33658
rect 12256 33594 12308 33600
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 11980 33380 12032 33386
rect 11980 33322 12032 33328
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 11716 31346 11744 31622
rect 11808 31482 11836 32370
rect 11888 32224 11940 32230
rect 11888 32166 11940 32172
rect 11796 31476 11848 31482
rect 11796 31418 11848 31424
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11716 30954 11744 31282
rect 11900 31278 11928 32166
rect 11992 31346 12020 33322
rect 12176 32910 12204 33458
rect 12268 33114 12296 33594
rect 12438 33552 12494 33561
rect 12438 33487 12440 33496
rect 12492 33487 12494 33496
rect 12440 33458 12492 33464
rect 12256 33108 12308 33114
rect 12256 33050 12308 33056
rect 12164 32904 12216 32910
rect 12164 32846 12216 32852
rect 12348 32360 12400 32366
rect 12348 32302 12400 32308
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 11888 31272 11940 31278
rect 12084 31249 12112 31758
rect 11888 31214 11940 31220
rect 12070 31240 12126 31249
rect 12360 31210 12388 32302
rect 12070 31175 12126 31184
rect 12348 31204 12400 31210
rect 12348 31146 12400 31152
rect 11716 30926 11928 30954
rect 11796 30252 11848 30258
rect 11796 30194 11848 30200
rect 11808 30161 11836 30194
rect 11794 30152 11850 30161
rect 11794 30087 11850 30096
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 11624 29714 11652 29990
rect 11612 29708 11664 29714
rect 11612 29650 11664 29656
rect 11796 29640 11848 29646
rect 11796 29582 11848 29588
rect 11808 29170 11836 29582
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11704 28960 11756 28966
rect 11704 28902 11756 28908
rect 11716 28422 11744 28902
rect 11808 28558 11836 29106
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11716 28150 11744 28358
rect 11704 28144 11756 28150
rect 11704 28086 11756 28092
rect 11520 27940 11572 27946
rect 11520 27882 11572 27888
rect 11612 27872 11664 27878
rect 11612 27814 11664 27820
rect 11336 27396 11388 27402
rect 11336 27338 11388 27344
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10968 27328 11020 27334
rect 10968 27270 11020 27276
rect 11244 27328 11296 27334
rect 11244 27270 11296 27276
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10600 26240 10652 26246
rect 10600 26182 10652 26188
rect 10692 26240 10744 26246
rect 10692 26182 10744 26188
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10612 24886 10640 25842
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 10600 24880 10652 24886
rect 10600 24822 10652 24828
rect 10520 24670 10640 24698
rect 10506 24576 10562 24585
rect 10506 24511 10562 24520
rect 10520 24206 10548 24511
rect 10508 24200 10560 24206
rect 10414 24168 10470 24177
rect 10508 24142 10560 24148
rect 10414 24103 10470 24112
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10336 22778 10364 22918
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10244 20942 10272 22714
rect 10428 22574 10456 24103
rect 10520 23730 10548 24142
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10506 22672 10562 22681
rect 10506 22607 10562 22616
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10324 21412 10376 21418
rect 10324 21354 10376 21360
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 10244 19514 10272 19722
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10336 19446 10364 21354
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 17649 10088 18022
rect 10244 17814 10272 18158
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10046 17640 10102 17649
rect 10046 17575 10102 17584
rect 10048 17536 10100 17542
rect 9968 17496 10048 17524
rect 10048 17478 10100 17484
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 9954 17368 10010 17377
rect 9772 17332 9824 17338
rect 10060 17338 10088 17478
rect 10152 17377 10180 17478
rect 10138 17368 10194 17377
rect 9954 17303 9956 17312
rect 9772 17274 9824 17280
rect 10008 17303 10010 17312
rect 10048 17332 10100 17338
rect 9956 17274 10008 17280
rect 10138 17303 10194 17312
rect 10048 17274 10100 17280
rect 9784 16794 9812 17274
rect 9954 17232 10010 17241
rect 9954 17167 9956 17176
rect 10008 17167 10010 17176
rect 9956 17138 10008 17144
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9508 15570 9536 16458
rect 9692 16250 9720 16458
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9508 14958 9536 15506
rect 9600 15162 9628 15982
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 9140 13938 9168 14894
rect 9324 14414 9352 14894
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9416 14618 9444 14826
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9404 14272 9456 14278
rect 9324 14232 9404 14260
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8680 13326 8708 13670
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8588 13144 8800 13172
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8024 12912 8076 12918
rect 8484 12912 8536 12918
rect 8024 12854 8076 12860
rect 8482 12880 8484 12889
rect 8536 12880 8538 12889
rect 8300 12844 8352 12850
rect 8352 12804 8432 12832
rect 8482 12815 8538 12824
rect 8300 12786 8352 12792
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7944 12374 7972 12582
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 8036 12322 8064 12378
rect 8220 12374 8248 12582
rect 8208 12368 8260 12374
rect 8036 12294 8156 12322
rect 8208 12310 8260 12316
rect 8024 12232 8076 12238
rect 8022 12200 8024 12209
rect 8076 12200 8078 12209
rect 8128 12186 8156 12294
rect 8208 12232 8260 12238
rect 8128 12180 8208 12186
rect 8128 12174 8260 12180
rect 8128 12158 8248 12174
rect 8022 12135 8078 12144
rect 8116 11824 8168 11830
rect 8168 11784 8248 11812
rect 8116 11766 8168 11772
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8128 10062 8156 10474
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7760 9382 7788 9590
rect 7852 9586 7880 9998
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7746 8664 7802 8673
rect 8036 8634 8064 9454
rect 8128 8906 8156 9862
rect 8220 9586 8248 11784
rect 8312 11762 8340 12650
rect 8404 11937 8432 12804
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8390 11928 8446 11937
rect 8390 11863 8446 11872
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8392 11756 8444 11762
rect 8496 11744 8524 12310
rect 8588 12170 8616 12922
rect 8772 12782 8800 13144
rect 8760 12776 8812 12782
rect 8680 12724 8760 12730
rect 8680 12718 8812 12724
rect 8680 12702 8800 12718
rect 8864 12714 8892 13670
rect 8956 12986 8984 13874
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8852 12708 8904 12714
rect 8680 12442 8708 12702
rect 8852 12650 8904 12656
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8680 11898 8708 12242
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8772 11762 8800 12378
rect 8444 11716 8524 11744
rect 8392 11698 8444 11704
rect 8390 11656 8446 11665
rect 8390 11591 8446 11600
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8312 10674 8340 11086
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8300 10192 8352 10198
rect 8298 10160 8300 10169
rect 8352 10160 8354 10169
rect 8298 10095 8354 10104
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8220 9450 8248 9522
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 7746 8599 7802 8608
rect 8024 8628 8076 8634
rect 7760 8566 7788 8599
rect 8024 8570 8076 8576
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7524 8452 7604 8480
rect 7656 8492 7708 8498
rect 7472 8434 7524 8440
rect 7656 8434 7708 8440
rect 7668 8090 7696 8434
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7300 7942 7420 7970
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7300 7750 7328 7822
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6390 7236 6598
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7300 5914 7328 7686
rect 7392 6118 7420 7942
rect 7760 7886 7788 8502
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7484 6798 7512 7482
rect 7944 7342 7972 7754
rect 8128 7750 8156 8842
rect 8220 8809 8248 9386
rect 8312 9178 8340 9930
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8206 8800 8262 8809
rect 8206 8735 8262 8744
rect 8404 7936 8432 11591
rect 8496 11286 8524 11716
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8588 11218 8616 11630
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 9994 8524 10950
rect 8588 10742 8616 11154
rect 8680 11082 8708 11222
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8680 10606 8708 11018
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8772 10554 8800 10678
rect 8864 10674 8892 11562
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 10674 8984 11494
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8496 8974 8524 9658
rect 8680 9568 8708 10542
rect 8772 10526 8892 10554
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8772 9722 8800 10066
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8864 9625 8892 10526
rect 8942 10160 8998 10169
rect 9048 10130 9076 13806
rect 9140 12850 9168 13874
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 11150 9168 12582
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9232 11014 9260 13398
rect 9324 11694 9352 14232
rect 9404 14214 9456 14220
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9416 13433 9444 13942
rect 9600 13938 9628 15098
rect 9784 15094 9812 16730
rect 10046 15600 10102 15609
rect 10046 15535 10102 15544
rect 10060 15502 10088 15535
rect 10152 15502 10180 16934
rect 10244 15570 10272 17750
rect 10336 17252 10364 19382
rect 10428 18193 10456 22510
rect 10520 22506 10548 22607
rect 10612 22545 10640 24670
rect 10704 24206 10732 25638
rect 10692 24200 10744 24206
rect 10692 24142 10744 24148
rect 10692 22568 10744 22574
rect 10598 22536 10654 22545
rect 10508 22500 10560 22506
rect 10692 22510 10744 22516
rect 10598 22471 10654 22480
rect 10508 22442 10560 22448
rect 10600 21888 10652 21894
rect 10598 21856 10600 21865
rect 10652 21856 10654 21865
rect 10598 21791 10654 21800
rect 10600 21140 10652 21146
rect 10600 21082 10652 21088
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10520 19292 10548 20946
rect 10612 19417 10640 21082
rect 10704 20466 10732 22510
rect 10796 21146 10824 25842
rect 10888 25226 10916 27066
rect 10980 26858 11008 27270
rect 11348 26994 11376 27338
rect 11336 26988 11388 26994
rect 11336 26930 11388 26936
rect 10968 26852 11020 26858
rect 10968 26794 11020 26800
rect 11152 26852 11204 26858
rect 11152 26794 11204 26800
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10980 25974 11008 26182
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 11058 25936 11114 25945
rect 11058 25871 11060 25880
rect 11112 25871 11114 25880
rect 11060 25842 11112 25848
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 10980 25498 11008 25638
rect 11164 25537 11192 26794
rect 11348 26586 11376 26930
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11520 26580 11572 26586
rect 11520 26522 11572 26528
rect 11336 26376 11388 26382
rect 11388 26336 11468 26364
rect 11336 26318 11388 26324
rect 11244 26240 11296 26246
rect 11244 26182 11296 26188
rect 11336 26240 11388 26246
rect 11336 26182 11388 26188
rect 11256 26042 11284 26182
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 11348 25974 11376 26182
rect 11336 25968 11388 25974
rect 11336 25910 11388 25916
rect 11150 25528 11206 25537
rect 10968 25492 11020 25498
rect 11150 25463 11206 25472
rect 10968 25434 11020 25440
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10876 25220 10928 25226
rect 10876 25162 10928 25168
rect 10874 24984 10930 24993
rect 10874 24919 10930 24928
rect 10888 24682 10916 24919
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 10980 24410 11008 25230
rect 11058 25120 11114 25129
rect 11058 25055 11114 25064
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10796 19446 10824 20810
rect 10888 20233 10916 24210
rect 11072 23662 11100 25055
rect 11164 24818 11192 25366
rect 11336 25220 11388 25226
rect 11336 25162 11388 25168
rect 11348 24818 11376 25162
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11336 24608 11388 24614
rect 11440 24596 11468 26336
rect 11532 25974 11560 26522
rect 11520 25968 11572 25974
rect 11520 25910 11572 25916
rect 11624 25514 11652 27814
rect 11808 27470 11836 28358
rect 11796 27464 11848 27470
rect 11796 27406 11848 27412
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 11388 24568 11468 24596
rect 11532 25486 11652 25514
rect 11336 24550 11388 24556
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10968 23248 11020 23254
rect 10968 23190 11020 23196
rect 10980 22710 11008 23190
rect 11164 23186 11192 24550
rect 11348 24256 11376 24550
rect 11532 24274 11560 25486
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11624 24954 11652 25230
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 11716 24698 11744 27270
rect 11796 26240 11848 26246
rect 11796 26182 11848 26188
rect 11808 24818 11836 26182
rect 11900 25362 11928 30926
rect 12360 30734 12388 31146
rect 11980 30728 12032 30734
rect 11980 30670 12032 30676
rect 12348 30728 12400 30734
rect 12348 30670 12400 30676
rect 11992 26450 12020 30670
rect 12636 29730 12664 34598
rect 12716 33992 12768 33998
rect 12716 33934 12768 33940
rect 12728 33697 12756 33934
rect 12714 33688 12770 33697
rect 12714 33623 12770 33632
rect 12728 33590 12756 33623
rect 12716 33584 12768 33590
rect 12716 33526 12768 33532
rect 12544 29702 12664 29730
rect 12256 29640 12308 29646
rect 12256 29582 12308 29588
rect 12268 29170 12296 29582
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 12440 29028 12492 29034
rect 12440 28970 12492 28976
rect 12348 28552 12400 28558
rect 12452 28529 12480 28970
rect 12348 28494 12400 28500
rect 12438 28520 12494 28529
rect 12164 28484 12216 28490
rect 12164 28426 12216 28432
rect 12176 27470 12204 28426
rect 12360 28082 12388 28494
rect 12438 28455 12494 28464
rect 12256 28076 12308 28082
rect 12256 28018 12308 28024
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12164 27464 12216 27470
rect 12164 27406 12216 27412
rect 12176 26994 12204 27406
rect 12268 27402 12296 28018
rect 12360 27538 12388 28018
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12440 27464 12492 27470
rect 12440 27406 12492 27412
rect 12256 27396 12308 27402
rect 12256 27338 12308 27344
rect 12452 27305 12480 27406
rect 12544 27402 12572 29702
rect 12624 29640 12676 29646
rect 12820 29628 12848 34682
rect 13004 33998 13032 35634
rect 13096 35562 13124 36128
rect 13176 36110 13228 36116
rect 13188 35630 13216 36110
rect 13372 35766 13400 36178
rect 13360 35760 13412 35766
rect 13360 35702 13412 35708
rect 13556 35698 13584 36178
rect 14108 36174 14136 36654
rect 14280 36644 14332 36650
rect 14280 36586 14332 36592
rect 14188 36576 14240 36582
rect 14188 36518 14240 36524
rect 14200 36242 14228 36518
rect 14188 36236 14240 36242
rect 14188 36178 14240 36184
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 13544 35692 13596 35698
rect 13544 35634 13596 35640
rect 14004 35692 14056 35698
rect 14004 35634 14056 35640
rect 13176 35624 13228 35630
rect 13176 35566 13228 35572
rect 13268 35624 13320 35630
rect 13268 35566 13320 35572
rect 13084 35556 13136 35562
rect 13084 35498 13136 35504
rect 13096 35034 13124 35498
rect 13176 35488 13228 35494
rect 13176 35430 13228 35436
rect 13188 35154 13216 35430
rect 13176 35148 13228 35154
rect 13176 35090 13228 35096
rect 13096 35006 13216 35034
rect 13084 34400 13136 34406
rect 13084 34342 13136 34348
rect 13096 34066 13124 34342
rect 13084 34060 13136 34066
rect 13084 34002 13136 34008
rect 12992 33992 13044 33998
rect 12992 33934 13044 33940
rect 13004 33454 13032 33934
rect 12992 33448 13044 33454
rect 12992 33390 13044 33396
rect 13188 33368 13216 35006
rect 13280 34610 13308 35566
rect 13268 34604 13320 34610
rect 13268 34546 13320 34552
rect 13556 34542 13584 35634
rect 13636 35488 13688 35494
rect 13636 35430 13688 35436
rect 13912 35488 13964 35494
rect 13912 35430 13964 35436
rect 13648 35222 13676 35430
rect 13636 35216 13688 35222
rect 13636 35158 13688 35164
rect 13924 35086 13952 35430
rect 14016 35154 14044 35634
rect 14200 35222 14228 36178
rect 14292 36174 14320 36586
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 14752 36106 14780 36654
rect 14844 36174 14872 36722
rect 14832 36168 14884 36174
rect 14832 36110 14884 36116
rect 14740 36100 14792 36106
rect 14740 36042 14792 36048
rect 14752 35714 14780 36042
rect 14752 35698 14872 35714
rect 14936 35698 14964 36722
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 15212 35698 15240 35974
rect 15304 35834 15332 36722
rect 15842 36136 15898 36145
rect 15842 36071 15898 36080
rect 15292 35828 15344 35834
rect 15292 35770 15344 35776
rect 15476 35828 15528 35834
rect 15476 35770 15528 35776
rect 14372 35692 14424 35698
rect 14752 35692 14884 35698
rect 14752 35686 14832 35692
rect 14372 35634 14424 35640
rect 14832 35634 14884 35640
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 15108 35692 15160 35698
rect 15108 35634 15160 35640
rect 15200 35692 15252 35698
rect 15200 35634 15252 35640
rect 14280 35488 14332 35494
rect 14280 35430 14332 35436
rect 14188 35216 14240 35222
rect 14188 35158 14240 35164
rect 14004 35148 14056 35154
rect 14004 35090 14056 35096
rect 13912 35080 13964 35086
rect 13912 35022 13964 35028
rect 14016 34950 14044 35090
rect 14096 35012 14148 35018
rect 14096 34954 14148 34960
rect 14004 34944 14056 34950
rect 14004 34886 14056 34892
rect 13912 34740 13964 34746
rect 13912 34682 13964 34688
rect 13636 34604 13688 34610
rect 13636 34546 13688 34552
rect 13544 34536 13596 34542
rect 13544 34478 13596 34484
rect 13648 34406 13676 34546
rect 13818 34504 13874 34513
rect 13818 34439 13874 34448
rect 13636 34400 13688 34406
rect 13636 34342 13688 34348
rect 13360 33516 13412 33522
rect 13360 33458 13412 33464
rect 13268 33380 13320 33386
rect 13188 33340 13268 33368
rect 13268 33322 13320 33328
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 12676 29600 12848 29628
rect 12624 29582 12676 29588
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12438 27296 12494 27305
rect 12360 27254 12438 27282
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 11980 26444 12032 26450
rect 11980 26386 12032 26392
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 12070 25936 12126 25945
rect 12070 25871 12126 25880
rect 11980 25832 12032 25838
rect 11980 25774 12032 25780
rect 11992 25430 12020 25774
rect 11980 25424 12032 25430
rect 11980 25366 12032 25372
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 11716 24670 11836 24698
rect 11256 24228 11376 24256
rect 11520 24268 11572 24274
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 11060 23112 11112 23118
rect 11058 23080 11060 23089
rect 11112 23080 11114 23089
rect 11058 23015 11114 23024
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 22030 11008 22510
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 11072 21486 11100 22918
rect 11164 21894 11192 23122
rect 11256 22930 11284 24228
rect 11520 24210 11572 24216
rect 11336 24132 11388 24138
rect 11336 24074 11388 24080
rect 11348 23633 11376 24074
rect 11334 23624 11390 23633
rect 11334 23559 11390 23568
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11348 23118 11376 23462
rect 11532 23118 11560 24210
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11520 23112 11572 23118
rect 11520 23054 11572 23060
rect 11610 23080 11666 23089
rect 11610 23015 11612 23024
rect 11664 23015 11666 23024
rect 11612 22986 11664 22992
rect 11256 22902 11468 22930
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11348 22030 11376 22714
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11164 21690 11192 21830
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11244 21616 11296 21622
rect 11164 21564 11244 21570
rect 11164 21558 11296 21564
rect 11164 21542 11284 21558
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11072 21078 11100 21422
rect 11060 21072 11112 21078
rect 11060 21014 11112 21020
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 10874 20224 10930 20233
rect 10874 20159 10930 20168
rect 11072 20058 11100 20878
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 10784 19440 10836 19446
rect 10598 19408 10654 19417
rect 10784 19382 10836 19388
rect 10598 19343 10654 19352
rect 10692 19304 10744 19310
rect 10520 19264 10640 19292
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 10520 18426 10548 18634
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10414 18184 10470 18193
rect 10414 18119 10470 18128
rect 10612 17977 10640 19264
rect 10692 19246 10744 19252
rect 10704 18970 10732 19246
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10704 18290 10732 18770
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10598 17968 10654 17977
rect 10598 17903 10654 17912
rect 10704 17814 10732 18022
rect 10692 17808 10744 17814
rect 10796 17785 10824 19382
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10888 18630 10916 19246
rect 11164 18834 11192 21542
rect 11348 21434 11376 21626
rect 11256 21406 11376 21434
rect 11256 21350 11284 21406
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11348 21146 11376 21286
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11440 20534 11468 22902
rect 11716 22778 11744 23462
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11610 22536 11666 22545
rect 11610 22471 11666 22480
rect 11624 22438 11652 22471
rect 11520 22432 11572 22438
rect 11520 22374 11572 22380
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11532 22030 11560 22374
rect 11716 22216 11744 22578
rect 11808 22409 11836 24670
rect 11900 23798 11928 25298
rect 11992 24342 12020 25366
rect 12084 24818 12112 25871
rect 12176 25226 12204 26250
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 12176 25129 12204 25162
rect 12162 25120 12218 25129
rect 12162 25055 12218 25064
rect 12360 24993 12388 27254
rect 12438 27231 12494 27240
rect 12544 27062 12572 27338
rect 12532 27056 12584 27062
rect 12532 26998 12584 27004
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12544 25838 12572 26318
rect 12636 26042 12664 29582
rect 12714 29336 12770 29345
rect 12714 29271 12770 29280
rect 12728 29170 12756 29271
rect 12912 29170 12940 32506
rect 12992 31748 13044 31754
rect 12992 31690 13044 31696
rect 12716 29164 12768 29170
rect 12716 29106 12768 29112
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 12808 29096 12860 29102
rect 12808 29038 12860 29044
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 12728 27538 12756 28562
rect 12820 27849 12848 29038
rect 12900 28620 12952 28626
rect 13004 28608 13032 31690
rect 13280 31142 13308 33322
rect 13372 33289 13400 33458
rect 13358 33280 13414 33289
rect 13358 33215 13414 33224
rect 13648 31906 13676 34342
rect 13832 34202 13860 34439
rect 13820 34196 13872 34202
rect 13820 34138 13872 34144
rect 13728 33992 13780 33998
rect 13728 33934 13780 33940
rect 13740 33833 13768 33934
rect 13924 33862 13952 34682
rect 14004 34468 14056 34474
rect 14004 34410 14056 34416
rect 14016 34066 14044 34410
rect 14108 34202 14136 34954
rect 14188 34944 14240 34950
rect 14188 34886 14240 34892
rect 14096 34196 14148 34202
rect 14096 34138 14148 34144
rect 14200 34082 14228 34886
rect 14292 34678 14320 35430
rect 14384 35290 14412 35634
rect 14648 35556 14700 35562
rect 14648 35498 14700 35504
rect 14372 35284 14424 35290
rect 14372 35226 14424 35232
rect 14556 35148 14608 35154
rect 14556 35090 14608 35096
rect 14280 34672 14332 34678
rect 14280 34614 14332 34620
rect 14372 34536 14424 34542
rect 14372 34478 14424 34484
rect 14004 34060 14056 34066
rect 14004 34002 14056 34008
rect 14108 34054 14228 34082
rect 14280 34128 14332 34134
rect 14280 34070 14332 34076
rect 13820 33856 13872 33862
rect 13726 33824 13782 33833
rect 13820 33798 13872 33804
rect 13912 33856 13964 33862
rect 13912 33798 13964 33804
rect 13726 33759 13782 33768
rect 13832 33522 13860 33798
rect 13820 33516 13872 33522
rect 13820 33458 13872 33464
rect 14004 33516 14056 33522
rect 14108 33504 14136 34054
rect 14292 33980 14320 34070
rect 14384 33998 14412 34478
rect 14568 34134 14596 35090
rect 14660 34950 14688 35498
rect 14648 34944 14700 34950
rect 14648 34886 14700 34892
rect 14740 34944 14792 34950
rect 14740 34886 14792 34892
rect 14752 34678 14780 34886
rect 14740 34672 14792 34678
rect 14740 34614 14792 34620
rect 14648 34400 14700 34406
rect 14648 34342 14700 34348
rect 14660 34134 14688 34342
rect 14556 34128 14608 34134
rect 14556 34070 14608 34076
rect 14648 34128 14700 34134
rect 14648 34070 14700 34076
rect 14740 34128 14792 34134
rect 14740 34070 14792 34076
rect 14200 33952 14320 33980
rect 14372 33992 14424 33998
rect 14200 33561 14228 33952
rect 14372 33934 14424 33940
rect 14462 33824 14518 33833
rect 14462 33759 14518 33768
rect 14278 33688 14334 33697
rect 14278 33623 14334 33632
rect 14056 33476 14136 33504
rect 14186 33552 14242 33561
rect 14186 33487 14188 33496
rect 14004 33458 14056 33464
rect 14240 33487 14242 33496
rect 14188 33458 14240 33464
rect 13728 33448 13780 33454
rect 13912 33448 13964 33454
rect 13728 33390 13780 33396
rect 13910 33416 13912 33425
rect 13964 33416 13966 33425
rect 13740 33300 13768 33390
rect 13910 33351 13966 33360
rect 13912 33312 13964 33318
rect 13740 33272 13912 33300
rect 13912 33254 13964 33260
rect 13912 32496 13964 32502
rect 13912 32438 13964 32444
rect 13924 32366 13952 32438
rect 13912 32360 13964 32366
rect 13912 32302 13964 32308
rect 13726 32056 13782 32065
rect 13726 31991 13728 32000
rect 13780 31991 13782 32000
rect 13728 31962 13780 31968
rect 13648 31878 13768 31906
rect 13452 31816 13504 31822
rect 13372 31776 13452 31804
rect 13268 31136 13320 31142
rect 13268 31078 13320 31084
rect 13176 30592 13228 30598
rect 13176 30534 13228 30540
rect 13268 30592 13320 30598
rect 13268 30534 13320 30540
rect 13082 30288 13138 30297
rect 13082 30223 13138 30232
rect 13096 29782 13124 30223
rect 13188 30190 13216 30534
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13280 30054 13308 30534
rect 13268 30048 13320 30054
rect 13268 29990 13320 29996
rect 13372 29782 13400 31776
rect 13452 31758 13504 31764
rect 13542 31104 13598 31113
rect 13542 31039 13598 31048
rect 13556 29832 13584 31039
rect 13464 29804 13584 29832
rect 13084 29776 13136 29782
rect 13084 29718 13136 29724
rect 13360 29776 13412 29782
rect 13360 29718 13412 29724
rect 13372 29617 13400 29718
rect 13358 29608 13414 29617
rect 13358 29543 13414 29552
rect 13176 29504 13228 29510
rect 13176 29446 13228 29452
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13360 29504 13412 29510
rect 13360 29446 13412 29452
rect 13082 29336 13138 29345
rect 13082 29271 13138 29280
rect 12952 28580 13032 28608
rect 12900 28562 12952 28568
rect 12912 27878 12940 28562
rect 13096 28558 13124 29271
rect 13188 29102 13216 29446
rect 13280 29170 13308 29446
rect 13268 29164 13320 29170
rect 13268 29106 13320 29112
rect 13176 29096 13228 29102
rect 13176 29038 13228 29044
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 13096 28150 13124 28494
rect 13188 28490 13216 29038
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 13188 28218 13216 28426
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13084 28144 13136 28150
rect 13084 28086 13136 28092
rect 12900 27872 12952 27878
rect 12806 27840 12862 27849
rect 12900 27814 12952 27820
rect 12806 27775 12862 27784
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 12900 27464 12952 27470
rect 13096 27452 13124 28086
rect 12952 27424 13124 27452
rect 12900 27406 12952 27412
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12728 26353 12756 26998
rect 12912 26994 12940 27406
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 12900 26988 12952 26994
rect 12900 26930 12952 26936
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12808 26376 12860 26382
rect 12714 26344 12770 26353
rect 12808 26318 12860 26324
rect 12714 26279 12770 26288
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12624 25900 12676 25906
rect 12728 25888 12756 26182
rect 12820 25945 12848 26318
rect 12912 26314 12940 26522
rect 13004 26314 13032 27066
rect 12900 26308 12952 26314
rect 12900 26250 12952 26256
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 12676 25860 12756 25888
rect 12806 25936 12862 25945
rect 12806 25871 12808 25880
rect 12624 25842 12676 25848
rect 12860 25871 12862 25880
rect 12808 25842 12860 25848
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 12346 24984 12402 24993
rect 12346 24919 12402 24928
rect 12254 24848 12310 24857
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 12176 24792 12254 24800
rect 12176 24772 12256 24792
rect 11980 24336 12032 24342
rect 11980 24278 12032 24284
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11992 23798 12020 24142
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11978 23352 12034 23361
rect 11978 23287 11980 23296
rect 12032 23287 12034 23296
rect 11980 23258 12032 23264
rect 11992 23118 12020 23258
rect 11980 23112 12032 23118
rect 11886 23080 11942 23089
rect 11980 23054 12032 23060
rect 12176 23066 12204 24772
rect 12308 24783 12310 24792
rect 12256 24754 12308 24760
rect 12452 24682 12480 25638
rect 12544 24954 12572 25774
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 12532 24948 12584 24954
rect 12584 24908 12664 24936
rect 12532 24890 12584 24896
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12440 24676 12492 24682
rect 12440 24618 12492 24624
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12268 23866 12296 24006
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12360 23662 12388 24550
rect 12544 24449 12572 24754
rect 12530 24440 12586 24449
rect 12636 24410 12664 24908
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12714 24712 12770 24721
rect 12714 24647 12770 24656
rect 12530 24375 12586 24384
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12268 23254 12296 23462
rect 12256 23248 12308 23254
rect 12636 23225 12664 24074
rect 12256 23190 12308 23196
rect 12622 23216 12678 23225
rect 12622 23151 12678 23160
rect 12348 23112 12400 23118
rect 12346 23080 12348 23089
rect 12624 23112 12676 23118
rect 12400 23080 12402 23089
rect 12176 23038 12296 23066
rect 11886 23015 11888 23024
rect 11940 23015 11942 23024
rect 11888 22986 11940 22992
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11794 22400 11850 22409
rect 11794 22335 11850 22344
rect 11796 22228 11848 22234
rect 11716 22188 11796 22216
rect 11796 22170 11848 22176
rect 11808 22030 11836 22170
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11532 21078 11560 21286
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11428 20528 11480 20534
rect 11428 20470 11480 20476
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 17977 10916 18566
rect 10968 18284 11020 18290
rect 11072 18272 11100 18702
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11020 18244 11100 18272
rect 10968 18226 11020 18232
rect 11152 18216 11204 18222
rect 11072 18176 11152 18204
rect 10874 17968 10930 17977
rect 10874 17903 10930 17912
rect 11072 17785 11100 18176
rect 11152 18158 11204 18164
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 10692 17750 10744 17756
rect 10782 17776 10838 17785
rect 10416 17740 10468 17746
rect 10782 17711 10838 17720
rect 11058 17776 11114 17785
rect 11058 17711 11114 17720
rect 10416 17682 10468 17688
rect 10428 17377 10456 17682
rect 10692 17672 10744 17678
rect 10744 17632 10824 17660
rect 10692 17614 10744 17620
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10414 17368 10470 17377
rect 10414 17303 10470 17312
rect 10416 17264 10468 17270
rect 10336 17224 10416 17252
rect 10416 17206 10468 17212
rect 10520 17202 10548 17478
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10324 17060 10376 17066
rect 10324 17002 10376 17008
rect 10336 16794 10364 17002
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10612 16522 10640 17274
rect 10704 17270 10732 17478
rect 10796 17377 10824 17632
rect 11164 17610 11192 18022
rect 11256 17882 11284 18634
rect 11428 18352 11480 18358
rect 11348 18300 11428 18306
rect 11348 18294 11480 18300
rect 11348 18278 11468 18294
rect 11348 18086 11376 18278
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11348 17954 11376 18022
rect 11348 17926 11560 17954
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11334 17776 11390 17785
rect 11334 17711 11390 17720
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11348 17524 11376 17711
rect 11440 17678 11468 17818
rect 11532 17678 11560 17926
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11256 17496 11376 17524
rect 11428 17536 11480 17542
rect 11426 17504 11428 17513
rect 11480 17504 11482 17513
rect 10782 17368 10838 17377
rect 10782 17303 10838 17312
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10966 17232 11022 17241
rect 10966 17167 11022 17176
rect 10782 16960 10838 16969
rect 10782 16895 10838 16904
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10612 15706 10640 15982
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9402 13424 9458 13433
rect 9402 13359 9458 13368
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12238 9444 13262
rect 9508 12374 9536 13670
rect 9692 12986 9720 14894
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9784 14482 9812 14554
rect 9954 14512 10010 14521
rect 9772 14476 9824 14482
rect 9954 14447 9956 14456
rect 9772 14418 9824 14424
rect 10008 14447 10010 14456
rect 9956 14418 10008 14424
rect 10060 14278 10088 15438
rect 10152 15162 10180 15438
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10152 14550 10180 15098
rect 10244 14958 10272 15302
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10520 14618 10548 15438
rect 10796 15366 10824 16895
rect 10980 16114 11008 17167
rect 11256 17134 11284 17496
rect 11426 17439 11482 17448
rect 11624 17377 11652 21966
rect 11900 21570 11928 22646
rect 11992 22574 12020 22918
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 12084 22420 12112 22918
rect 12176 22778 12204 22918
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12162 22672 12218 22681
rect 12162 22607 12164 22616
rect 12216 22607 12218 22616
rect 12164 22578 12216 22584
rect 11992 22392 12112 22420
rect 11992 22030 12020 22392
rect 12070 22264 12126 22273
rect 12070 22199 12126 22208
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11900 21554 12020 21570
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11796 21548 11848 21554
rect 11900 21548 12032 21554
rect 11900 21542 11980 21548
rect 11796 21490 11848 21496
rect 11980 21490 12032 21496
rect 11716 21418 11744 21490
rect 11704 21412 11756 21418
rect 11704 21354 11756 21360
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 11610 17368 11666 17377
rect 11336 17332 11388 17338
rect 11716 17338 11744 20878
rect 11808 20058 11836 21490
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11808 19378 11836 19994
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11900 18766 11928 19178
rect 11796 18760 11848 18766
rect 11794 18728 11796 18737
rect 11888 18760 11940 18766
rect 11848 18728 11850 18737
rect 11888 18702 11940 18708
rect 11794 18663 11850 18672
rect 11900 18426 11928 18702
rect 11888 18420 11940 18426
rect 11808 18380 11888 18408
rect 11808 17610 11836 18380
rect 11888 18362 11940 18368
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11900 17678 11928 18226
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11610 17303 11666 17312
rect 11704 17332 11756 17338
rect 11336 17274 11388 17280
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11072 16590 11100 17070
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11348 16250 11376 17274
rect 11624 16946 11652 17303
rect 11704 17274 11756 17280
rect 11532 16918 11652 16946
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10690 15192 10746 15201
rect 10690 15127 10746 15136
rect 10704 15026 10732 15127
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10520 14482 10548 14554
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9876 13530 9904 13806
rect 10428 13734 10456 14214
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9416 11898 9444 12174
rect 9508 11898 9536 12310
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9600 11762 9628 12854
rect 9692 12714 9720 12922
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9324 11150 9352 11630
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 8942 10095 8998 10104
rect 9036 10124 9088 10130
rect 8956 10062 8984 10095
rect 9036 10066 9088 10072
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8850 9616 8906 9625
rect 8680 9540 8800 9568
rect 8850 9551 8852 9560
rect 8576 9376 8628 9382
rect 8772 9353 8800 9540
rect 8904 9551 8906 9560
rect 8852 9522 8904 9528
rect 8576 9318 8628 9324
rect 8758 9344 8814 9353
rect 8588 9042 8616 9318
rect 8758 9279 8814 9288
rect 8772 9110 8800 9279
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8956 8974 8984 9862
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9048 9217 9076 9522
rect 9140 9382 9168 10610
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9324 9722 9352 9930
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9034 9208 9090 9217
rect 9034 9143 9090 9152
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8496 8566 8524 8910
rect 8680 8634 8708 8910
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8680 7954 8708 8570
rect 8772 7954 8800 8774
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8668 7948 8720 7954
rect 8404 7908 8524 7936
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8404 7478 8432 7754
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7944 6798 7972 7278
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 6934 8248 7142
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8404 6866 8432 7414
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7656 6792 7708 6798
rect 7932 6792 7984 6798
rect 7656 6734 7708 6740
rect 7746 6760 7802 6769
rect 7472 6656 7524 6662
rect 7470 6624 7472 6633
rect 7524 6624 7526 6633
rect 7470 6559 7526 6568
rect 7668 6458 7696 6734
rect 7932 6734 7984 6740
rect 7746 6695 7802 6704
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7760 6390 7788 6695
rect 8496 6662 8524 7908
rect 8668 7890 8720 7896
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8680 7818 8708 7890
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8758 7576 8814 7585
rect 8758 7511 8814 7520
rect 8772 7478 8800 7511
rect 8864 7478 8892 8230
rect 8956 7546 8984 8366
rect 9048 8090 9076 8366
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8760 7472 8812 7478
rect 8666 7440 8722 7449
rect 8760 7414 8812 7420
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8666 7375 8668 7384
rect 8720 7375 8722 7384
rect 8668 7346 8720 7352
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8588 7002 8616 7210
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8574 6896 8630 6905
rect 8574 6831 8630 6840
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 7760 5302 7788 6326
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8128 5370 8156 5782
rect 8588 5710 8616 6831
rect 8772 6458 8800 7414
rect 9036 7404 9088 7410
rect 9140 7392 9168 9318
rect 9232 8634 9260 9522
rect 9416 9450 9444 10610
rect 9508 10470 9536 10610
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9088 7364 9168 7392
rect 9036 7346 9088 7352
rect 9048 7313 9076 7346
rect 9232 7324 9260 8570
rect 9324 8498 9352 8774
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9508 7954 9536 8910
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9416 7478 9444 7890
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9034 7304 9090 7313
rect 9034 7239 9090 7248
rect 9140 7296 9260 7324
rect 8852 6792 8904 6798
rect 9140 6780 9168 7296
rect 9218 6896 9274 6905
rect 9508 6866 9536 7890
rect 9600 7410 9628 9454
rect 9678 8528 9734 8537
rect 9678 8463 9680 8472
rect 9732 8463 9734 8472
rect 9680 8434 9732 8440
rect 9784 7478 9812 13466
rect 10230 13424 10286 13433
rect 10230 13359 10286 13368
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9968 12646 9996 13126
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 10060 12442 10088 12786
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10060 12306 10088 12378
rect 10152 12374 10180 13262
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 10060 11898 10088 12106
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9968 11150 9996 11834
rect 10152 11200 10180 12174
rect 10060 11172 10180 11200
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 9586 9904 10406
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 10060 8838 10088 11172
rect 10244 11098 10272 13359
rect 10324 13252 10376 13258
rect 10324 13194 10376 13200
rect 10336 12986 10364 13194
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10336 11898 10364 12718
rect 10428 12714 10456 13670
rect 10704 13462 10732 14554
rect 10796 14074 10824 15302
rect 10888 15026 10916 15370
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10152 11070 10272 11098
rect 10152 9160 10180 11070
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10606 10272 10950
rect 10428 10742 10456 12650
rect 10520 12084 10548 12854
rect 10612 12782 10640 13262
rect 10704 12850 10732 13398
rect 10888 12889 10916 14826
rect 10980 13938 11008 16050
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15570 11284 15846
rect 11348 15570 11376 16186
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10874 12880 10930 12889
rect 10692 12844 10744 12850
rect 10874 12815 10930 12824
rect 10692 12786 10744 12792
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10612 12238 10640 12718
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10520 12056 10640 12084
rect 10612 11762 10640 12056
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10598 11656 10654 11665
rect 10520 11558 10548 11630
rect 10598 11591 10654 11600
rect 10612 11558 10640 11591
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10520 11082 10548 11494
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10612 10962 10640 11086
rect 10520 10934 10640 10962
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10336 9382 10364 10610
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10232 9172 10284 9178
rect 10152 9132 10232 9160
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10060 8090 10088 8570
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10152 7970 10180 9132
rect 10232 9114 10284 9120
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8480 10272 8774
rect 10428 8634 10456 9522
rect 10520 9466 10548 10934
rect 10704 10674 10732 11834
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 9512 10652 9518
rect 10520 9460 10600 9466
rect 10520 9454 10652 9460
rect 10520 9438 10640 9454
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9042 10548 9318
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10612 8498 10640 9438
rect 10324 8492 10376 8498
rect 10244 8452 10324 8480
rect 10244 8362 10272 8452
rect 10324 8434 10376 8440
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10060 7942 10180 7970
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9784 7290 9812 7414
rect 10060 7410 10088 7942
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9692 7262 9812 7290
rect 9218 6831 9274 6840
rect 9496 6860 9548 6866
rect 9232 6798 9260 6831
rect 9496 6802 9548 6808
rect 8904 6752 9168 6780
rect 9220 6792 9272 6798
rect 8852 6734 8904 6740
rect 9220 6734 9272 6740
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8680 5574 8708 6190
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8036 2446 8064 4558
rect 8128 3466 8156 5306
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 3602 8340 3878
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8404 3534 8432 5510
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8312 2514 8340 2994
rect 8496 2990 8524 3538
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8680 2922 8708 4014
rect 8864 3738 8892 4014
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 3194 8800 3334
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9048 3126 9076 6598
rect 9508 6322 9536 6802
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9692 6202 9720 7262
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9784 6390 9812 7142
rect 9968 7002 9996 7142
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6458 9996 6598
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9600 6186 9720 6202
rect 9588 6180 9720 6186
rect 9640 6174 9720 6180
rect 9588 6122 9640 6128
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5710 9444 6054
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5302 9352 5510
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9600 4078 9628 5714
rect 9692 4214 9720 6174
rect 9784 4282 9812 6326
rect 9968 5846 9996 6394
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 10060 5642 10088 6054
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10152 5234 10180 7822
rect 10244 7206 10272 7822
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7478 10364 7686
rect 10520 7546 10548 7822
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10336 6866 10364 7142
rect 10428 7002 10456 7346
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10244 6474 10272 6666
rect 10428 6662 10456 6802
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10704 6474 10732 9998
rect 10796 8378 10824 12582
rect 10888 12374 10916 12815
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11354 10916 12174
rect 10980 11914 11008 13874
rect 11072 12102 11100 14758
rect 11242 14512 11298 14521
rect 11242 14447 11298 14456
rect 11256 14414 11284 14447
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10980 11886 11100 11914
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10888 11132 10916 11290
rect 10968 11144 11020 11150
rect 10888 11104 10968 11132
rect 10968 11086 11020 11092
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9722 10916 9998
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10888 8498 10916 9386
rect 10980 9178 11008 9522
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10980 8566 11008 9114
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11072 8401 11100 11886
rect 11256 11762 11284 14350
rect 11532 14074 11560 16918
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11624 16590 11652 16730
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16114 11744 16526
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 13258 11560 13670
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11440 12434 11468 12922
rect 11440 12406 11560 12434
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11164 11354 11192 11698
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11058 8392 11114 8401
rect 10796 8350 11008 8378
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 8090 10824 8230
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10796 7818 10824 8026
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10244 6446 10732 6474
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10244 5166 10272 6446
rect 10796 5914 10824 7278
rect 10888 6254 10916 7482
rect 10980 7342 11008 8350
rect 11058 8327 11114 8336
rect 11164 7818 11192 8842
rect 11348 8634 11376 12038
rect 11532 11694 11560 12406
rect 11716 12306 11744 16050
rect 11992 12434 12020 21490
rect 12084 21146 12112 22199
rect 12268 21978 12296 23038
rect 12624 23054 12676 23060
rect 12346 23015 12402 23024
rect 12532 23044 12584 23050
rect 12532 22986 12584 22992
rect 12544 22506 12572 22986
rect 12636 22710 12664 23054
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12348 22500 12400 22506
rect 12348 22442 12400 22448
rect 12532 22500 12584 22506
rect 12532 22442 12584 22448
rect 12360 22234 12388 22442
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 12176 21962 12296 21978
rect 12164 21956 12296 21962
rect 12216 21950 12296 21956
rect 12346 21992 12402 22001
rect 12346 21927 12348 21936
rect 12164 21898 12216 21904
rect 12400 21927 12402 21936
rect 12348 21898 12400 21904
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12254 21176 12310 21185
rect 12072 21140 12124 21146
rect 12254 21111 12256 21120
rect 12072 21082 12124 21088
rect 12308 21111 12310 21120
rect 12256 21082 12308 21088
rect 12084 20602 12112 21082
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 12084 19718 12112 20334
rect 12268 19922 12296 20946
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 12084 19145 12112 19654
rect 12360 19174 12388 21422
rect 12544 21350 12572 22442
rect 12728 21842 12756 24647
rect 12820 23866 12848 24754
rect 12912 24721 12940 24754
rect 12898 24712 12954 24721
rect 12898 24647 12954 24656
rect 13004 24206 13032 25638
rect 13084 25220 13136 25226
rect 13084 25162 13136 25168
rect 13096 24818 13124 25162
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13176 24744 13228 24750
rect 13176 24686 13228 24692
rect 13188 24342 13216 24686
rect 13280 24682 13308 28494
rect 13372 27130 13400 29446
rect 13464 29209 13492 29804
rect 13740 29730 13768 31878
rect 13924 31482 13952 32302
rect 14016 31958 14044 33458
rect 14096 33380 14148 33386
rect 14096 33322 14148 33328
rect 14108 33289 14136 33322
rect 14094 33280 14150 33289
rect 14094 33215 14150 33224
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 14004 31952 14056 31958
rect 14004 31894 14056 31900
rect 13912 31476 13964 31482
rect 13912 31418 13964 31424
rect 13912 31272 13964 31278
rect 13912 31214 13964 31220
rect 13924 30122 13952 31214
rect 14016 30122 14044 31894
rect 14108 31890 14136 32846
rect 14200 32774 14228 33458
rect 14292 33454 14320 33623
rect 14476 33522 14504 33759
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14464 33516 14516 33522
rect 14464 33458 14516 33464
rect 14280 33448 14332 33454
rect 14280 33390 14332 33396
rect 14384 32842 14412 33458
rect 14568 33130 14596 34070
rect 14648 33856 14700 33862
rect 14648 33798 14700 33804
rect 14660 33318 14688 33798
rect 14752 33522 14780 34070
rect 14740 33516 14792 33522
rect 14740 33458 14792 33464
rect 14648 33312 14700 33318
rect 14648 33254 14700 33260
rect 14476 33102 14596 33130
rect 14372 32836 14424 32842
rect 14372 32778 14424 32784
rect 14188 32768 14240 32774
rect 14188 32710 14240 32716
rect 14096 31884 14148 31890
rect 14096 31826 14148 31832
rect 14096 30660 14148 30666
rect 14096 30602 14148 30608
rect 14108 30394 14136 30602
rect 14096 30388 14148 30394
rect 14096 30330 14148 30336
rect 14094 30152 14150 30161
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 14004 30116 14056 30122
rect 14094 30087 14150 30096
rect 14004 30058 14056 30064
rect 14108 29832 14136 30087
rect 13556 29702 13768 29730
rect 14016 29804 14136 29832
rect 13450 29200 13506 29209
rect 13450 29135 13506 29144
rect 13464 29102 13492 29135
rect 13452 29096 13504 29102
rect 13452 29038 13504 29044
rect 13556 28558 13584 29702
rect 13636 29640 13688 29646
rect 13820 29640 13872 29646
rect 13636 29582 13688 29588
rect 13726 29608 13782 29617
rect 13648 29510 13676 29582
rect 13820 29582 13872 29588
rect 13726 29543 13782 29552
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13648 29345 13676 29446
rect 13634 29336 13690 29345
rect 13634 29271 13690 29280
rect 13648 29170 13676 29271
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13740 29050 13768 29543
rect 13832 29102 13860 29582
rect 14016 29578 14044 29804
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 14004 29572 14056 29578
rect 14004 29514 14056 29520
rect 14016 29209 14044 29514
rect 14002 29200 14058 29209
rect 14002 29135 14058 29144
rect 13648 29022 13768 29050
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13452 28008 13504 28014
rect 13452 27950 13504 27956
rect 13464 27470 13492 27950
rect 13556 27470 13584 28018
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13544 27464 13596 27470
rect 13544 27406 13596 27412
rect 13360 27124 13412 27130
rect 13360 27066 13412 27072
rect 13464 26994 13492 27406
rect 13452 26988 13504 26994
rect 13452 26930 13504 26936
rect 13360 26784 13412 26790
rect 13360 26726 13412 26732
rect 13372 26450 13400 26726
rect 13648 26602 13676 29022
rect 13832 28994 13860 29038
rect 13740 28966 13860 28994
rect 13740 28558 13768 28966
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13740 28014 13768 28494
rect 13912 28416 13964 28422
rect 13912 28358 13964 28364
rect 13728 28008 13780 28014
rect 13728 27950 13780 27956
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13556 26574 13676 26602
rect 13360 26444 13412 26450
rect 13360 26386 13412 26392
rect 13452 26240 13504 26246
rect 13452 26182 13504 26188
rect 13464 25226 13492 26182
rect 13452 25220 13504 25226
rect 13452 25162 13504 25168
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 13268 24676 13320 24682
rect 13268 24618 13320 24624
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13176 24336 13228 24342
rect 13082 24304 13138 24313
rect 13176 24278 13228 24284
rect 13082 24239 13138 24248
rect 13096 24206 13124 24239
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12820 23050 12848 23666
rect 13096 23610 13124 24142
rect 13188 23730 13216 24278
rect 13280 24206 13308 24346
rect 13268 24200 13320 24206
rect 13372 24188 13400 24822
rect 13320 24160 13400 24188
rect 13268 24142 13320 24148
rect 13372 23730 13400 24160
rect 13556 23730 13584 26574
rect 13636 26512 13688 26518
rect 13636 26454 13688 26460
rect 13648 23730 13676 26454
rect 13740 26382 13768 26726
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13820 26308 13872 26314
rect 13820 26250 13872 26256
rect 13832 26042 13860 26250
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13832 25226 13860 25978
rect 13820 25220 13872 25226
rect 13820 25162 13872 25168
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 13740 24410 13768 25094
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13004 23582 13124 23610
rect 12808 23044 12860 23050
rect 12808 22986 12860 22992
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 12820 22166 12848 22646
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12636 21814 12756 21842
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12636 21162 12664 21814
rect 12716 21684 12768 21690
rect 12820 21672 12848 22102
rect 12912 22030 12940 22918
rect 13004 22094 13032 23582
rect 13084 23520 13136 23526
rect 13280 23497 13308 23666
rect 13556 23526 13584 23666
rect 13740 23633 13768 24074
rect 13726 23624 13782 23633
rect 13726 23559 13782 23568
rect 13544 23520 13596 23526
rect 13084 23462 13136 23468
rect 13266 23488 13322 23497
rect 13096 22438 13124 23462
rect 13544 23462 13596 23468
rect 13266 23423 13322 23432
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 13188 22710 13216 23258
rect 13634 23216 13690 23225
rect 13452 23180 13504 23186
rect 13372 23140 13452 23168
rect 13372 22710 13400 23140
rect 13634 23151 13690 23160
rect 13452 23122 13504 23128
rect 13176 22704 13228 22710
rect 13176 22646 13228 22652
rect 13360 22704 13412 22710
rect 13360 22646 13412 22652
rect 13450 22672 13506 22681
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 13004 22066 13124 22094
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12768 21644 12848 21672
rect 12716 21626 12768 21632
rect 13096 21622 13124 22066
rect 13372 22030 13400 22646
rect 13450 22607 13452 22616
rect 13504 22607 13506 22616
rect 13544 22636 13596 22642
rect 13452 22578 13504 22584
rect 13544 22578 13596 22584
rect 13464 22030 13492 22578
rect 13556 22234 13584 22578
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 13268 21956 13320 21962
rect 13268 21898 13320 21904
rect 13280 21690 13308 21898
rect 13648 21706 13676 23151
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13740 22574 13768 22918
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13832 22234 13860 22986
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 13832 21894 13860 22170
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13268 21684 13320 21690
rect 13648 21678 13768 21706
rect 13268 21626 13320 21632
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 12544 21134 12664 21162
rect 12990 21176 13046 21185
rect 12544 20874 12572 21134
rect 12990 21111 13046 21120
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12636 20942 12664 21014
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12544 20058 12572 20334
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12544 19530 12572 19858
rect 12452 19514 12572 19530
rect 12440 19508 12572 19514
rect 12492 19502 12572 19508
rect 12440 19450 12492 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12348 19168 12400 19174
rect 12070 19136 12126 19145
rect 12348 19110 12400 19116
rect 12070 19071 12126 19080
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12084 18766 12112 18906
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12084 18290 12112 18702
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12176 17882 12204 18226
rect 12268 18222 12296 18634
rect 12360 18630 12388 19110
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12452 17882 12480 18838
rect 12636 18170 12664 19314
rect 12728 19174 12756 20878
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12820 19310 12848 20810
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12728 18290 12756 18838
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12820 18426 12848 18702
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12532 18148 12584 18154
rect 12636 18142 12756 18170
rect 12532 18090 12584 18096
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12254 17776 12310 17785
rect 12254 17711 12310 17720
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 17338 12204 17614
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 16114 12112 16390
rect 12268 16182 12296 17711
rect 12452 17678 12480 17818
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12544 17270 12572 18090
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12636 17338 12664 17614
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12544 16726 12572 17206
rect 12728 16726 12756 18142
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16794 12848 17138
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12532 16720 12584 16726
rect 12716 16720 12768 16726
rect 12532 16662 12584 16668
rect 12622 16688 12678 16697
rect 12716 16662 12768 16668
rect 12622 16623 12678 16632
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11900 12406 12020 12434
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11532 10062 11560 11630
rect 11624 10130 11652 12174
rect 11716 11286 11744 12242
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11900 10198 11928 12406
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11992 11150 12020 11766
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11992 9654 12020 10678
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12084 10266 12112 10474
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11624 8974 11652 9386
rect 11716 9178 11744 9522
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10980 6866 11008 7278
rect 11072 7002 11100 7278
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10980 6186 11008 6802
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9876 4554 9904 5034
rect 10796 5030 10824 5510
rect 10888 5114 10916 5578
rect 11072 5302 11100 6734
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10888 5086 11100 5114
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 8220 2106 8248 2246
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 8404 800 8432 2790
rect 8680 2774 8708 2858
rect 8956 2854 8984 2994
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8588 2746 8708 2774
rect 8588 2446 8616 2746
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9140 2378 9168 3674
rect 9232 3534 9260 4014
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9232 2990 9260 3470
rect 9324 2990 9352 3470
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9232 2378 9260 2790
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9784 1714 9812 3606
rect 9876 3466 9904 4490
rect 9968 4146 9996 4626
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10152 3942 10180 4490
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10796 3602 10824 4218
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 3602 10916 3878
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9876 3058 9904 3402
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9876 2394 9904 2994
rect 10796 2650 10824 3538
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10232 2440 10284 2446
rect 9876 2388 10232 2394
rect 9876 2382 10284 2388
rect 9876 2378 10272 2382
rect 9864 2372 10272 2378
rect 9916 2366 10272 2372
rect 9864 2314 9916 2320
rect 9692 1686 9812 1714
rect 9692 800 9720 1686
rect 10336 800 10364 2586
rect 10980 800 11008 4490
rect 11072 4146 11100 5086
rect 11164 4690 11192 6598
rect 11256 5302 11284 6666
rect 11348 5642 11376 8570
rect 11624 8498 11652 8910
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8498 12020 8774
rect 12176 8634 12204 15302
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 10062 12296 12174
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11624 8294 11652 8434
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11440 7954 11468 8230
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11440 5386 11468 7346
rect 11518 6896 11574 6905
rect 11518 6831 11520 6840
rect 11572 6831 11574 6840
rect 11520 6802 11572 6808
rect 11624 6633 11652 7346
rect 11716 7206 11744 8434
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11796 7336 11848 7342
rect 11794 7304 11796 7313
rect 11848 7304 11850 7313
rect 11794 7239 11850 7248
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11900 6730 11928 8230
rect 12254 7440 12310 7449
rect 12254 7375 12256 7384
rect 12308 7375 12310 7384
rect 12256 7346 12308 7352
rect 12360 7290 12388 14418
rect 12452 13802 12480 16050
rect 12636 15502 12664 16623
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12544 14890 12572 15438
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12728 13938 12756 16526
rect 12806 16144 12862 16153
rect 12806 16079 12808 16088
rect 12860 16079 12862 16088
rect 12808 16050 12860 16056
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12820 15638 12848 15914
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12452 11354 12480 11630
rect 12544 11354 12572 13466
rect 12728 13326 12756 13738
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12820 13190 12848 15438
rect 12912 14482 12940 20198
rect 13004 19174 13032 21111
rect 13280 20942 13308 21354
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 13096 20602 13124 20810
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13188 19378 13216 20742
rect 13280 20262 13308 20878
rect 13372 20874 13400 21014
rect 13360 20868 13412 20874
rect 13360 20810 13412 20816
rect 13372 20602 13400 20810
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13280 19378 13308 20198
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13084 18760 13136 18766
rect 12990 18728 13046 18737
rect 13084 18702 13136 18708
rect 12990 18663 13046 18672
rect 13004 18290 13032 18663
rect 13096 18426 13124 18702
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13188 18306 13216 18634
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13096 18278 13216 18306
rect 13096 18154 13124 18278
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 17134 13032 17614
rect 13188 17610 13216 18158
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13082 17368 13138 17377
rect 13280 17354 13308 19110
rect 13082 17303 13138 17312
rect 13188 17326 13308 17354
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12912 13326 12940 13942
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 13004 12322 13032 16186
rect 13096 14226 13124 17303
rect 13188 14482 13216 17326
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13280 14618 13308 15982
rect 13372 15366 13400 20538
rect 13464 19242 13492 21014
rect 13556 19446 13584 21286
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13648 19446 13676 19994
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18766 13492 19178
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13544 18284 13596 18290
rect 13464 18244 13544 18272
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13268 14408 13320 14414
rect 13464 14362 13492 18244
rect 13648 18272 13676 18906
rect 13596 18244 13676 18272
rect 13544 18226 13596 18232
rect 13740 17898 13768 21678
rect 13924 19446 13952 28358
rect 14108 27470 14136 29650
rect 14200 29170 14228 32710
rect 14372 31748 14424 31754
rect 14372 31690 14424 31696
rect 14384 31482 14412 31690
rect 14372 31476 14424 31482
rect 14372 31418 14424 31424
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14292 30938 14320 31078
rect 14280 30932 14332 30938
rect 14280 30874 14332 30880
rect 14280 30320 14332 30326
rect 14280 30262 14332 30268
rect 14292 30190 14320 30262
rect 14280 30184 14332 30190
rect 14280 30126 14332 30132
rect 14372 29640 14424 29646
rect 14476 29628 14504 33102
rect 14648 32428 14700 32434
rect 14648 32370 14700 32376
rect 14660 30666 14688 32370
rect 14844 31754 14872 35634
rect 14936 35222 14964 35634
rect 15120 35290 15148 35634
rect 15384 35624 15436 35630
rect 15488 35612 15516 35770
rect 15436 35584 15516 35612
rect 15384 35566 15436 35572
rect 15382 35320 15438 35329
rect 15108 35284 15160 35290
rect 15382 35255 15438 35264
rect 15108 35226 15160 35232
rect 14924 35216 14976 35222
rect 14924 35158 14976 35164
rect 14936 34542 14964 35158
rect 15396 35086 15424 35255
rect 15016 35080 15068 35086
rect 15016 35022 15068 35028
rect 15384 35080 15436 35086
rect 15384 35022 15436 35028
rect 14924 34536 14976 34542
rect 14924 34478 14976 34484
rect 15028 34474 15056 35022
rect 15292 34944 15344 34950
rect 15292 34886 15344 34892
rect 15304 34746 15332 34886
rect 15292 34740 15344 34746
rect 15292 34682 15344 34688
rect 15200 34604 15252 34610
rect 15200 34546 15252 34552
rect 15016 34468 15068 34474
rect 15016 34410 15068 34416
rect 14922 34096 14978 34105
rect 14922 34031 14924 34040
rect 14976 34031 14978 34040
rect 14924 34002 14976 34008
rect 14924 33924 14976 33930
rect 14924 33866 14976 33872
rect 14936 33658 14964 33866
rect 15028 33674 15056 34410
rect 15212 33998 15240 34546
rect 15200 33992 15252 33998
rect 15292 33992 15344 33998
rect 15200 33934 15252 33940
rect 15290 33960 15292 33969
rect 15344 33960 15346 33969
rect 15396 33946 15424 35022
rect 15212 33833 15240 33934
rect 15346 33918 15424 33946
rect 15290 33895 15346 33904
rect 15198 33824 15254 33833
rect 15198 33759 15254 33768
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 15028 33646 15332 33674
rect 15396 33658 15424 33918
rect 14924 32836 14976 32842
rect 14924 32778 14976 32784
rect 14936 32366 14964 32778
rect 14924 32360 14976 32366
rect 14924 32302 14976 32308
rect 14924 31884 14976 31890
rect 14924 31826 14976 31832
rect 14752 31726 14872 31754
rect 14648 30660 14700 30666
rect 14648 30602 14700 30608
rect 14660 30394 14688 30602
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 14424 29600 14504 29628
rect 14372 29582 14424 29588
rect 14384 29238 14412 29582
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 14464 29164 14516 29170
rect 14464 29106 14516 29112
rect 14372 29096 14424 29102
rect 14372 29038 14424 29044
rect 14280 29028 14332 29034
rect 14280 28970 14332 28976
rect 14188 28484 14240 28490
rect 14188 28426 14240 28432
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14200 27112 14228 28426
rect 14292 27606 14320 28970
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 14200 27084 14320 27112
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14096 26308 14148 26314
rect 14096 26250 14148 26256
rect 14108 25702 14136 26250
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14002 23488 14058 23497
rect 14002 23423 14058 23432
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13832 18426 13860 19178
rect 13820 18420 13872 18426
rect 14016 18408 14044 23423
rect 14108 21418 14136 24006
rect 14200 22094 14228 26930
rect 14292 26353 14320 27084
rect 14384 26926 14412 29038
rect 14476 28082 14504 29106
rect 14464 28076 14516 28082
rect 14516 28036 14596 28064
rect 14464 28018 14516 28024
rect 14372 26920 14424 26926
rect 14372 26862 14424 26868
rect 14278 26344 14334 26353
rect 14278 26279 14334 26288
rect 14280 25220 14332 25226
rect 14280 25162 14332 25168
rect 14292 24818 14320 25162
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14292 24188 14320 24754
rect 14384 24290 14412 26862
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 14476 25294 14504 25842
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14476 24410 14504 25230
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14384 24262 14504 24290
rect 14292 24160 14412 24188
rect 14280 23248 14332 23254
rect 14280 23190 14332 23196
rect 14292 22642 14320 23190
rect 14384 23118 14412 24160
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14370 22944 14426 22953
rect 14370 22879 14426 22888
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 14200 22066 14320 22094
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14292 20942 14320 22066
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14108 20398 14136 20742
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14200 19514 14228 20878
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14292 20058 14320 20470
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14384 19802 14412 22879
rect 14476 21350 14504 24262
rect 14568 23254 14596 28036
rect 14752 27130 14780 31726
rect 14936 31346 14964 31826
rect 14924 31340 14976 31346
rect 14924 31282 14976 31288
rect 15028 30870 15056 33646
rect 15198 33552 15254 33561
rect 15198 33487 15200 33496
rect 15252 33487 15254 33496
rect 15200 33458 15252 33464
rect 15108 31816 15160 31822
rect 15106 31784 15108 31793
rect 15160 31784 15162 31793
rect 15106 31719 15162 31728
rect 15016 30864 15068 30870
rect 15016 30806 15068 30812
rect 14832 30728 14884 30734
rect 14832 30670 14884 30676
rect 14844 30258 14872 30670
rect 15212 30598 15240 33458
rect 15304 33454 15332 33646
rect 15384 33652 15436 33658
rect 15384 33594 15436 33600
rect 15292 33448 15344 33454
rect 15292 33390 15344 33396
rect 15488 33402 15516 35584
rect 15856 34610 15884 36071
rect 16132 35698 16160 36858
rect 16592 36854 16620 37130
rect 16580 36848 16632 36854
rect 16580 36790 16632 36796
rect 16488 36780 16540 36786
rect 16488 36722 16540 36728
rect 16500 36666 16528 36722
rect 16500 36638 16712 36666
rect 16684 36378 16712 36638
rect 16672 36372 16724 36378
rect 16672 36314 16724 36320
rect 16488 36100 16540 36106
rect 16488 36042 16540 36048
rect 16500 35834 16528 36042
rect 16488 35828 16540 35834
rect 16488 35770 16540 35776
rect 16120 35692 16172 35698
rect 16120 35634 16172 35640
rect 16672 35692 16724 35698
rect 16672 35634 16724 35640
rect 16304 35624 16356 35630
rect 16580 35624 16632 35630
rect 16304 35566 16356 35572
rect 16500 35584 16580 35612
rect 16316 35290 16344 35566
rect 16500 35494 16528 35584
rect 16580 35566 16632 35572
rect 16488 35488 16540 35494
rect 16488 35430 16540 35436
rect 16580 35488 16632 35494
rect 16580 35430 16632 35436
rect 16304 35284 16356 35290
rect 16304 35226 16356 35232
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 16488 35080 16540 35086
rect 16488 35022 16540 35028
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 16224 34649 16252 34682
rect 16210 34640 16266 34649
rect 15844 34604 15896 34610
rect 16210 34575 16266 34584
rect 15844 34546 15896 34552
rect 15568 34536 15620 34542
rect 15568 34478 15620 34484
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 15752 34536 15804 34542
rect 15752 34478 15804 34484
rect 15580 33590 15608 34478
rect 15672 34202 15700 34478
rect 15660 34196 15712 34202
rect 15660 34138 15712 34144
rect 15764 33862 15792 34478
rect 16316 34474 16344 35022
rect 16396 34944 16448 34950
rect 16396 34886 16448 34892
rect 16408 34474 16436 34886
rect 16500 34542 16528 35022
rect 16488 34536 16540 34542
rect 16488 34478 16540 34484
rect 16212 34468 16264 34474
rect 16212 34410 16264 34416
rect 16304 34468 16356 34474
rect 16304 34410 16356 34416
rect 16396 34468 16448 34474
rect 16396 34410 16448 34416
rect 16224 34354 16252 34410
rect 16224 34326 16344 34354
rect 16120 34196 16172 34202
rect 16120 34138 16172 34144
rect 15844 33924 15896 33930
rect 15844 33866 15896 33872
rect 15752 33856 15804 33862
rect 15752 33798 15804 33804
rect 15856 33590 15884 33866
rect 16028 33856 16080 33862
rect 16028 33798 16080 33804
rect 15568 33584 15620 33590
rect 15568 33526 15620 33532
rect 15844 33584 15896 33590
rect 15844 33526 15896 33532
rect 15566 33416 15622 33425
rect 15488 33374 15566 33402
rect 15566 33351 15568 33360
rect 15620 33351 15622 33360
rect 15568 33322 15620 33328
rect 15844 33040 15896 33046
rect 15844 32982 15896 32988
rect 15856 32434 15884 32982
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15476 32224 15528 32230
rect 15476 32166 15528 32172
rect 15488 31958 15516 32166
rect 15476 31952 15528 31958
rect 15476 31894 15528 31900
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15384 31340 15436 31346
rect 15384 31282 15436 31288
rect 15396 31249 15424 31282
rect 15382 31240 15438 31249
rect 15382 31175 15438 31184
rect 15292 30864 15344 30870
rect 15292 30806 15344 30812
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 15108 30252 15160 30258
rect 15108 30194 15160 30200
rect 14922 29064 14978 29073
rect 14922 28999 14924 29008
rect 14976 28999 14978 29008
rect 14924 28970 14976 28976
rect 14832 28960 14884 28966
rect 14832 28902 14884 28908
rect 14844 28082 14872 28902
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 15028 28558 15056 28698
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 14832 28076 14884 28082
rect 14884 28036 14964 28064
rect 14832 28018 14884 28024
rect 14740 27124 14792 27130
rect 14740 27066 14792 27072
rect 14740 26852 14792 26858
rect 14740 26794 14792 26800
rect 14752 26217 14780 26794
rect 14830 26344 14886 26353
rect 14830 26279 14886 26288
rect 14738 26208 14794 26217
rect 14738 26143 14794 26152
rect 14752 24206 14780 26143
rect 14844 25906 14872 26279
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14844 24750 14872 25094
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 14844 24206 14872 24686
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 14556 23248 14608 23254
rect 14556 23190 14608 23196
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14568 22012 14596 23054
rect 14660 22778 14688 24074
rect 14752 23594 14780 24142
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14740 23588 14792 23594
rect 14740 23530 14792 23536
rect 14738 23216 14794 23225
rect 14738 23151 14740 23160
rect 14792 23151 14794 23160
rect 14740 23122 14792 23128
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14752 22710 14780 23122
rect 14844 22953 14872 23802
rect 14830 22944 14886 22953
rect 14830 22879 14886 22888
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14660 22545 14688 22578
rect 14832 22568 14884 22574
rect 14646 22536 14702 22545
rect 14832 22510 14884 22516
rect 14646 22471 14702 22480
rect 14844 22166 14872 22510
rect 14832 22160 14884 22166
rect 14832 22102 14884 22108
rect 14740 22024 14792 22030
rect 14568 21984 14740 22012
rect 14740 21966 14792 21972
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14556 20256 14608 20262
rect 14660 20233 14688 21490
rect 14556 20198 14608 20204
rect 14646 20224 14702 20233
rect 14292 19774 14412 19802
rect 14568 19786 14596 20198
rect 14646 20159 14702 20168
rect 14556 19780 14608 19786
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14108 18970 14136 19314
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14200 18698 14228 19450
rect 14292 19446 14320 19774
rect 14556 19722 14608 19728
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14554 19680 14610 19689
rect 14384 19514 14412 19654
rect 14554 19615 14610 19624
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14568 19378 14596 19615
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14016 18380 14136 18408
rect 13820 18362 13872 18368
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13648 17870 13768 17898
rect 14016 17882 14044 18226
rect 14004 17876 14056 17882
rect 13542 17368 13598 17377
rect 13542 17303 13598 17312
rect 13556 17270 13584 17303
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13556 16114 13584 16458
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13648 15910 13676 17870
rect 14004 17818 14056 17824
rect 13726 17096 13782 17105
rect 13726 17031 13782 17040
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13320 14356 13492 14362
rect 13268 14350 13492 14356
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13280 14334 13492 14350
rect 13096 14198 13308 14226
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13096 12442 13124 13806
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13004 12294 13124 12322
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12544 11014 12572 11154
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12728 10810 12756 11086
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12544 9674 12572 10066
rect 12820 9994 12848 11630
rect 12912 11558 12940 12038
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 13004 11370 13032 12174
rect 12912 11354 13032 11370
rect 12900 11348 13032 11354
rect 12952 11342 13032 11348
rect 12900 11290 12952 11296
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12728 9722 12756 9930
rect 12716 9716 12768 9722
rect 12544 9646 12664 9674
rect 12716 9658 12768 9664
rect 12912 9654 12940 11290
rect 12530 9480 12586 9489
rect 12530 9415 12532 9424
rect 12584 9415 12586 9424
rect 12532 9386 12584 9392
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 9042 12480 9318
rect 12544 9110 12572 9386
rect 12636 9364 12664 9646
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12716 9376 12768 9382
rect 12636 9336 12716 9364
rect 12716 9318 12768 9324
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8634 12664 8774
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12728 7954 12756 9318
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 8362 12848 8774
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 7948 12768 7954
rect 12636 7908 12716 7936
rect 12636 7478 12664 7908
rect 12716 7890 12768 7896
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12728 7342 12756 7482
rect 12912 7478 12940 7686
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12176 7262 12388 7290
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11610 6624 11666 6633
rect 11610 6559 11666 6568
rect 11518 6488 11574 6497
rect 12084 6474 12112 7142
rect 12176 6798 12204 7262
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 11518 6423 11520 6432
rect 11572 6423 11574 6432
rect 11808 6446 12112 6474
rect 11520 6394 11572 6400
rect 11532 6118 11560 6394
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11624 5642 11652 6258
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11440 5358 11652 5386
rect 11716 5370 11744 6258
rect 11808 5778 11836 6446
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11796 5772 11848 5778
rect 11848 5732 11928 5760
rect 11796 5714 11848 5720
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11256 4826 11284 5102
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11348 4758 11376 5170
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 11256 4078 11284 4626
rect 11244 4072 11296 4078
rect 11150 4040 11206 4049
rect 11244 4014 11296 4020
rect 11150 3975 11206 3984
rect 11164 2446 11192 3975
rect 11440 3602 11468 5170
rect 11624 4826 11652 5358
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11716 4622 11744 5306
rect 11808 5030 11836 5306
rect 11900 5302 11928 5732
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11900 5166 11928 5238
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4758 11928 4966
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 12084 4622 12112 6326
rect 12176 4690 12204 6734
rect 12268 6202 12296 7142
rect 12636 7002 12664 7278
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12452 6322 12480 6666
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12716 6248 12768 6254
rect 12268 6186 12388 6202
rect 12716 6190 12768 6196
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12268 6180 12400 6186
rect 12268 6174 12348 6180
rect 12348 6122 12400 6128
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5914 12480 6054
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12728 5778 12756 6190
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12912 5681 12940 6190
rect 12898 5672 12954 5681
rect 12532 5636 12584 5642
rect 12584 5596 12848 5624
rect 12898 5607 12954 5616
rect 12532 5578 12584 5584
rect 12820 5302 12848 5596
rect 12808 5296 12860 5302
rect 12728 5256 12808 5284
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 12072 4616 12124 4622
rect 12360 4570 12388 4626
rect 12072 4558 12124 4564
rect 11716 4146 11744 4558
rect 11808 4486 11836 4558
rect 12268 4542 12388 4570
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11716 3738 11744 4082
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11256 3058 11284 3538
rect 11808 3482 11836 3674
rect 11624 3454 11836 3482
rect 11624 3398 11652 3454
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11256 2514 11284 2994
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11888 2508 11940 2514
rect 11992 2496 12020 4422
rect 12164 4208 12216 4214
rect 12268 4196 12296 4542
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12216 4168 12296 4196
rect 12164 4150 12216 4156
rect 12268 2854 12296 4168
rect 12360 3126 12388 4422
rect 12728 4214 12756 5256
rect 12808 5238 12860 5244
rect 13004 5030 13032 6734
rect 13096 5302 13124 12294
rect 13188 11762 13216 13126
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13280 9194 13308 14198
rect 13372 11694 13400 14334
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13464 11150 13492 11698
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13464 11014 13492 11086
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13188 9166 13308 9194
rect 13188 8566 13216 9166
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13188 8362 13216 8502
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13188 7886 13216 8298
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13188 6458 13216 6734
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13280 6322 13308 8026
rect 13372 7886 13400 9658
rect 13464 9586 13492 9998
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13556 9450 13584 14350
rect 13740 14346 13768 17031
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16182 13860 16934
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13924 14074 13952 14350
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14016 13326 14044 13874
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13648 12170 13676 13262
rect 14108 12434 14136 18380
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 14200 16114 14228 16458
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14200 12918 14228 15846
rect 14292 15570 14320 19246
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14292 12986 14320 13194
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14384 12866 14412 15914
rect 14476 15910 14504 17614
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14476 13326 14504 15846
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14384 12838 14504 12866
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 13924 12406 14136 12434
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13648 11626 13676 12106
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13740 9058 13768 11154
rect 13924 10282 13952 12406
rect 14384 12374 14412 12718
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11830 14228 12038
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13832 10254 13952 10282
rect 13832 9160 13860 10254
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13924 9586 13952 10066
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 14016 9518 14044 11086
rect 14292 10044 14320 12106
rect 14384 11150 14412 12310
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14476 10713 14504 12838
rect 14568 12102 14596 18634
rect 14660 17882 14688 20159
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14660 15570 14688 17818
rect 14752 17814 14780 21966
rect 14844 21962 14872 22102
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14936 21622 14964 28036
rect 15120 26042 15148 30194
rect 15304 29714 15332 30806
rect 15488 29850 15516 31758
rect 15660 31272 15712 31278
rect 15566 31240 15622 31249
rect 15660 31214 15712 31220
rect 15566 31175 15622 31184
rect 15580 30433 15608 31175
rect 15672 30666 15700 31214
rect 15752 31204 15804 31210
rect 15752 31146 15804 31152
rect 15764 30734 15792 31146
rect 15752 30728 15804 30734
rect 15752 30670 15804 30676
rect 15660 30660 15712 30666
rect 15660 30602 15712 30608
rect 15566 30424 15622 30433
rect 15566 30359 15622 30368
rect 15476 29844 15528 29850
rect 15476 29786 15528 29792
rect 15292 29708 15344 29714
rect 15292 29650 15344 29656
rect 15304 29238 15332 29650
rect 15292 29232 15344 29238
rect 15292 29174 15344 29180
rect 15488 29102 15516 29786
rect 15568 29572 15620 29578
rect 15568 29514 15620 29520
rect 15580 29102 15608 29514
rect 15672 29102 15700 30602
rect 15752 29640 15804 29646
rect 15856 29628 15884 32370
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15948 32026 15976 32166
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 15948 31929 15976 31962
rect 15934 31920 15990 31929
rect 15934 31855 15990 31864
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 15948 30870 15976 31622
rect 15936 30864 15988 30870
rect 15936 30806 15988 30812
rect 16040 29782 16068 33798
rect 16132 33522 16160 34138
rect 16316 33930 16344 34326
rect 16304 33924 16356 33930
rect 16304 33866 16356 33872
rect 16316 33590 16344 33866
rect 16408 33658 16436 34410
rect 16488 34400 16540 34406
rect 16486 34368 16488 34377
rect 16540 34368 16542 34377
rect 16486 34303 16542 34312
rect 16396 33652 16448 33658
rect 16396 33594 16448 33600
rect 16304 33584 16356 33590
rect 16304 33526 16356 33532
rect 16120 33516 16172 33522
rect 16120 33458 16172 33464
rect 16500 33436 16528 34303
rect 16316 33408 16528 33436
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 16132 32298 16160 32914
rect 16212 32428 16264 32434
rect 16212 32370 16264 32376
rect 16120 32292 16172 32298
rect 16120 32234 16172 32240
rect 16132 30734 16160 32234
rect 16224 31278 16252 32370
rect 16212 31272 16264 31278
rect 16212 31214 16264 31220
rect 16210 30832 16266 30841
rect 16210 30767 16212 30776
rect 16264 30767 16266 30776
rect 16212 30738 16264 30744
rect 16120 30728 16172 30734
rect 16120 30670 16172 30676
rect 16212 30660 16264 30666
rect 16212 30602 16264 30608
rect 16224 30569 16252 30602
rect 16210 30560 16266 30569
rect 16210 30495 16266 30504
rect 16028 29776 16080 29782
rect 16028 29718 16080 29724
rect 15804 29600 16068 29628
rect 15752 29582 15804 29588
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15292 29096 15344 29102
rect 15476 29096 15528 29102
rect 15292 29038 15344 29044
rect 15382 29064 15438 29073
rect 15304 28762 15332 29038
rect 15476 29038 15528 29044
rect 15568 29096 15620 29102
rect 15568 29038 15620 29044
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 15382 28999 15384 29008
rect 15436 28999 15438 29008
rect 15384 28970 15436 28976
rect 15764 28762 15792 29106
rect 15856 29102 15884 29446
rect 16040 29306 16068 29600
rect 16224 29578 16252 30495
rect 16212 29572 16264 29578
rect 16212 29514 16264 29520
rect 16120 29504 16172 29510
rect 16120 29446 16172 29452
rect 16028 29300 16080 29306
rect 16028 29242 16080 29248
rect 15844 29096 15896 29102
rect 15844 29038 15896 29044
rect 15292 28756 15344 28762
rect 15292 28698 15344 28704
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 15200 28688 15252 28694
rect 15200 28630 15252 28636
rect 15212 27674 15240 28630
rect 15200 27668 15252 27674
rect 15200 27610 15252 27616
rect 15200 26512 15252 26518
rect 15200 26454 15252 26460
rect 15108 26036 15160 26042
rect 15108 25978 15160 25984
rect 15212 25906 15240 26454
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15028 25362 15056 25842
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 15016 25356 15068 25362
rect 15016 25298 15068 25304
rect 15120 25294 15148 25774
rect 15108 25288 15160 25294
rect 15108 25230 15160 25236
rect 15106 24848 15162 24857
rect 15106 24783 15162 24792
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 15028 23866 15056 24074
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15028 22506 15056 23054
rect 15016 22500 15068 22506
rect 15016 22442 15068 22448
rect 14924 21616 14976 21622
rect 14924 21558 14976 21564
rect 15028 21468 15056 22442
rect 14936 21457 15056 21468
rect 14936 21448 15070 21457
rect 14936 21440 15014 21448
rect 14936 19334 14964 21440
rect 15014 21383 15070 21392
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 15028 20398 15056 20538
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15028 19922 15056 20334
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 15120 19718 15148 24783
rect 15212 24682 15240 25842
rect 15304 25294 15332 28698
rect 16040 28558 16068 29242
rect 15384 28552 15436 28558
rect 15568 28552 15620 28558
rect 15384 28494 15436 28500
rect 15566 28520 15568 28529
rect 15660 28552 15712 28558
rect 15620 28520 15622 28529
rect 15396 28218 15424 28494
rect 15660 28494 15712 28500
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 15566 28455 15622 28464
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15474 28248 15530 28257
rect 15384 28212 15436 28218
rect 15474 28183 15530 28192
rect 15384 28154 15436 28160
rect 15396 27538 15424 28154
rect 15488 28082 15516 28183
rect 15476 28076 15528 28082
rect 15476 28018 15528 28024
rect 15384 27532 15436 27538
rect 15384 27474 15436 27480
rect 15488 27402 15516 28018
rect 15580 27402 15608 28358
rect 15672 28014 15700 28494
rect 15660 28008 15712 28014
rect 15660 27950 15712 27956
rect 15476 27396 15528 27402
rect 15476 27338 15528 27344
rect 15568 27396 15620 27402
rect 15568 27338 15620 27344
rect 15672 27282 15700 27950
rect 15580 27254 15700 27282
rect 15292 25288 15344 25294
rect 15344 25248 15424 25276
rect 15292 25230 15344 25236
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15290 23352 15346 23361
rect 15290 23287 15346 23296
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 15212 21486 15240 22986
rect 15304 22778 15332 23287
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15304 22216 15332 22510
rect 15396 22409 15424 25248
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15488 23633 15516 23666
rect 15474 23624 15530 23633
rect 15474 23559 15530 23568
rect 15580 23508 15608 27254
rect 16028 26920 16080 26926
rect 16028 26862 16080 26868
rect 16040 26382 16068 26862
rect 15844 26376 15896 26382
rect 16028 26376 16080 26382
rect 15844 26318 15896 26324
rect 15948 26324 16028 26330
rect 15948 26318 16080 26324
rect 15856 26246 15884 26318
rect 15948 26302 16068 26318
rect 15844 26240 15896 26246
rect 15844 26182 15896 26188
rect 15856 25838 15884 26182
rect 15948 25906 15976 26302
rect 16028 26240 16080 26246
rect 16028 26182 16080 26188
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 15844 25832 15896 25838
rect 15844 25774 15896 25780
rect 15856 25430 15884 25774
rect 15844 25424 15896 25430
rect 15844 25366 15896 25372
rect 15948 25226 15976 25842
rect 16040 25226 16068 26182
rect 15936 25220 15988 25226
rect 15936 25162 15988 25168
rect 16028 25220 16080 25226
rect 16028 25162 16080 25168
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15856 24206 15884 25094
rect 16028 24336 16080 24342
rect 16028 24278 16080 24284
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15672 23769 15700 23802
rect 15936 23792 15988 23798
rect 15658 23760 15714 23769
rect 15936 23734 15988 23740
rect 15658 23695 15714 23704
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15488 23480 15608 23508
rect 15382 22400 15438 22409
rect 15382 22335 15438 22344
rect 15304 22188 15424 22216
rect 15396 22137 15424 22188
rect 15382 22128 15438 22137
rect 15382 22063 15438 22072
rect 15382 21584 15438 21593
rect 15382 21519 15438 21528
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15396 21010 15424 21519
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15212 19378 15240 20198
rect 14844 19306 14964 19334
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14740 17808 14792 17814
rect 14740 17750 14792 17756
rect 14844 16096 14872 19306
rect 14922 18184 14978 18193
rect 14922 18119 14978 18128
rect 14936 17814 14964 18119
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14924 16108 14976 16114
rect 14844 16068 14924 16096
rect 14924 16050 14976 16056
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14844 15502 14872 15574
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14936 15366 14964 16050
rect 15028 15502 15056 17614
rect 15120 17542 15148 17818
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15120 15638 15148 17478
rect 15212 17218 15240 19314
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15396 17678 15424 18906
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15290 17368 15346 17377
rect 15290 17303 15292 17312
rect 15344 17303 15346 17312
rect 15292 17274 15344 17280
rect 15212 17190 15332 17218
rect 15396 17202 15424 17478
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15212 16017 15240 17002
rect 15198 16008 15254 16017
rect 15198 15943 15254 15952
rect 15200 15904 15252 15910
rect 15304 15892 15332 17190
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15488 16114 15516 23480
rect 15856 23186 15884 23666
rect 15844 23180 15896 23186
rect 15844 23122 15896 23128
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15672 22522 15700 23054
rect 15752 22976 15804 22982
rect 15752 22918 15804 22924
rect 15764 22642 15792 22918
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15856 22545 15884 23122
rect 15948 23118 15976 23734
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15936 22772 15988 22778
rect 15936 22714 15988 22720
rect 15842 22536 15898 22545
rect 15672 22494 15792 22522
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15658 22400 15714 22409
rect 15580 22166 15608 22374
rect 15658 22335 15714 22344
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15580 21554 15608 21966
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15672 20942 15700 22335
rect 15764 22098 15792 22494
rect 15842 22471 15898 22480
rect 15948 22216 15976 22714
rect 15856 22188 15976 22216
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15750 21992 15806 22001
rect 15750 21927 15752 21936
rect 15804 21927 15806 21936
rect 15752 21898 15804 21904
rect 15856 21894 15884 22188
rect 16040 22094 16068 24278
rect 15948 22066 16068 22094
rect 15948 22012 15976 22066
rect 15948 21984 16068 22012
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15672 20398 15700 20742
rect 15764 20534 15792 20742
rect 15948 20534 15976 20878
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 15936 20528 15988 20534
rect 15936 20470 15988 20476
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15948 20058 15976 20470
rect 16040 20262 16068 21984
rect 16132 20534 16160 29446
rect 16212 29096 16264 29102
rect 16212 29038 16264 29044
rect 16224 22094 16252 29038
rect 16316 28200 16344 33408
rect 16592 32910 16620 35430
rect 16684 34746 16712 35634
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 16764 35012 16816 35018
rect 16764 34954 16816 34960
rect 16672 34740 16724 34746
rect 16672 34682 16724 34688
rect 16672 34060 16724 34066
rect 16672 34002 16724 34008
rect 16684 33590 16712 34002
rect 16672 33584 16724 33590
rect 16672 33526 16724 33532
rect 16580 32904 16632 32910
rect 16580 32846 16632 32852
rect 16776 32570 16804 34954
rect 16868 33522 16896 35022
rect 16960 34105 16988 37198
rect 17052 36378 17080 37198
rect 17316 37188 17368 37194
rect 17316 37130 17368 37136
rect 18880 37188 18932 37194
rect 18880 37130 18932 37136
rect 17224 36712 17276 36718
rect 17224 36654 17276 36660
rect 17132 36576 17184 36582
rect 17132 36518 17184 36524
rect 17040 36372 17092 36378
rect 17040 36314 17092 36320
rect 17052 35766 17080 36314
rect 17040 35760 17092 35766
rect 17040 35702 17092 35708
rect 17040 34536 17092 34542
rect 17040 34478 17092 34484
rect 17052 34377 17080 34478
rect 17038 34368 17094 34377
rect 17038 34303 17094 34312
rect 16946 34096 17002 34105
rect 16946 34031 17002 34040
rect 17144 33998 17172 36518
rect 17236 34610 17264 36654
rect 17328 35154 17356 37130
rect 17500 37120 17552 37126
rect 17500 37062 17552 37068
rect 18788 37120 18840 37126
rect 18788 37062 18840 37068
rect 17512 36786 17540 37062
rect 17776 36848 17828 36854
rect 17776 36790 17828 36796
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 17592 36780 17644 36786
rect 17592 36722 17644 36728
rect 17406 36680 17462 36689
rect 17406 36615 17462 36624
rect 17420 35630 17448 36615
rect 17408 35624 17460 35630
rect 17408 35566 17460 35572
rect 17408 35284 17460 35290
rect 17408 35226 17460 35232
rect 17316 35148 17368 35154
rect 17316 35090 17368 35096
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 17328 34202 17356 35090
rect 17420 34746 17448 35226
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 17512 34610 17540 36722
rect 17604 35222 17632 36722
rect 17684 36032 17736 36038
rect 17684 35974 17736 35980
rect 17696 35630 17724 35974
rect 17788 35698 17816 36790
rect 18800 36786 18828 37062
rect 18236 36780 18288 36786
rect 18236 36722 18288 36728
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 17868 36712 17920 36718
rect 18144 36712 18196 36718
rect 17920 36672 18144 36700
rect 17868 36654 17920 36660
rect 18144 36654 18196 36660
rect 17776 35692 17828 35698
rect 17776 35634 17828 35640
rect 17684 35624 17736 35630
rect 17684 35566 17736 35572
rect 17788 35290 17816 35634
rect 17880 35630 17908 36654
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 18144 36576 18196 36582
rect 18144 36518 18196 36524
rect 17972 36378 18000 36518
rect 17960 36372 18012 36378
rect 17960 36314 18012 36320
rect 17868 35624 17920 35630
rect 17868 35566 17920 35572
rect 17776 35284 17828 35290
rect 17776 35226 17828 35232
rect 17592 35216 17644 35222
rect 17592 35158 17644 35164
rect 17880 35086 17908 35566
rect 17868 35080 17920 35086
rect 17868 35022 17920 35028
rect 18050 34640 18106 34649
rect 17500 34604 17552 34610
rect 18050 34575 18052 34584
rect 17500 34546 17552 34552
rect 18104 34575 18106 34584
rect 18052 34546 18104 34552
rect 17316 34196 17368 34202
rect 17316 34138 17368 34144
rect 18156 33998 18184 36518
rect 18248 35834 18276 36722
rect 18328 36712 18380 36718
rect 18420 36712 18472 36718
rect 18328 36654 18380 36660
rect 18418 36680 18420 36689
rect 18696 36712 18748 36718
rect 18472 36680 18474 36689
rect 18340 36582 18368 36654
rect 18696 36654 18748 36660
rect 18418 36615 18474 36624
rect 18604 36644 18656 36650
rect 18604 36586 18656 36592
rect 18328 36576 18380 36582
rect 18328 36518 18380 36524
rect 18420 36236 18472 36242
rect 18420 36178 18472 36184
rect 18328 36100 18380 36106
rect 18328 36042 18380 36048
rect 18236 35828 18288 35834
rect 18236 35770 18288 35776
rect 18340 35766 18368 36042
rect 18328 35760 18380 35766
rect 18328 35702 18380 35708
rect 18432 35698 18460 36178
rect 18512 36100 18564 36106
rect 18512 36042 18564 36048
rect 18420 35692 18472 35698
rect 18420 35634 18472 35640
rect 18432 35154 18460 35634
rect 18420 35148 18472 35154
rect 18420 35090 18472 35096
rect 18432 34610 18460 35090
rect 18420 34604 18472 34610
rect 18420 34546 18472 34552
rect 18524 34082 18552 36042
rect 18616 36038 18644 36586
rect 18708 36242 18736 36654
rect 18788 36576 18840 36582
rect 18788 36518 18840 36524
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 18604 36032 18656 36038
rect 18604 35974 18656 35980
rect 18800 35766 18828 36518
rect 18788 35760 18840 35766
rect 18788 35702 18840 35708
rect 18892 35612 18920 37130
rect 20168 37120 20220 37126
rect 20168 37062 20220 37068
rect 19616 36712 19668 36718
rect 19616 36654 19668 36660
rect 19628 36378 19656 36654
rect 19616 36372 19668 36378
rect 19616 36314 19668 36320
rect 18984 36230 19196 36258
rect 20180 36242 20208 37062
rect 18984 36038 19012 36230
rect 19064 36168 19116 36174
rect 19064 36110 19116 36116
rect 18972 36032 19024 36038
rect 18972 35974 19024 35980
rect 19076 35986 19104 36110
rect 19168 36106 19196 36230
rect 19248 36236 19300 36242
rect 19248 36178 19300 36184
rect 19800 36236 19852 36242
rect 19800 36178 19852 36184
rect 20168 36236 20220 36242
rect 20168 36178 20220 36184
rect 20260 36236 20312 36242
rect 20260 36178 20312 36184
rect 19260 36145 19288 36178
rect 19340 36168 19392 36174
rect 19246 36136 19302 36145
rect 19156 36100 19208 36106
rect 19524 36168 19576 36174
rect 19392 36128 19524 36156
rect 19340 36110 19392 36116
rect 19246 36071 19302 36080
rect 19156 36042 19208 36048
rect 19248 36032 19300 36038
rect 19076 35980 19248 35986
rect 19076 35974 19300 35980
rect 19076 35958 19288 35974
rect 18800 35584 18920 35612
rect 18696 35216 18748 35222
rect 18696 35158 18748 35164
rect 18604 34468 18656 34474
rect 18604 34410 18656 34416
rect 18328 34060 18380 34066
rect 18328 34002 18380 34008
rect 18432 34054 18552 34082
rect 17132 33992 17184 33998
rect 17132 33934 17184 33940
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 18156 33561 18184 33934
rect 18142 33552 18198 33561
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 18052 33516 18104 33522
rect 18142 33487 18198 33496
rect 18052 33458 18104 33464
rect 16764 32564 16816 32570
rect 16764 32506 16816 32512
rect 16580 32496 16632 32502
rect 16580 32438 16632 32444
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 16408 30569 16436 32370
rect 16486 30832 16542 30841
rect 16486 30767 16542 30776
rect 16394 30560 16450 30569
rect 16394 30495 16450 30504
rect 16396 29232 16448 29238
rect 16396 29174 16448 29180
rect 16408 28558 16436 29174
rect 16500 28762 16528 30767
rect 16592 29714 16620 32438
rect 16868 31142 16896 33458
rect 18064 33153 18092 33458
rect 18050 33144 18106 33153
rect 18248 33114 18276 33934
rect 18340 33658 18368 34002
rect 18328 33652 18380 33658
rect 18328 33594 18380 33600
rect 18432 33454 18460 34054
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 18524 33658 18552 33934
rect 18512 33652 18564 33658
rect 18512 33594 18564 33600
rect 18524 33522 18552 33594
rect 18616 33522 18644 34410
rect 18708 33522 18736 35158
rect 18800 34377 18828 35584
rect 19260 34746 19288 35958
rect 19248 34740 19300 34746
rect 19248 34682 19300 34688
rect 19444 34610 19472 36128
rect 19812 36145 19840 36178
rect 19524 36110 19576 36116
rect 19798 36136 19854 36145
rect 20272 36106 20300 36178
rect 19798 36071 19854 36080
rect 20260 36100 20312 36106
rect 20260 36042 20312 36048
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 19892 35488 19944 35494
rect 19892 35430 19944 35436
rect 19616 35148 19668 35154
rect 19616 35090 19668 35096
rect 19628 35018 19656 35090
rect 19616 35012 19668 35018
rect 19616 34954 19668 34960
rect 19156 34604 19208 34610
rect 19156 34546 19208 34552
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 18880 34536 18932 34542
rect 18880 34478 18932 34484
rect 18786 34368 18842 34377
rect 18786 34303 18842 34312
rect 18512 33516 18564 33522
rect 18512 33458 18564 33464
rect 18604 33516 18656 33522
rect 18604 33458 18656 33464
rect 18696 33516 18748 33522
rect 18696 33458 18748 33464
rect 18420 33448 18472 33454
rect 18420 33390 18472 33396
rect 18050 33079 18106 33088
rect 18236 33108 18288 33114
rect 18236 33050 18288 33056
rect 18328 33108 18380 33114
rect 18328 33050 18380 33056
rect 18340 32502 18368 33050
rect 18616 33017 18644 33458
rect 18800 33454 18828 34303
rect 18892 33522 18920 34478
rect 18972 34400 19024 34406
rect 18972 34342 19024 34348
rect 18984 33998 19012 34342
rect 18972 33992 19024 33998
rect 18972 33934 19024 33940
rect 18984 33590 19012 33934
rect 19168 33590 19196 34546
rect 19628 34490 19656 34954
rect 19904 34678 19932 35430
rect 20168 35012 20220 35018
rect 20168 34954 20220 34960
rect 20180 34921 20208 34954
rect 20166 34912 20222 34921
rect 20166 34847 20222 34856
rect 20364 34678 20392 35634
rect 21100 35630 21128 37266
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 21916 37120 21968 37126
rect 21916 37062 21968 37068
rect 21928 36242 21956 37062
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 21916 36236 21968 36242
rect 21916 36178 21968 36184
rect 22112 36106 22140 36722
rect 22204 36582 22232 37130
rect 22192 36576 22244 36582
rect 22192 36518 22244 36524
rect 22190 36272 22246 36281
rect 22190 36207 22192 36216
rect 22244 36207 22246 36216
rect 22192 36178 22244 36184
rect 22100 36100 22152 36106
rect 22100 36042 22152 36048
rect 21548 36032 21600 36038
rect 21548 35974 21600 35980
rect 21364 35692 21416 35698
rect 21364 35634 21416 35640
rect 21088 35624 21140 35630
rect 21088 35566 21140 35572
rect 19892 34672 19944 34678
rect 19892 34614 19944 34620
rect 20352 34672 20404 34678
rect 20352 34614 20404 34620
rect 19536 34474 19656 34490
rect 19524 34468 19656 34474
rect 19576 34462 19656 34468
rect 19524 34410 19576 34416
rect 19248 34400 19300 34406
rect 19248 34342 19300 34348
rect 19260 33658 19288 34342
rect 19536 34066 19564 34410
rect 19524 34060 19576 34066
rect 19524 34002 19576 34008
rect 19248 33652 19300 33658
rect 19248 33594 19300 33600
rect 18972 33584 19024 33590
rect 18972 33526 19024 33532
rect 19156 33584 19208 33590
rect 19156 33526 19208 33532
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 18788 33448 18840 33454
rect 18788 33390 18840 33396
rect 19156 33448 19208 33454
rect 19156 33390 19208 33396
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 18696 33380 18748 33386
rect 18696 33322 18748 33328
rect 18602 33008 18658 33017
rect 18602 32943 18658 32952
rect 17500 32496 17552 32502
rect 18328 32496 18380 32502
rect 17552 32456 17908 32484
rect 17500 32438 17552 32444
rect 17880 32450 17908 32456
rect 17880 32434 18092 32450
rect 18328 32438 18380 32444
rect 17880 32428 18104 32434
rect 17880 32422 18052 32428
rect 18052 32370 18104 32376
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 17684 32360 17736 32366
rect 17684 32302 17736 32308
rect 17960 32360 18012 32366
rect 17960 32302 18012 32308
rect 17500 32224 17552 32230
rect 17500 32166 17552 32172
rect 17408 31952 17460 31958
rect 17408 31894 17460 31900
rect 17316 31748 17368 31754
rect 17316 31690 17368 31696
rect 17328 31142 17356 31690
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 17316 31136 17368 31142
rect 17316 31078 17368 31084
rect 16868 30122 16896 31078
rect 17132 30592 17184 30598
rect 17132 30534 17184 30540
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 16856 30116 16908 30122
rect 16856 30058 16908 30064
rect 16868 29974 17080 30002
rect 16670 29880 16726 29889
rect 16670 29815 16726 29824
rect 16580 29708 16632 29714
rect 16580 29650 16632 29656
rect 16684 29510 16712 29815
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16764 29504 16816 29510
rect 16764 29446 16816 29452
rect 16776 29238 16804 29446
rect 16764 29232 16816 29238
rect 16764 29174 16816 29180
rect 16580 28960 16632 28966
rect 16580 28902 16632 28908
rect 16488 28756 16540 28762
rect 16488 28698 16540 28704
rect 16396 28552 16448 28558
rect 16396 28494 16448 28500
rect 16408 28422 16436 28494
rect 16396 28416 16448 28422
rect 16396 28358 16448 28364
rect 16316 28172 16436 28200
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16316 27470 16344 28018
rect 16408 27985 16436 28172
rect 16500 28014 16528 28698
rect 16592 28558 16620 28902
rect 16776 28626 16804 29174
rect 16868 29170 16896 29974
rect 16946 29880 17002 29889
rect 16946 29815 17002 29824
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16856 28688 16908 28694
rect 16856 28630 16908 28636
rect 16764 28620 16816 28626
rect 16764 28562 16816 28568
rect 16580 28552 16632 28558
rect 16672 28552 16724 28558
rect 16580 28494 16632 28500
rect 16670 28520 16672 28529
rect 16724 28520 16726 28529
rect 16670 28455 16726 28464
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 16488 28008 16540 28014
rect 16394 27976 16450 27985
rect 16488 27950 16540 27956
rect 16394 27911 16450 27920
rect 16592 27826 16620 28358
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16500 27798 16620 27826
rect 16304 27464 16356 27470
rect 16304 27406 16356 27412
rect 16316 27334 16344 27406
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 16500 27130 16528 27798
rect 16488 27124 16540 27130
rect 16488 27066 16540 27072
rect 16394 27024 16450 27033
rect 16394 26959 16396 26968
rect 16448 26959 16450 26968
rect 16396 26930 16448 26936
rect 16396 26240 16448 26246
rect 16396 26182 16448 26188
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16316 24954 16344 25230
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16302 24168 16358 24177
rect 16302 24103 16358 24112
rect 16316 23118 16344 24103
rect 16408 23866 16436 26182
rect 16500 25770 16528 27066
rect 16580 26988 16632 26994
rect 16580 26930 16632 26936
rect 16488 25764 16540 25770
rect 16488 25706 16540 25712
rect 16592 24857 16620 26930
rect 16684 26081 16712 28018
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16670 26072 16726 26081
rect 16670 26007 16726 26016
rect 16672 25968 16724 25974
rect 16672 25910 16724 25916
rect 16684 25226 16712 25910
rect 16776 25294 16804 26182
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16578 24848 16634 24857
rect 16684 24818 16712 25162
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16578 24783 16634 24792
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16670 24712 16726 24721
rect 16670 24647 16726 24656
rect 16488 24268 16540 24274
rect 16488 24210 16540 24216
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16500 23254 16528 24210
rect 16488 23248 16540 23254
rect 16488 23190 16540 23196
rect 16304 23112 16356 23118
rect 16302 23080 16304 23089
rect 16356 23080 16358 23089
rect 16302 23015 16358 23024
rect 16500 22574 16528 23190
rect 16684 23100 16712 24647
rect 16592 23072 16712 23100
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16224 22066 16344 22094
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16224 20641 16252 21830
rect 16210 20632 16266 20641
rect 16210 20567 16266 20576
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 16316 20346 16344 22066
rect 16500 22030 16528 22374
rect 16592 22137 16620 23072
rect 16578 22128 16634 22137
rect 16776 22094 16804 25094
rect 16868 23118 16896 28630
rect 16960 28082 16988 29815
rect 17052 29646 17080 29974
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 17052 29102 17080 29446
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17144 28490 17172 30534
rect 17236 29730 17264 30534
rect 17328 29850 17356 31078
rect 17316 29844 17368 29850
rect 17316 29786 17368 29792
rect 17236 29702 17356 29730
rect 17420 29714 17448 31894
rect 17512 31822 17540 32166
rect 17696 32026 17724 32302
rect 17684 32020 17736 32026
rect 17684 31962 17736 31968
rect 17868 31952 17920 31958
rect 17604 31900 17868 31906
rect 17604 31894 17920 31900
rect 17604 31878 17908 31894
rect 17500 31816 17552 31822
rect 17500 31758 17552 31764
rect 17604 31414 17632 31878
rect 17868 31816 17920 31822
rect 17868 31758 17920 31764
rect 17776 31680 17828 31686
rect 17776 31622 17828 31628
rect 17788 31414 17816 31622
rect 17592 31408 17644 31414
rect 17592 31350 17644 31356
rect 17776 31408 17828 31414
rect 17776 31350 17828 31356
rect 17592 31136 17644 31142
rect 17592 31078 17644 31084
rect 17604 30258 17632 31078
rect 17684 30660 17736 30666
rect 17684 30602 17736 30608
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17222 29200 17278 29209
rect 17222 29135 17224 29144
rect 17276 29135 17278 29144
rect 17224 29106 17276 29112
rect 17224 29028 17276 29034
rect 17224 28970 17276 28976
rect 17132 28484 17184 28490
rect 17132 28426 17184 28432
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 16948 27600 17000 27606
rect 16948 27542 17000 27548
rect 16960 26790 16988 27542
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17040 27396 17092 27402
rect 17040 27338 17092 27344
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 16960 26586 16988 26726
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 17052 26518 17080 27338
rect 17040 26512 17092 26518
rect 17040 26454 17092 26460
rect 16948 26376 17000 26382
rect 16946 26344 16948 26353
rect 17000 26344 17002 26353
rect 16946 26279 17002 26288
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16960 24721 16988 25230
rect 16946 24712 17002 24721
rect 16946 24647 17002 24656
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 16960 24449 16988 24550
rect 16946 24440 17002 24449
rect 16946 24375 17002 24384
rect 17052 23594 17080 24550
rect 17040 23588 17092 23594
rect 17040 23530 17092 23536
rect 17052 23361 17080 23530
rect 17038 23352 17094 23361
rect 17038 23287 17040 23296
rect 17092 23287 17094 23296
rect 17040 23258 17092 23264
rect 16856 23112 16908 23118
rect 16948 23112 17000 23118
rect 16856 23054 16908 23060
rect 16946 23080 16948 23089
rect 17000 23080 17002 23089
rect 16946 23015 17002 23024
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 17052 22953 17080 22986
rect 17038 22944 17094 22953
rect 17038 22879 17094 22888
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 16578 22063 16634 22072
rect 16684 22066 16804 22094
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16408 21865 16436 21898
rect 16394 21856 16450 21865
rect 16394 21791 16450 21800
rect 16396 21072 16448 21078
rect 16396 21014 16448 21020
rect 16408 20874 16436 21014
rect 16396 20868 16448 20874
rect 16396 20810 16448 20816
rect 16224 20318 16344 20346
rect 16408 20330 16436 20810
rect 16500 20534 16528 21966
rect 16580 21548 16632 21554
rect 16684 21536 16712 22066
rect 16762 21992 16818 22001
rect 16762 21927 16818 21936
rect 16632 21508 16712 21536
rect 16580 21490 16632 21496
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16396 20324 16448 20330
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15252 15864 15332 15892
rect 15200 15846 15252 15852
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14936 15094 14964 15302
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 14936 14618 14964 15030
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 13938 14780 14214
rect 15014 13968 15070 13977
rect 14740 13932 14792 13938
rect 15014 13903 15070 13912
rect 14740 13874 14792 13880
rect 14752 13530 14780 13874
rect 15028 13870 15056 13903
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 13734 15056 13806
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13569 15056 13670
rect 15014 13560 15070 13569
rect 14740 13524 14792 13530
rect 15014 13495 15070 13504
rect 14740 13466 14792 13472
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14660 12646 14688 13330
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14844 12696 14872 12786
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 14752 12668 14872 12696
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11762 14596 12038
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14554 11520 14610 11529
rect 14554 11455 14610 11464
rect 14568 11150 14596 11455
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14462 10704 14518 10713
rect 14462 10639 14518 10648
rect 14292 10016 14412 10044
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 13832 9132 13952 9160
rect 13818 9072 13874 9081
rect 13740 9030 13818 9058
rect 13818 9007 13874 9016
rect 13832 8022 13860 9007
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13832 7818 13860 7958
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 7002 13400 7686
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6662 13400 6734
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13096 4672 13124 5238
rect 13360 4684 13412 4690
rect 13096 4644 13360 4672
rect 13360 4626 13412 4632
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12728 3534 12756 4150
rect 12820 4078 12848 4422
rect 13464 4214 13492 7482
rect 13818 7304 13874 7313
rect 13818 7239 13874 7248
rect 13832 7002 13860 7239
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13556 6458 13584 6870
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13634 6624 13690 6633
rect 13634 6559 13690 6568
rect 13648 6458 13676 6559
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13832 6361 13860 6802
rect 13924 6662 13952 9132
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13818 6352 13874 6361
rect 13818 6287 13820 6296
rect 13872 6287 13874 6296
rect 13820 6258 13872 6264
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13542 5672 13598 5681
rect 13542 5607 13598 5616
rect 13556 5574 13584 5607
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12452 2650 12480 2994
rect 12728 2774 12756 3470
rect 12636 2746 12756 2774
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12636 2496 12664 2746
rect 11940 2468 12020 2496
rect 12544 2468 12664 2496
rect 11888 2450 11940 2456
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 12544 2378 12572 2468
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 11624 800 11652 2042
rect 12176 1170 12204 2246
rect 12176 1142 12296 1170
rect 12268 800 12296 1142
rect 12912 800 12940 3674
rect 13360 3596 13412 3602
rect 13280 3556 13360 3584
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3194 13032 3470
rect 13280 3398 13308 3556
rect 13360 3538 13412 3544
rect 13464 3534 13492 3878
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13280 3126 13308 3334
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13556 2774 13584 4966
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13648 4282 13676 4558
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13740 3602 13768 6190
rect 13924 6186 13952 6598
rect 14108 6458 14136 9522
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 9110 14228 9318
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14186 7984 14242 7993
rect 14186 7919 14242 7928
rect 14200 7886 14228 7919
rect 14292 7886 14320 8230
rect 14384 8090 14412 10016
rect 14476 9738 14504 10639
rect 14568 9926 14596 11086
rect 14660 11014 14688 11086
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14476 9710 14596 9738
rect 14660 9722 14688 10950
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14476 8498 14504 9318
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14200 7546 14228 7822
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14568 7478 14596 9710
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14752 9586 14780 12668
rect 14936 12594 14964 12718
rect 14844 12566 14964 12594
rect 14844 9586 14872 12566
rect 15028 10470 15056 13126
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15028 9722 15056 9998
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14752 7954 14780 9522
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14752 7478 14780 7890
rect 15120 7886 15148 15574
rect 15212 14958 15240 15846
rect 15488 15502 15516 16050
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15212 11762 15240 12174
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11082 15240 11494
rect 15304 11218 15332 13670
rect 15396 12442 15424 15302
rect 15488 15026 15516 15438
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 9586 15240 11018
rect 15304 10674 15332 11154
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15396 10062 15424 12378
rect 15488 12322 15516 14758
rect 15580 12442 15608 19314
rect 15672 18222 15700 19926
rect 16132 19922 16160 20198
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15750 19272 15806 19281
rect 15750 19207 15806 19216
rect 15764 18766 15792 19207
rect 15948 18834 15976 19790
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15764 17678 15792 18362
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15672 16522 15700 17138
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15750 16144 15806 16153
rect 15750 16079 15806 16088
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15672 15026 15700 15370
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15764 14074 15792 16079
rect 15948 15910 15976 18770
rect 16040 17796 16068 19654
rect 16224 19446 16252 20318
rect 16396 20266 16448 20272
rect 16304 20256 16356 20262
rect 16592 20210 16620 21490
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16684 20369 16712 20402
rect 16776 20398 16804 21927
rect 16764 20392 16816 20398
rect 16670 20360 16726 20369
rect 16764 20334 16816 20340
rect 16670 20295 16726 20304
rect 16960 20262 16988 22714
rect 17144 21146 17172 27406
rect 17236 26994 17264 28970
rect 17328 28082 17356 29702
rect 17408 29708 17460 29714
rect 17408 29650 17460 29656
rect 17408 28484 17460 28490
rect 17408 28426 17460 28432
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 17420 26994 17448 28426
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 17512 27606 17540 28018
rect 17500 27600 17552 27606
rect 17500 27542 17552 27548
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 17316 26920 17368 26926
rect 17512 26874 17540 26930
rect 17316 26862 17368 26868
rect 17224 26512 17276 26518
rect 17224 26454 17276 26460
rect 17236 24138 17264 26454
rect 17328 26353 17356 26862
rect 17420 26846 17540 26874
rect 17314 26344 17370 26353
rect 17314 26279 17316 26288
rect 17368 26279 17370 26288
rect 17316 26250 17368 26256
rect 17314 26072 17370 26081
rect 17314 26007 17370 26016
rect 17328 24682 17356 26007
rect 17316 24676 17368 24682
rect 17316 24618 17368 24624
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17236 23338 17264 24074
rect 17420 23526 17448 26846
rect 17498 26344 17554 26353
rect 17498 26279 17500 26288
rect 17552 26279 17554 26288
rect 17500 26250 17552 26256
rect 17604 26194 17632 30194
rect 17696 30190 17724 30602
rect 17684 30184 17736 30190
rect 17684 30126 17736 30132
rect 17696 29646 17724 30126
rect 17684 29640 17736 29646
rect 17684 29582 17736 29588
rect 17696 29102 17724 29582
rect 17788 29578 17816 31350
rect 17880 31346 17908 31758
rect 17972 31754 18000 32302
rect 18432 31754 18460 32370
rect 18708 31890 18736 33322
rect 18880 32564 18932 32570
rect 18880 32506 18932 32512
rect 18696 31884 18748 31890
rect 18696 31826 18748 31832
rect 17972 31726 18184 31754
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17880 30938 17908 31282
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17868 30660 17920 30666
rect 17868 30602 17920 30608
rect 17880 30569 17908 30602
rect 17866 30560 17922 30569
rect 17866 30495 17922 30504
rect 17972 29646 18000 30670
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 17776 29572 17828 29578
rect 17776 29514 17828 29520
rect 17868 29572 17920 29578
rect 17868 29514 17920 29520
rect 17788 29170 17816 29514
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17684 29096 17736 29102
rect 17684 29038 17736 29044
rect 17880 28218 17908 29514
rect 17972 29510 18000 29582
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 18064 29170 18092 31214
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18064 29034 18092 29106
rect 18052 29028 18104 29034
rect 18052 28970 18104 28976
rect 18156 28914 18184 31726
rect 18420 31748 18472 31754
rect 18420 31690 18472 31696
rect 18604 30320 18656 30326
rect 18604 30262 18656 30268
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 18340 29782 18368 30126
rect 18328 29776 18380 29782
rect 18328 29718 18380 29724
rect 18524 29730 18552 30194
rect 18616 29850 18644 30262
rect 18604 29844 18656 29850
rect 18604 29786 18656 29792
rect 18524 29702 18644 29730
rect 18512 29640 18564 29646
rect 18512 29582 18564 29588
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 18236 29504 18288 29510
rect 18236 29446 18288 29452
rect 18248 29209 18276 29446
rect 18234 29200 18290 29209
rect 18234 29135 18290 29144
rect 18064 28886 18184 28914
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17512 26166 17632 26194
rect 17408 23520 17460 23526
rect 17406 23488 17408 23497
rect 17460 23488 17462 23497
rect 17406 23423 17462 23432
rect 17236 23310 17448 23338
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17236 21690 17264 22170
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17328 21622 17356 22102
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17328 21146 17356 21286
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 17040 20936 17092 20942
rect 17038 20904 17040 20913
rect 17092 20904 17094 20913
rect 17038 20839 17094 20848
rect 17040 20392 17092 20398
rect 17040 20334 17092 20340
rect 16304 20198 16356 20204
rect 16212 19440 16264 19446
rect 16212 19382 16264 19388
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16132 18057 16160 18702
rect 16224 18630 16252 19382
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16118 18048 16174 18057
rect 16118 17983 16174 17992
rect 16040 17768 16160 17796
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 16040 15706 16068 17614
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15764 12782 15792 13262
rect 15856 12850 15884 15438
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15764 12374 15792 12718
rect 15752 12368 15804 12374
rect 15488 12294 15700 12322
rect 15752 12310 15804 12316
rect 15488 11830 15516 12294
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15488 10266 15516 10610
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15580 10266 15608 10542
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15580 9518 15608 10202
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 6798 14320 7346
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14660 6662 14688 7278
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14660 6322 14688 6598
rect 15120 6390 15148 7822
rect 15212 7478 15240 9318
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15396 7886 15424 8026
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15198 6896 15254 6905
rect 15198 6831 15254 6840
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13832 4146 13860 5102
rect 13924 5098 13952 5782
rect 15212 5710 15240 6831
rect 15396 6118 15424 7142
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13832 3126 13860 4082
rect 14016 3670 14044 5646
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14188 5296 14240 5302
rect 14372 5296 14424 5302
rect 14240 5256 14372 5284
rect 14188 5238 14240 5244
rect 14372 5238 14424 5244
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14384 4758 14412 4966
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13556 2746 13676 2774
rect 13648 2446 13676 2746
rect 13740 2650 13768 2926
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13832 2514 13860 3062
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 14016 2446 14044 3606
rect 14200 3466 14228 3606
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 14292 2990 14320 4558
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 13556 800 13584 2382
rect 14384 2378 14412 4150
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14476 3738 14504 4014
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14568 3602 14596 5510
rect 14752 3602 14780 5646
rect 15304 5166 15332 6054
rect 15488 5710 15516 6054
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15580 5574 15608 7754
rect 15672 6322 15700 12294
rect 15764 11762 15792 12310
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15856 9382 15884 12786
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15948 8378 15976 12378
rect 16132 8634 16160 17768
rect 16316 17202 16344 20198
rect 16500 20182 16620 20210
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16408 19514 16436 19790
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16408 19174 16436 19450
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16500 18714 16528 20182
rect 16762 20088 16818 20097
rect 16580 20052 16632 20058
rect 16762 20023 16818 20032
rect 16580 19994 16632 20000
rect 16592 18834 16620 19994
rect 16776 19786 16804 20023
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16960 19666 16988 20198
rect 17052 19786 17080 20334
rect 17144 19854 17172 21082
rect 17224 20256 17276 20262
rect 17222 20224 17224 20233
rect 17276 20224 17278 20233
rect 17222 20159 17278 20168
rect 17328 19938 17356 21082
rect 17420 20058 17448 23310
rect 17512 22778 17540 26166
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17604 24342 17632 24686
rect 17592 24336 17644 24342
rect 17592 24278 17644 24284
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17604 23322 17632 24006
rect 17696 23866 17724 28018
rect 17880 25838 17908 28154
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17972 26994 18000 27814
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 18064 25786 18092 28886
rect 18248 28529 18276 29135
rect 18234 28520 18290 28529
rect 18234 28455 18290 28464
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 18156 26586 18184 26930
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 18248 26489 18276 28086
rect 18328 27328 18380 27334
rect 18328 27270 18380 27276
rect 18234 26480 18290 26489
rect 18144 26444 18196 26450
rect 18234 26415 18290 26424
rect 18144 26386 18196 26392
rect 18156 25906 18184 26386
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18064 25758 18276 25786
rect 17868 25696 17920 25702
rect 17920 25644 18000 25650
rect 17868 25638 18000 25644
rect 17880 25622 18000 25638
rect 17972 24818 18000 25622
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17880 24410 17908 24550
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 17776 24336 17828 24342
rect 17776 24278 17828 24284
rect 17788 24138 17816 24278
rect 17972 24274 18000 24550
rect 17960 24268 18012 24274
rect 17960 24210 18012 24216
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 18064 24018 18092 24210
rect 17788 23990 18092 24018
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17696 23322 17724 23802
rect 17788 23594 17816 23990
rect 18144 23860 18196 23866
rect 17972 23820 18144 23848
rect 17868 23792 17920 23798
rect 17972 23746 18000 23820
rect 18144 23802 18196 23808
rect 18248 23746 18276 25758
rect 17920 23740 18000 23746
rect 17868 23734 18000 23740
rect 17880 23718 18000 23734
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17868 23520 17920 23526
rect 17774 23488 17830 23497
rect 17868 23462 17920 23468
rect 17774 23423 17830 23432
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17604 22658 17632 23258
rect 17788 23168 17816 23423
rect 17880 23361 17908 23462
rect 17866 23352 17922 23361
rect 17866 23287 17922 23296
rect 17972 23186 18000 23718
rect 18064 23718 18276 23746
rect 17696 23140 17816 23168
rect 17960 23180 18012 23186
rect 17696 22982 17724 23140
rect 17960 23122 18012 23128
rect 17776 23044 17828 23050
rect 17776 22986 17828 22992
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17512 22630 17632 22658
rect 17512 20262 17540 22630
rect 17696 22556 17724 22918
rect 17604 22528 17724 22556
rect 17604 20534 17632 22528
rect 17682 22128 17738 22137
rect 17682 22063 17738 22072
rect 17696 21622 17724 22063
rect 17788 22001 17816 22986
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17774 21992 17830 22001
rect 17774 21927 17830 21936
rect 17880 21706 17908 22646
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17972 22234 18000 22578
rect 17960 22228 18012 22234
rect 17960 22170 18012 22176
rect 17788 21678 17908 21706
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 17592 20528 17644 20534
rect 17590 20496 17592 20505
rect 17644 20496 17646 20505
rect 17590 20431 17646 20440
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17328 19910 17448 19938
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17132 19712 17184 19718
rect 16960 19660 17132 19666
rect 16960 19654 17184 19660
rect 16684 18902 16712 19654
rect 16960 19638 17172 19654
rect 16762 19408 16818 19417
rect 16762 19343 16818 19352
rect 16776 19310 16804 19343
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16776 19009 16804 19110
rect 16762 19000 16818 19009
rect 16762 18935 16764 18944
rect 16816 18935 16818 18944
rect 16764 18906 16816 18912
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16672 18760 16724 18766
rect 16500 18686 16620 18714
rect 16672 18702 16724 18708
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16224 14550 16252 14894
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 15856 8350 15976 8378
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15764 7546 15792 7754
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15856 6186 15884 8350
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15948 7886 15976 8230
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15672 5302 15700 5646
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 14832 3936 14884 3942
rect 15028 3924 15056 5102
rect 15672 4826 15700 5238
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 14884 3896 15056 3924
rect 14832 3878 14884 3884
rect 15028 3602 15056 3896
rect 15304 3738 15332 4762
rect 15672 4078 15700 4762
rect 15764 4690 15792 6122
rect 15856 5642 15884 6122
rect 16224 5914 16252 6326
rect 16316 6254 16344 13874
rect 16408 9178 16436 17002
rect 16592 13326 16620 18686
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16500 12918 16528 13262
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11393 16528 12106
rect 16486 11384 16542 11393
rect 16486 11319 16542 11328
rect 16500 11218 16528 11319
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16592 9908 16620 13262
rect 16684 12102 16712 18702
rect 16776 12434 16804 18906
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16868 18358 16896 18566
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16960 17610 16988 19638
rect 17038 19544 17094 19553
rect 17038 19479 17094 19488
rect 17052 18766 17080 19479
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17144 17954 17172 19314
rect 17144 17926 17264 17954
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16960 15434 16988 15914
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16960 14074 16988 15370
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16960 13938 16988 14010
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16776 12406 16896 12434
rect 16762 12200 16818 12209
rect 16762 12135 16818 12144
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16670 11928 16726 11937
rect 16776 11898 16804 12135
rect 16670 11863 16672 11872
rect 16724 11863 16726 11872
rect 16764 11892 16816 11898
rect 16672 11834 16724 11840
rect 16868 11880 16896 12406
rect 16868 11852 16988 11880
rect 16764 11834 16816 11840
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16776 11558 16804 11630
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16672 11144 16724 11150
rect 16670 11112 16672 11121
rect 16724 11112 16726 11121
rect 16670 11047 16726 11056
rect 16500 9880 16620 9908
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16394 8392 16450 8401
rect 16394 8327 16450 8336
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16316 5914 16344 6190
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16408 5710 16436 8327
rect 16500 7410 16528 9880
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16486 7304 16542 7313
rect 16486 7239 16542 7248
rect 16500 5710 16528 7239
rect 16592 7206 16620 9046
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16684 7546 16712 8366
rect 16776 8362 16804 11494
rect 16868 11354 16896 11698
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16960 8616 16988 11852
rect 17052 10198 17080 17478
rect 17130 16280 17186 16289
rect 17130 16215 17132 16224
rect 17184 16215 17186 16224
rect 17132 16186 17184 16192
rect 17236 16182 17264 17926
rect 17420 17678 17448 19910
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17696 19378 17724 19722
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17788 18850 17816 21678
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17880 20806 17908 21558
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17880 19922 17908 20742
rect 17972 20097 18000 20878
rect 17958 20088 18014 20097
rect 17958 20023 18014 20032
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17972 19394 18000 20023
rect 17512 18822 17816 18850
rect 17880 19366 18000 19394
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17144 13530 17172 13874
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17130 12336 17186 12345
rect 17236 12306 17264 15982
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17328 13938 17356 15302
rect 17420 15026 17448 17614
rect 17512 15434 17540 18822
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17604 17270 17632 17682
rect 17696 17678 17724 18634
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17592 17264 17644 17270
rect 17592 17206 17644 17212
rect 17604 16114 17632 17206
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17696 15162 17724 17614
rect 17880 15366 17908 19366
rect 18064 18154 18092 23718
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18156 23225 18184 23462
rect 18236 23248 18288 23254
rect 18142 23216 18198 23225
rect 18236 23190 18288 23196
rect 18142 23151 18198 23160
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 18156 20482 18184 22918
rect 18248 22681 18276 23190
rect 18234 22672 18290 22681
rect 18234 22607 18236 22616
rect 18288 22607 18290 22616
rect 18236 22578 18288 22584
rect 18340 22574 18368 27270
rect 18432 26058 18460 29514
rect 18524 29306 18552 29582
rect 18512 29300 18564 29306
rect 18512 29242 18564 29248
rect 18616 28626 18644 29702
rect 18604 28620 18656 28626
rect 18604 28562 18656 28568
rect 18708 27402 18736 31826
rect 18892 31346 18920 32506
rect 19168 31754 19196 33390
rect 19444 33318 19472 33390
rect 19536 33386 19564 34002
rect 20364 33946 20392 34614
rect 20272 33930 20392 33946
rect 20260 33924 20392 33930
rect 20312 33918 20392 33924
rect 20260 33866 20312 33872
rect 20272 33658 20300 33866
rect 20260 33652 20312 33658
rect 20260 33594 20312 33600
rect 19524 33380 19576 33386
rect 19524 33322 19576 33328
rect 19432 33312 19484 33318
rect 19432 33254 19484 33260
rect 19248 32836 19300 32842
rect 19248 32778 19300 32784
rect 19260 32434 19288 32778
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19352 32434 19380 32710
rect 19444 32552 19472 33254
rect 20074 33008 20130 33017
rect 19892 32972 19944 32978
rect 20074 32943 20130 32952
rect 19892 32914 19944 32920
rect 19904 32570 19932 32914
rect 20088 32910 20116 32943
rect 20076 32904 20128 32910
rect 20260 32904 20312 32910
rect 20076 32846 20128 32852
rect 20258 32872 20260 32881
rect 20312 32872 20314 32881
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19800 32564 19852 32570
rect 19444 32524 19564 32552
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19260 31890 19288 32370
rect 19340 32292 19392 32298
rect 19340 32234 19392 32240
rect 19248 31884 19300 31890
rect 19248 31826 19300 31832
rect 19168 31726 19288 31754
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 18880 31340 18932 31346
rect 18880 31282 18932 31288
rect 18800 31142 18828 31282
rect 18788 31136 18840 31142
rect 18788 31078 18840 31084
rect 18892 30734 18920 31282
rect 19156 31204 19208 31210
rect 19156 31146 19208 31152
rect 18880 30728 18932 30734
rect 18932 30688 19012 30716
rect 18880 30670 18932 30676
rect 18880 30592 18932 30598
rect 18880 30534 18932 30540
rect 18892 30258 18920 30534
rect 18984 30326 19012 30688
rect 19168 30598 19196 31146
rect 19260 30666 19288 31726
rect 19352 31482 19380 32234
rect 19444 31958 19472 32370
rect 19432 31952 19484 31958
rect 19432 31894 19484 31900
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19248 30660 19300 30666
rect 19248 30602 19300 30608
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 19260 30410 19288 30602
rect 19064 30388 19116 30394
rect 19064 30330 19116 30336
rect 19168 30382 19288 30410
rect 18972 30320 19024 30326
rect 18972 30262 19024 30268
rect 18880 30252 18932 30258
rect 18880 30194 18932 30200
rect 18788 29776 18840 29782
rect 18788 29718 18840 29724
rect 18800 28558 18828 29718
rect 18892 28642 18920 30194
rect 18972 30184 19024 30190
rect 18972 30126 19024 30132
rect 18984 29850 19012 30126
rect 18972 29844 19024 29850
rect 18972 29786 19024 29792
rect 19076 29306 19104 30330
rect 19064 29300 19116 29306
rect 19064 29242 19116 29248
rect 19168 29186 19196 30382
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 18972 29164 19024 29170
rect 18972 29106 19024 29112
rect 19076 29158 19196 29186
rect 18984 29073 19012 29106
rect 18970 29064 19026 29073
rect 18970 28999 19026 29008
rect 19076 28994 19104 29158
rect 19076 28966 19196 28994
rect 18892 28614 19104 28642
rect 18788 28552 18840 28558
rect 18788 28494 18840 28500
rect 18972 28552 19024 28558
rect 18972 28494 19024 28500
rect 18880 28416 18932 28422
rect 18786 28384 18842 28393
rect 18880 28358 18932 28364
rect 18786 28319 18842 28328
rect 18604 27396 18656 27402
rect 18604 27338 18656 27344
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18524 27062 18552 27270
rect 18616 27130 18644 27338
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18602 27024 18658 27033
rect 18708 26994 18736 27338
rect 18602 26959 18604 26968
rect 18656 26959 18658 26968
rect 18696 26988 18748 26994
rect 18604 26930 18656 26936
rect 18696 26930 18748 26936
rect 18510 26480 18566 26489
rect 18510 26415 18512 26424
rect 18564 26415 18566 26424
rect 18512 26386 18564 26392
rect 18616 26382 18644 26930
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18432 26030 18736 26058
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 18432 25498 18460 25842
rect 18420 25492 18472 25498
rect 18420 25434 18472 25440
rect 18604 25220 18656 25226
rect 18604 25162 18656 25168
rect 18616 24886 18644 25162
rect 18512 24880 18564 24886
rect 18512 24822 18564 24828
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18420 24676 18472 24682
rect 18420 24618 18472 24624
rect 18432 22760 18460 24618
rect 18524 22930 18552 24822
rect 18616 23050 18644 24822
rect 18708 23730 18736 26030
rect 18800 25838 18828 28319
rect 18892 25906 18920 28358
rect 18984 27946 19012 28494
rect 18972 27940 19024 27946
rect 18972 27882 19024 27888
rect 18984 27713 19012 27882
rect 18970 27704 19026 27713
rect 18970 27639 19026 27648
rect 18972 27532 19024 27538
rect 18972 27474 19024 27480
rect 18984 27062 19012 27474
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18788 25832 18840 25838
rect 18788 25774 18840 25780
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18892 25430 18920 25638
rect 18880 25424 18932 25430
rect 18880 25366 18932 25372
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 18880 25288 18932 25294
rect 18984 25276 19012 25366
rect 18932 25248 19012 25276
rect 18880 25230 18932 25236
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18892 24800 18920 25230
rect 18972 24812 19024 24818
rect 18892 24772 18972 24800
rect 18800 24682 18828 24754
rect 18788 24676 18840 24682
rect 18788 24618 18840 24624
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 18708 23118 18736 23666
rect 18696 23112 18748 23118
rect 18800 23089 18828 24142
rect 18892 23186 18920 24772
rect 18972 24754 19024 24760
rect 18972 24200 19024 24206
rect 18972 24142 19024 24148
rect 18984 23662 19012 24142
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18972 23520 19024 23526
rect 18972 23462 19024 23468
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18984 23089 19012 23462
rect 19076 23225 19104 28614
rect 19168 28218 19196 28966
rect 19260 28762 19288 30194
rect 19352 30190 19380 30670
rect 19340 30184 19392 30190
rect 19340 30126 19392 30132
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19246 28248 19302 28257
rect 19156 28212 19208 28218
rect 19246 28183 19248 28192
rect 19156 28154 19208 28160
rect 19300 28183 19302 28192
rect 19248 28154 19300 28160
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19168 24410 19196 28018
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 19260 24177 19288 26250
rect 19246 24168 19302 24177
rect 19246 24103 19302 24112
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19168 23594 19196 24006
rect 19260 23798 19288 24006
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19352 23730 19380 29990
rect 19430 28792 19486 28801
rect 19430 28727 19486 28736
rect 19444 28014 19472 28727
rect 19536 28014 19564 32524
rect 19800 32506 19852 32512
rect 19892 32564 19944 32570
rect 19892 32506 19944 32512
rect 19812 31822 19840 32506
rect 19904 32473 19932 32506
rect 19890 32464 19946 32473
rect 19996 32434 20024 32710
rect 19890 32399 19946 32408
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19892 32292 19944 32298
rect 19892 32234 19944 32240
rect 19708 31816 19760 31822
rect 19708 31758 19760 31764
rect 19800 31816 19852 31822
rect 19800 31758 19852 31764
rect 19614 30560 19670 30569
rect 19614 30495 19670 30504
rect 19628 30394 19656 30495
rect 19616 30388 19668 30394
rect 19616 30330 19668 30336
rect 19628 30054 19656 30330
rect 19616 30048 19668 30054
rect 19616 29990 19668 29996
rect 19720 29782 19748 31758
rect 19800 30728 19852 30734
rect 19800 30670 19852 30676
rect 19708 29776 19760 29782
rect 19708 29718 19760 29724
rect 19708 29640 19760 29646
rect 19708 29582 19760 29588
rect 19616 29572 19668 29578
rect 19616 29514 19668 29520
rect 19628 29481 19656 29514
rect 19614 29472 19670 29481
rect 19614 29407 19670 29416
rect 19432 28008 19484 28014
rect 19432 27950 19484 27956
rect 19524 28008 19576 28014
rect 19524 27950 19576 27956
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19444 26246 19472 27406
rect 19536 26790 19564 27950
rect 19616 27940 19668 27946
rect 19616 27882 19668 27888
rect 19628 27470 19656 27882
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19616 26240 19668 26246
rect 19616 26182 19668 26188
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 19444 24614 19472 25978
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19536 24290 19564 25774
rect 19628 25702 19656 26182
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19444 24262 19564 24290
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19260 23304 19288 23598
rect 19168 23276 19288 23304
rect 19338 23352 19394 23361
rect 19444 23338 19472 24262
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19394 23310 19472 23338
rect 19338 23287 19340 23296
rect 19062 23216 19118 23225
rect 19062 23151 19118 23160
rect 18696 23054 18748 23060
rect 18786 23080 18842 23089
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18524 22902 18644 22930
rect 18432 22732 18552 22760
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18236 22500 18288 22506
rect 18236 22442 18288 22448
rect 18248 21554 18276 22442
rect 18432 22030 18460 22578
rect 18524 22137 18552 22732
rect 18616 22574 18644 22902
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18510 22128 18566 22137
rect 18510 22063 18566 22072
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18248 20874 18276 21490
rect 18524 21146 18552 21490
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 18156 20454 18276 20482
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18156 19922 18184 20266
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18248 19258 18276 20454
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18326 20360 18382 20369
rect 18326 20295 18382 20304
rect 18340 19854 18368 20295
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18432 19514 18460 20402
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18156 19230 18276 19258
rect 18156 18873 18184 19230
rect 18234 19136 18290 19145
rect 18234 19071 18290 19080
rect 18142 18864 18198 18873
rect 18142 18799 18198 18808
rect 18248 18766 18276 19071
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 17960 17604 18012 17610
rect 17960 17546 18012 17552
rect 17972 17270 18000 17546
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17696 14414 17724 15098
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17130 12271 17186 12280
rect 17224 12300 17276 12306
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 17144 9160 17172 12271
rect 17224 12242 17276 12248
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17236 11286 17264 11698
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17222 11112 17278 11121
rect 17222 11047 17224 11056
rect 17276 11047 17278 11056
rect 17224 11018 17276 11024
rect 17052 9132 17172 9160
rect 17052 8974 17080 9132
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16868 8588 16988 8616
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14556 2848 14608 2854
rect 14752 2836 14780 3538
rect 15396 3534 15424 4014
rect 15764 3942 15792 4626
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15856 4185 15884 4558
rect 15842 4176 15898 4185
rect 15842 4111 15844 4120
rect 15896 4111 15898 4120
rect 15844 4082 15896 4088
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15120 3126 15148 3334
rect 15672 3126 15700 3878
rect 15856 3602 15884 4082
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15948 3058 15976 4694
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16040 4282 16068 4558
rect 16868 4554 16896 8588
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16960 7818 16988 8434
rect 17052 8430 17080 8910
rect 17144 8498 17172 8978
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 17052 7954 17080 8366
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16960 6390 16988 7754
rect 16948 6384 17000 6390
rect 16948 6326 17000 6332
rect 17052 4690 17080 7890
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17144 6866 17172 7346
rect 17236 7342 17264 11018
rect 17328 8498 17356 13874
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17604 13462 17632 13806
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17420 12714 17448 13262
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17512 12782 17540 13194
rect 17604 12889 17632 13262
rect 17590 12880 17646 12889
rect 17590 12815 17646 12824
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17408 12708 17460 12714
rect 17408 12650 17460 12656
rect 17512 12442 17540 12718
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17696 12345 17724 14010
rect 17880 14006 17908 15302
rect 17972 15042 18000 17206
rect 18052 17128 18104 17134
rect 18050 17096 18052 17105
rect 18104 17096 18106 17105
rect 18050 17031 18106 17040
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 18064 15162 18092 16458
rect 18156 15178 18184 18702
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18052 15156 18104 15162
rect 18156 15150 18276 15178
rect 18052 15098 18104 15104
rect 17972 15014 18184 15042
rect 17972 14414 18000 15014
rect 18156 14958 18184 15014
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17972 13394 18000 14350
rect 18064 14278 18092 14894
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18248 13734 18276 15150
rect 18340 14958 18368 16526
rect 18432 15570 18460 19450
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 17960 13388 18012 13394
rect 18012 13348 18092 13376
rect 17960 13330 18012 13336
rect 17776 12368 17828 12374
rect 17682 12336 17738 12345
rect 17776 12310 17828 12316
rect 17682 12271 17738 12280
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 10554 17448 12038
rect 17788 11914 17816 12310
rect 18064 12238 18092 13348
rect 18248 12442 18276 13670
rect 18340 13326 18368 13670
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18326 12336 18382 12345
rect 18248 12280 18326 12288
rect 18248 12260 18328 12280
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 17788 11886 17908 11914
rect 17498 11792 17554 11801
rect 17880 11762 17908 11886
rect 17498 11727 17554 11736
rect 17592 11756 17644 11762
rect 17512 11694 17540 11727
rect 17592 11698 17644 11704
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17604 11529 17632 11698
rect 17590 11520 17646 11529
rect 17590 11455 17646 11464
rect 17696 11393 17724 11698
rect 17972 11642 18000 11698
rect 17880 11626 18000 11642
rect 17868 11620 18012 11626
rect 17920 11614 17960 11620
rect 17868 11562 17920 11568
rect 17960 11562 18012 11568
rect 17682 11384 17738 11393
rect 17682 11319 17738 11328
rect 18156 11286 18184 12174
rect 17684 11280 17736 11286
rect 17498 11248 17554 11257
rect 17684 11222 17736 11228
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 17498 11183 17554 11192
rect 17512 11150 17540 11183
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17696 10606 17724 11222
rect 18248 11098 18276 12260
rect 18380 12271 18382 12280
rect 18328 12242 18380 12248
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 17880 11070 18276 11098
rect 17774 10704 17830 10713
rect 17774 10639 17776 10648
rect 17828 10639 17830 10648
rect 17776 10610 17828 10616
rect 17684 10600 17736 10606
rect 17420 10526 17540 10554
rect 17684 10542 17736 10548
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 10169 17448 10406
rect 17406 10160 17462 10169
rect 17406 10095 17462 10104
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17420 8498 17448 9862
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17328 7478 17356 7890
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17236 7002 17264 7278
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17144 6254 17172 6802
rect 17236 6730 17264 6938
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17328 6458 17356 6802
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17420 5642 17448 6394
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17512 5386 17540 10526
rect 17696 9586 17724 10542
rect 17880 10470 17908 11070
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 17958 10704 18014 10713
rect 18064 10674 18092 10950
rect 17958 10639 17960 10648
rect 18012 10639 18014 10648
rect 18052 10668 18104 10674
rect 17960 10610 18012 10616
rect 18052 10610 18104 10616
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17590 9208 17646 9217
rect 17590 9143 17646 9152
rect 17604 9110 17632 9143
rect 17788 9110 17816 9998
rect 18064 9926 18092 10610
rect 18248 10062 18276 10950
rect 18340 10470 18368 12038
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 17868 9920 17920 9926
rect 18052 9920 18104 9926
rect 17868 9862 17920 9868
rect 17972 9880 18052 9908
rect 17880 9654 17908 9862
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17592 9104 17644 9110
rect 17592 9046 17644 9052
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17788 8974 17816 9046
rect 17880 8974 17908 9590
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17420 5358 17540 5386
rect 17420 4826 17448 5358
rect 17498 5264 17554 5273
rect 17498 5199 17554 5208
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 17420 4554 17448 4762
rect 17512 4758 17540 5199
rect 17500 4752 17552 4758
rect 17500 4694 17552 4700
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 16132 4146 16160 4490
rect 16212 4480 16264 4486
rect 16264 4440 16344 4468
rect 16212 4422 16264 4428
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16224 3942 16252 4082
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16040 3194 16068 3538
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 14608 2808 14780 2836
rect 14556 2790 14608 2796
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 800 14228 2246
rect 14844 800 14872 2586
rect 15200 2372 15252 2378
rect 15396 2366 15608 2394
rect 15396 2360 15424 2366
rect 15252 2332 15424 2360
rect 15200 2314 15252 2320
rect 15580 2310 15608 2366
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15488 800 15516 2246
rect 16132 800 16160 3674
rect 16224 3058 16252 3878
rect 16316 3058 16344 4440
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 16408 3194 16436 4014
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16394 3088 16450 3097
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16304 3052 16356 3058
rect 16394 3023 16396 3032
rect 16304 2994 16356 3000
rect 16448 3023 16450 3032
rect 16396 2994 16448 3000
rect 16500 2922 16528 4014
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16316 2394 16344 2518
rect 16684 2514 16712 3062
rect 17144 2922 17172 4014
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17328 3602 17356 3878
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16316 2366 16528 2394
rect 17420 2378 17448 3878
rect 17604 3670 17632 8434
rect 17880 8378 17908 8910
rect 17972 8498 18000 9880
rect 18052 9862 18104 9868
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 9382 18092 9454
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 8974 18092 9318
rect 18156 8974 18184 9522
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18234 8936 18290 8945
rect 18156 8650 18184 8910
rect 18234 8871 18236 8880
rect 18288 8871 18290 8880
rect 18236 8842 18288 8848
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18156 8622 18276 8650
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17880 8350 18000 8378
rect 17972 8242 18000 8350
rect 17972 8214 18092 8242
rect 18064 7478 18092 8214
rect 18156 7546 18184 8502
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17880 6866 17908 6938
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 18064 6730 18092 7414
rect 18248 7410 18276 8622
rect 18340 8566 18368 8774
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 18236 7404 18288 7410
rect 18288 7364 18368 7392
rect 18236 7346 18288 7352
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 17682 6488 17738 6497
rect 17682 6423 17684 6432
rect 17736 6423 17738 6432
rect 17684 6394 17736 6400
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17880 6066 17908 6258
rect 17880 6038 18000 6066
rect 17972 5642 18000 6038
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17972 4622 18000 5578
rect 18064 5574 18092 6666
rect 18248 6254 18276 6666
rect 18340 6458 18368 7364
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18236 4752 18288 4758
rect 18236 4694 18288 4700
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 4078 17724 4422
rect 18064 4146 18092 4490
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17512 2990 17540 3334
rect 17604 3126 17632 3470
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17696 2854 17724 4014
rect 18248 3602 18276 4694
rect 18432 4622 18460 14554
rect 18524 11558 18552 19790
rect 18708 19718 18736 23054
rect 18786 23015 18842 23024
rect 18970 23080 19026 23089
rect 18970 23015 19026 23024
rect 19168 22953 19196 23276
rect 19392 23287 19394 23296
rect 19340 23258 19392 23264
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19154 22944 19210 22953
rect 19154 22879 19210 22888
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18616 19446 18644 19654
rect 18800 19514 18828 21830
rect 19168 21672 19196 22879
rect 19076 21644 19196 21672
rect 19076 19922 19104 21644
rect 19260 21554 19288 23122
rect 19352 22710 19380 23122
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19338 21992 19394 22001
rect 19338 21927 19340 21936
rect 19392 21927 19394 21936
rect 19340 21898 19392 21904
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19168 21146 19196 21490
rect 19260 21457 19288 21490
rect 19246 21448 19302 21457
rect 19246 21383 19302 21392
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19352 20618 19380 21286
rect 19260 20590 19380 20618
rect 19260 20369 19288 20590
rect 19246 20360 19302 20369
rect 19246 20295 19302 20304
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19246 19816 19302 19825
rect 18972 19780 19024 19786
rect 19246 19751 19248 19760
rect 18972 19722 19024 19728
rect 19300 19751 19302 19760
rect 19248 19722 19300 19728
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18616 18698 18644 19246
rect 18604 18692 18656 18698
rect 18604 18634 18656 18640
rect 18602 18320 18658 18329
rect 18602 18255 18658 18264
rect 18616 17882 18644 18255
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18708 15638 18736 15982
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18616 12209 18644 14962
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18708 14278 18736 14418
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18602 12200 18658 12209
rect 18602 12135 18658 12144
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18524 10742 18552 10950
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 9761 18552 10406
rect 18616 10282 18644 12038
rect 18708 10606 18736 14214
rect 18800 10742 18828 19450
rect 18984 19378 19012 19722
rect 19352 19514 19380 20266
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 18892 16726 18920 17818
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18892 13297 18920 16662
rect 18984 15042 19012 17614
rect 19076 15910 19104 19314
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 15162 19104 15438
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 18984 15014 19104 15042
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18878 13288 18934 13297
rect 18878 13223 18934 13232
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18788 10736 18840 10742
rect 18788 10678 18840 10684
rect 18696 10600 18748 10606
rect 18694 10568 18696 10577
rect 18748 10568 18750 10577
rect 18694 10503 18750 10512
rect 18616 10254 18736 10282
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18510 9752 18566 9761
rect 18510 9687 18566 9696
rect 18524 8838 18552 9687
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18512 8560 18564 8566
rect 18616 8548 18644 10134
rect 18564 8520 18644 8548
rect 18512 8502 18564 8508
rect 18708 7818 18736 10254
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18800 8634 18828 8910
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18616 6866 18644 7482
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18512 6792 18564 6798
rect 18510 6760 18512 6769
rect 18564 6760 18566 6769
rect 18510 6695 18566 6704
rect 18708 6662 18736 7754
rect 18892 7546 18920 13126
rect 18984 12442 19012 14826
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 19076 12238 19104 15014
rect 19168 13938 19196 15914
rect 19260 15201 19288 19178
rect 19352 17134 19380 19246
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16658 19380 16934
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19246 15192 19302 15201
rect 19246 15127 19302 15136
rect 19352 15026 19380 16186
rect 19444 15502 19472 22578
rect 19536 21690 19564 24142
rect 19628 23905 19656 24754
rect 19614 23896 19670 23905
rect 19614 23831 19670 23840
rect 19616 23792 19668 23798
rect 19616 23734 19668 23740
rect 19628 23118 19656 23734
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19628 22658 19656 23054
rect 19720 22778 19748 29582
rect 19812 25498 19840 30670
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19800 24404 19852 24410
rect 19800 24346 19852 24352
rect 19812 24138 19840 24346
rect 19904 24274 19932 32234
rect 19984 32020 20036 32026
rect 19984 31962 20036 31968
rect 19996 31822 20024 31962
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 20088 30054 20116 32846
rect 20258 32807 20314 32816
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20444 32224 20496 32230
rect 20444 32166 20496 32172
rect 20456 31754 20484 32166
rect 20536 31884 20588 31890
rect 20536 31826 20588 31832
rect 20364 31726 20484 31754
rect 20168 31680 20220 31686
rect 20168 31622 20220 31628
rect 20180 31346 20208 31622
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20260 31340 20312 31346
rect 20260 31282 20312 31288
rect 20180 30802 20208 31282
rect 20168 30796 20220 30802
rect 20168 30738 20220 30744
rect 20272 30734 20300 31282
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20168 29776 20220 29782
rect 20168 29718 20220 29724
rect 20180 29034 20208 29718
rect 20260 29232 20312 29238
rect 20260 29174 20312 29180
rect 20168 29028 20220 29034
rect 20168 28970 20220 28976
rect 20180 28490 20208 28970
rect 20272 28558 20300 29174
rect 20260 28552 20312 28558
rect 20260 28494 20312 28500
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 19984 27940 20036 27946
rect 19984 27882 20036 27888
rect 19996 27713 20024 27882
rect 19982 27704 20038 27713
rect 19982 27639 20038 27648
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19996 26790 20024 27406
rect 20364 26858 20392 31726
rect 20444 31340 20496 31346
rect 20444 31282 20496 31288
rect 20352 26852 20404 26858
rect 20352 26794 20404 26800
rect 19984 26784 20036 26790
rect 19984 26726 20036 26732
rect 19996 26314 20024 26726
rect 20260 26512 20312 26518
rect 20258 26480 20260 26489
rect 20312 26480 20314 26489
rect 20258 26415 20314 26424
rect 20364 26382 20392 26794
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 19984 25968 20036 25974
rect 19984 25910 20036 25916
rect 20168 25968 20220 25974
rect 20168 25910 20220 25916
rect 19996 25838 20024 25910
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19984 25696 20036 25702
rect 19984 25638 20036 25644
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19800 24132 19852 24138
rect 19800 24074 19852 24080
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19904 23798 19932 24006
rect 19892 23792 19944 23798
rect 19892 23734 19944 23740
rect 19904 23497 19932 23734
rect 19890 23488 19946 23497
rect 19890 23423 19946 23432
rect 19996 23304 20024 25638
rect 20076 25424 20128 25430
rect 20076 25366 20128 25372
rect 19812 23276 20024 23304
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19628 22630 19748 22658
rect 19614 22128 19670 22137
rect 19614 22063 19670 22072
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 19524 21004 19576 21010
rect 19524 20946 19576 20952
rect 19536 15706 19564 20946
rect 19628 20874 19656 22063
rect 19720 21554 19748 22630
rect 19812 22030 19840 23276
rect 19982 23216 20038 23225
rect 19982 23151 20038 23160
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19904 22166 19932 22374
rect 19892 22160 19944 22166
rect 19892 22102 19944 22108
rect 19800 22024 19852 22030
rect 19800 21966 19852 21972
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19616 20868 19668 20874
rect 19616 20810 19668 20816
rect 19628 16250 19656 20810
rect 19720 19786 19748 21082
rect 19708 19780 19760 19786
rect 19708 19722 19760 19728
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19720 18329 19748 19314
rect 19706 18320 19762 18329
rect 19706 18255 19762 18264
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19812 15706 19840 21966
rect 19904 21078 19932 21966
rect 19892 21072 19944 21078
rect 19892 21014 19944 21020
rect 19996 21010 20024 23151
rect 20088 21486 20116 25366
rect 20180 25226 20208 25910
rect 20168 25220 20220 25226
rect 20168 25162 20220 25168
rect 20180 21894 20208 25162
rect 20272 24698 20300 26250
rect 20456 26042 20484 31282
rect 20548 31142 20576 31826
rect 20732 31346 20760 32778
rect 20904 32020 20956 32026
rect 20904 31962 20956 31968
rect 20916 31346 20944 31962
rect 21100 31482 21128 35566
rect 21376 35329 21404 35634
rect 21362 35320 21418 35329
rect 21362 35255 21418 35264
rect 21560 35018 21588 35974
rect 21640 35556 21692 35562
rect 21640 35498 21692 35504
rect 21652 35290 21680 35498
rect 21640 35284 21692 35290
rect 21640 35226 21692 35232
rect 21548 35012 21600 35018
rect 21548 34954 21600 34960
rect 21652 34678 21680 35226
rect 22112 34746 22140 36042
rect 22204 35630 22232 36178
rect 22296 36174 22324 37198
rect 22480 36786 22508 37198
rect 22572 36922 22600 38926
rect 22560 36916 22612 36922
rect 22560 36858 22612 36864
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 22572 36224 22600 36858
rect 23216 36582 23244 38926
rect 23860 37346 23888 38926
rect 23768 37318 23888 37346
rect 23768 37126 23796 37318
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 23756 37120 23808 37126
rect 23756 37062 23808 37068
rect 23296 36848 23348 36854
rect 23296 36790 23348 36796
rect 23308 36666 23336 36790
rect 23860 36786 23888 37198
rect 23848 36780 23900 36786
rect 23848 36722 23900 36728
rect 23480 36712 23532 36718
rect 23308 36660 23480 36666
rect 23308 36654 23532 36660
rect 23308 36638 23520 36654
rect 23204 36576 23256 36582
rect 23204 36518 23256 36524
rect 22744 36236 22796 36242
rect 22572 36196 22744 36224
rect 22744 36178 22796 36184
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22572 36106 22784 36122
rect 22572 36100 22796 36106
rect 22572 36094 22744 36100
rect 22572 35834 22600 36094
rect 22744 36042 22796 36048
rect 23308 36038 23336 36638
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 23400 36038 23428 36518
rect 23478 36272 23534 36281
rect 23534 36216 23704 36224
rect 23478 36207 23480 36216
rect 23532 36196 23704 36216
rect 23480 36178 23532 36184
rect 22652 36032 22704 36038
rect 22652 35974 22704 35980
rect 23296 36032 23348 36038
rect 23296 35974 23348 35980
rect 23388 36032 23440 36038
rect 23388 35974 23440 35980
rect 22560 35828 22612 35834
rect 22560 35770 22612 35776
rect 22664 35630 22692 35974
rect 22192 35624 22244 35630
rect 22192 35566 22244 35572
rect 22284 35624 22336 35630
rect 22284 35566 22336 35572
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 23020 35624 23072 35630
rect 23020 35566 23072 35572
rect 22296 35154 22324 35566
rect 22284 35148 22336 35154
rect 22284 35090 22336 35096
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 21640 34672 21692 34678
rect 21640 34614 21692 34620
rect 22296 34542 22324 35090
rect 23032 35086 23060 35566
rect 23020 35080 23072 35086
rect 23020 35022 23072 35028
rect 22560 35012 22612 35018
rect 22560 34954 22612 34960
rect 22572 34746 22600 34954
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 23572 34740 23624 34746
rect 23572 34682 23624 34688
rect 22284 34536 22336 34542
rect 22284 34478 22336 34484
rect 22296 33998 22324 34478
rect 21640 33992 21692 33998
rect 22008 33992 22060 33998
rect 21640 33934 21692 33940
rect 22006 33960 22008 33969
rect 22284 33992 22336 33998
rect 22060 33960 22062 33969
rect 21652 32570 21680 33934
rect 22284 33934 22336 33940
rect 22006 33895 22062 33904
rect 22008 33856 22060 33862
rect 22296 33844 22324 33934
rect 22008 33798 22060 33804
rect 22112 33816 22324 33844
rect 22376 33856 22428 33862
rect 21824 33652 21876 33658
rect 21824 33594 21876 33600
rect 21836 32910 21864 33594
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21916 32836 21968 32842
rect 21916 32778 21968 32784
rect 21732 32768 21784 32774
rect 21732 32710 21784 32716
rect 21744 32570 21772 32710
rect 21822 32600 21878 32609
rect 21640 32564 21692 32570
rect 21640 32506 21692 32512
rect 21732 32564 21784 32570
rect 21822 32535 21878 32544
rect 21732 32506 21784 32512
rect 21272 32496 21324 32502
rect 21272 32438 21324 32444
rect 21284 32026 21312 32438
rect 21836 32434 21864 32535
rect 21928 32434 21956 32778
rect 22020 32570 22048 33798
rect 22112 33114 22140 33816
rect 22376 33798 22428 33804
rect 22284 33312 22336 33318
rect 22284 33254 22336 33260
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 22008 32564 22060 32570
rect 22008 32506 22060 32512
rect 22296 32473 22324 33254
rect 22388 32978 22416 33798
rect 22572 33590 22600 34682
rect 22836 34536 22888 34542
rect 22836 34478 22888 34484
rect 22848 34202 22876 34478
rect 22836 34196 22888 34202
rect 22836 34138 22888 34144
rect 22652 34128 22704 34134
rect 22652 34070 22704 34076
rect 22560 33584 22612 33590
rect 22560 33526 22612 33532
rect 22468 33108 22520 33114
rect 22468 33050 22520 33056
rect 22376 32972 22428 32978
rect 22376 32914 22428 32920
rect 22480 32609 22508 33050
rect 22466 32600 22522 32609
rect 22466 32535 22522 32544
rect 22560 32496 22612 32502
rect 22098 32464 22154 32473
rect 21640 32428 21692 32434
rect 21640 32370 21692 32376
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 21916 32428 21968 32434
rect 22098 32399 22154 32408
rect 22282 32464 22338 32473
rect 22664 32484 22692 34070
rect 23204 33992 23256 33998
rect 23110 33960 23166 33969
rect 23204 33934 23256 33940
rect 23110 33895 23166 33904
rect 23020 33652 23072 33658
rect 23020 33594 23072 33600
rect 22744 33448 22796 33454
rect 22744 33390 22796 33396
rect 22756 32570 22784 33390
rect 22744 32564 22796 32570
rect 22744 32506 22796 32512
rect 22928 32564 22980 32570
rect 22928 32506 22980 32512
rect 22612 32456 22692 32484
rect 22560 32438 22612 32444
rect 22282 32399 22338 32408
rect 21916 32370 21968 32376
rect 21652 32337 21680 32370
rect 21638 32328 21694 32337
rect 21638 32263 21694 32272
rect 21272 32020 21324 32026
rect 21272 31962 21324 31968
rect 21364 31952 21416 31958
rect 21364 31894 21416 31900
rect 21272 31748 21324 31754
rect 21272 31690 21324 31696
rect 21088 31476 21140 31482
rect 21088 31418 21140 31424
rect 21180 31476 21232 31482
rect 21180 31418 21232 31424
rect 21192 31362 21220 31418
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20904 31340 20956 31346
rect 20904 31282 20956 31288
rect 21008 31334 21220 31362
rect 21284 31346 21312 31690
rect 21272 31340 21324 31346
rect 20628 31272 20680 31278
rect 20628 31214 20680 31220
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20640 30666 20668 31214
rect 20732 31142 20760 31282
rect 20812 31204 20864 31210
rect 20812 31146 20864 31152
rect 20720 31136 20772 31142
rect 20720 31078 20772 31084
rect 20732 30734 20760 31078
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20628 30660 20680 30666
rect 20628 30602 20680 30608
rect 20640 30258 20668 30602
rect 20732 30394 20760 30670
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 20628 30252 20680 30258
rect 20628 30194 20680 30200
rect 20720 30252 20772 30258
rect 20720 30194 20772 30200
rect 20628 29164 20680 29170
rect 20628 29106 20680 29112
rect 20536 28552 20588 28558
rect 20536 28494 20588 28500
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20352 25832 20404 25838
rect 20352 25774 20404 25780
rect 20364 25702 20392 25774
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 20548 25265 20576 28494
rect 20534 25256 20590 25265
rect 20534 25191 20590 25200
rect 20444 25152 20496 25158
rect 20444 25094 20496 25100
rect 20536 25152 20588 25158
rect 20536 25094 20588 25100
rect 20272 24670 20392 24698
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 20272 21962 20300 24550
rect 20364 24070 20392 24670
rect 20352 24064 20404 24070
rect 20352 24006 20404 24012
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20258 21856 20314 21865
rect 20258 21791 20314 21800
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 20088 20890 20116 21422
rect 19904 20862 20116 20890
rect 19904 19514 19932 20862
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19984 19984 20036 19990
rect 19984 19926 20036 19932
rect 19996 19514 20024 19926
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19982 19408 20038 19417
rect 19982 19343 19984 19352
rect 20036 19343 20038 19352
rect 19984 19314 20036 19320
rect 19892 17604 19944 17610
rect 19892 17546 19944 17552
rect 19904 17202 19932 17546
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19996 17082 20024 19314
rect 19904 17066 20024 17082
rect 19892 17060 20024 17066
rect 19944 17054 20024 17060
rect 19892 17002 19944 17008
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19524 15700 19576 15706
rect 19800 15700 19852 15706
rect 19576 15660 19748 15688
rect 19524 15642 19576 15648
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19248 14952 19300 14958
rect 19352 14929 19380 14962
rect 19432 14952 19484 14958
rect 19248 14894 19300 14900
rect 19338 14920 19394 14929
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 13258 19196 13874
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19154 13152 19210 13161
rect 19154 13087 19210 13096
rect 19168 12374 19196 13087
rect 19156 12368 19208 12374
rect 19156 12310 19208 12316
rect 19064 12232 19116 12238
rect 19116 12180 19196 12186
rect 19064 12174 19196 12180
rect 19076 12158 19196 12174
rect 19168 11762 19196 12158
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19260 10690 19288 14894
rect 19432 14894 19484 14900
rect 19338 14855 19394 14864
rect 19444 14550 19472 14894
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19352 13433 19380 13466
rect 19536 13462 19564 15098
rect 19524 13456 19576 13462
rect 19338 13424 19394 13433
rect 19338 13359 19394 13368
rect 19444 13416 19524 13444
rect 19338 13288 19394 13297
rect 19338 13223 19340 13232
rect 19392 13223 19394 13232
rect 19340 13194 19392 13200
rect 19338 13016 19394 13025
rect 19338 12951 19340 12960
rect 19392 12951 19394 12960
rect 19340 12922 19392 12928
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19352 12617 19380 12650
rect 19338 12608 19394 12617
rect 19338 12543 19394 12552
rect 19168 10674 19288 10690
rect 19352 10674 19380 12543
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 19156 10668 19288 10674
rect 19208 10662 19288 10668
rect 19340 10668 19392 10674
rect 19156 10610 19208 10616
rect 19340 10610 19392 10616
rect 18984 9217 19012 10610
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19076 9722 19104 10406
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18970 9208 19026 9217
rect 18970 9143 19026 9152
rect 18984 8974 19012 9143
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 19076 8838 19104 9046
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18972 8424 19024 8430
rect 19076 8401 19104 8434
rect 18972 8366 19024 8372
rect 19062 8392 19118 8401
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18892 6866 18920 7482
rect 18984 7313 19012 8366
rect 19062 8327 19118 8336
rect 19064 7880 19116 7886
rect 19062 7848 19064 7857
rect 19116 7848 19118 7857
rect 19062 7783 19118 7792
rect 19168 7410 19196 10610
rect 19444 9654 19472 13416
rect 19524 13398 19576 13404
rect 19628 11354 19656 15506
rect 19720 13977 19748 15660
rect 19800 15642 19852 15648
rect 19706 13968 19762 13977
rect 19706 13903 19762 13912
rect 19720 13274 19748 13903
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19812 13444 19840 13806
rect 19904 13802 19932 15982
rect 20088 14890 20116 20402
rect 20272 20058 20300 21791
rect 20364 21690 20392 22374
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20364 20534 20392 21490
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20456 20466 20484 25094
rect 20548 24993 20576 25094
rect 20534 24984 20590 24993
rect 20534 24919 20590 24928
rect 20536 24676 20588 24682
rect 20536 24618 20588 24624
rect 20548 24410 20576 24618
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20640 24290 20668 29106
rect 20732 28626 20760 30194
rect 20824 29646 20852 31146
rect 20916 30802 20944 31282
rect 21008 30870 21036 31334
rect 21272 31282 21324 31288
rect 21376 30938 21404 31894
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21364 30932 21416 30938
rect 21284 30892 21364 30920
rect 20996 30864 21048 30870
rect 20996 30806 21048 30812
rect 20904 30796 20956 30802
rect 20904 30738 20956 30744
rect 20916 29646 20944 30738
rect 21284 29782 21312 30892
rect 21364 30874 21416 30880
rect 21364 30592 21416 30598
rect 21362 30560 21364 30569
rect 21416 30560 21418 30569
rect 21362 30495 21418 30504
rect 21272 29776 21324 29782
rect 21272 29718 21324 29724
rect 21284 29646 21312 29718
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20904 29640 20956 29646
rect 20996 29640 21048 29646
rect 20904 29582 20956 29588
rect 20994 29608 20996 29617
rect 21272 29640 21324 29646
rect 21048 29608 21050 29617
rect 21272 29582 21324 29588
rect 20994 29543 21050 29552
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 21008 29170 21036 29446
rect 21270 29336 21326 29345
rect 21270 29271 21326 29280
rect 20812 29164 20864 29170
rect 20996 29164 21048 29170
rect 20864 29124 20944 29152
rect 20812 29106 20864 29112
rect 20720 28620 20772 28626
rect 20720 28562 20772 28568
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20732 26994 20760 27542
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20732 26625 20760 26930
rect 20718 26616 20774 26625
rect 20718 26551 20774 26560
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20732 25294 20760 26250
rect 20824 25922 20852 28358
rect 20916 28150 20944 29124
rect 20996 29106 21048 29112
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21008 28558 21036 29106
rect 21086 28928 21142 28937
rect 21086 28863 21142 28872
rect 21100 28558 21128 28863
rect 21192 28762 21220 29106
rect 21180 28756 21232 28762
rect 21180 28698 21232 28704
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 21088 28552 21140 28558
rect 21088 28494 21140 28500
rect 21284 28234 21312 29271
rect 21376 29034 21404 30495
rect 21652 30326 21680 31758
rect 21732 30932 21784 30938
rect 21732 30874 21784 30880
rect 21744 30734 21772 30874
rect 21732 30728 21784 30734
rect 21732 30670 21784 30676
rect 21836 30546 21864 32370
rect 21928 31890 21956 32370
rect 22112 32026 22140 32399
rect 22296 32042 22324 32399
rect 22100 32020 22152 32026
rect 22020 31980 22100 32008
rect 21916 31884 21968 31890
rect 21916 31826 21968 31832
rect 21916 30864 21968 30870
rect 21916 30806 21968 30812
rect 21744 30518 21864 30546
rect 21640 30320 21692 30326
rect 21640 30262 21692 30268
rect 21548 29776 21600 29782
rect 21548 29718 21600 29724
rect 21456 29572 21508 29578
rect 21456 29514 21508 29520
rect 21468 29170 21496 29514
rect 21560 29209 21588 29718
rect 21744 29646 21772 30518
rect 21824 30388 21876 30394
rect 21824 30330 21876 30336
rect 21732 29640 21784 29646
rect 21732 29582 21784 29588
rect 21640 29504 21692 29510
rect 21744 29481 21772 29582
rect 21640 29446 21692 29452
rect 21730 29472 21786 29481
rect 21652 29306 21680 29446
rect 21730 29407 21786 29416
rect 21836 29306 21864 30330
rect 21640 29300 21692 29306
rect 21640 29242 21692 29248
rect 21824 29300 21876 29306
rect 21824 29242 21876 29248
rect 21546 29200 21602 29209
rect 21456 29164 21508 29170
rect 21652 29170 21680 29242
rect 21546 29135 21602 29144
rect 21640 29164 21692 29170
rect 21456 29106 21508 29112
rect 21640 29106 21692 29112
rect 21364 29028 21416 29034
rect 21364 28970 21416 28976
rect 21362 28656 21418 28665
rect 21362 28591 21418 28600
rect 21376 28558 21404 28591
rect 21364 28552 21416 28558
rect 21364 28494 21416 28500
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21100 28206 21312 28234
rect 20904 28144 20956 28150
rect 20904 28086 20956 28092
rect 20996 27872 21048 27878
rect 20996 27814 21048 27820
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20916 26994 20944 27270
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20824 25894 20944 25922
rect 20812 25764 20864 25770
rect 20812 25706 20864 25712
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20824 24886 20852 25706
rect 20812 24880 20864 24886
rect 20812 24822 20864 24828
rect 20916 24342 20944 25894
rect 21008 24410 21036 27814
rect 21100 27112 21128 28206
rect 21180 28144 21232 28150
rect 21180 28086 21232 28092
rect 21192 27538 21220 28086
rect 21180 27532 21232 27538
rect 21180 27474 21232 27480
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21100 27084 21220 27112
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 21100 26586 21128 26930
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21192 26217 21220 27084
rect 21178 26208 21234 26217
rect 21178 26143 21234 26152
rect 21180 25832 21232 25838
rect 21180 25774 21232 25780
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 20548 24262 20668 24290
rect 20904 24336 20956 24342
rect 20904 24278 20956 24284
rect 20548 24070 20576 24262
rect 20812 24200 20864 24206
rect 20810 24168 20812 24177
rect 20904 24200 20956 24206
rect 20864 24168 20866 24177
rect 20628 24132 20680 24138
rect 20904 24142 20956 24148
rect 20810 24103 20866 24112
rect 20628 24074 20680 24080
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20640 23866 20668 24074
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20536 23316 20588 23322
rect 20536 23258 20588 23264
rect 20548 22642 20576 23258
rect 20640 23186 20668 23666
rect 20732 23526 20760 23666
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20916 22710 20944 24142
rect 21100 24138 21128 25298
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 21008 23322 21036 23598
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20272 19378 20300 19722
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20168 17060 20220 17066
rect 20168 17002 20220 17008
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 20180 14770 20208 17002
rect 19996 14742 20208 14770
rect 19892 13796 19944 13802
rect 19892 13738 19944 13744
rect 19892 13456 19944 13462
rect 19812 13416 19892 13444
rect 19892 13398 19944 13404
rect 19892 13320 19944 13326
rect 19890 13288 19892 13297
rect 19944 13288 19946 13297
rect 19720 13246 19840 13274
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19720 12850 19748 13126
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19720 12628 19748 12786
rect 19812 12696 19840 13246
rect 19890 13223 19946 13232
rect 19812 12668 19932 12696
rect 19720 12600 19840 12628
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19720 11898 19748 12106
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19720 11354 19748 11494
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19246 8936 19302 8945
rect 19246 8871 19248 8880
rect 19300 8871 19302 8880
rect 19248 8842 19300 8848
rect 19352 7886 19380 8978
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19260 7410 19288 7754
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 18970 7304 19026 7313
rect 18970 7239 19026 7248
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18878 6760 18934 6769
rect 18878 6695 18880 6704
rect 18932 6695 18934 6704
rect 18880 6666 18932 6672
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 6322 18736 6598
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18984 6118 19012 6258
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 19168 5370 19196 7210
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 5778 19288 6598
rect 19352 6390 19380 7822
rect 19536 7546 19564 10542
rect 19628 10441 19656 11154
rect 19614 10432 19670 10441
rect 19614 10367 19670 10376
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19352 5658 19380 6326
rect 19444 5710 19472 7414
rect 19628 6780 19656 10202
rect 19720 9042 19748 11154
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19812 8634 19840 12600
rect 19904 11898 19932 12668
rect 19996 12458 20024 14742
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20088 12646 20116 14350
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20180 13433 20208 13466
rect 20166 13424 20222 13433
rect 20166 13359 20222 13368
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20180 12850 20208 13262
rect 20272 13138 20300 17614
rect 20352 15428 20404 15434
rect 20352 15370 20404 15376
rect 20364 15094 20392 15370
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20456 14414 20484 19110
rect 20548 17746 20576 22578
rect 21100 22166 21128 23598
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20640 21146 20668 21422
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20732 19904 20760 22102
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20916 20534 20944 21286
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 20810 20360 20866 20369
rect 20810 20295 20866 20304
rect 20824 19922 20852 20295
rect 20916 19922 20944 20470
rect 20640 19876 20760 19904
rect 20812 19916 20864 19922
rect 20640 19446 20668 19876
rect 20812 19858 20864 19864
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20916 19378 20944 19858
rect 21008 19854 21036 21898
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 21100 20874 21128 21558
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 21086 20496 21142 20505
rect 21086 20431 21142 20440
rect 21100 20262 21128 20431
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20916 18970 20944 19314
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20640 16794 20668 18022
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20732 17134 20760 17818
rect 21008 17202 21036 19790
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 21100 17542 21128 18226
rect 21192 18154 21220 25774
rect 21284 20602 21312 27406
rect 21376 26314 21404 28358
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 21560 27130 21588 27338
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21456 26920 21508 26926
rect 21456 26862 21508 26868
rect 21364 26308 21416 26314
rect 21364 26250 21416 26256
rect 21376 25974 21404 26250
rect 21364 25968 21416 25974
rect 21364 25910 21416 25916
rect 21362 25256 21418 25265
rect 21362 25191 21418 25200
rect 21376 24410 21404 25191
rect 21468 25140 21496 26862
rect 21652 26330 21680 29106
rect 21928 28966 21956 30806
rect 22020 30734 22048 31980
rect 22296 32014 22416 32042
rect 22100 31962 22152 31968
rect 22388 31754 22416 32014
rect 22560 31952 22612 31958
rect 22560 31894 22612 31900
rect 22468 31816 22520 31822
rect 22468 31758 22520 31764
rect 22376 31748 22428 31754
rect 22376 31690 22428 31696
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 22006 30288 22062 30297
rect 22006 30223 22008 30232
rect 22060 30223 22062 30232
rect 22008 30194 22060 30200
rect 22112 30138 22140 31350
rect 22388 30190 22416 31690
rect 22480 30258 22508 31758
rect 22572 31657 22600 31894
rect 22558 31648 22614 31657
rect 22558 31583 22614 31592
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22020 30110 22140 30138
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 22284 30116 22336 30122
rect 22020 29714 22048 30110
rect 22284 30058 22336 30064
rect 22100 30048 22152 30054
rect 22100 29990 22152 29996
rect 22112 29782 22140 29990
rect 22296 29782 22324 30058
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 22100 29776 22152 29782
rect 22100 29718 22152 29724
rect 22192 29776 22244 29782
rect 22192 29718 22244 29724
rect 22284 29776 22336 29782
rect 22284 29718 22336 29724
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 21824 28960 21876 28966
rect 21916 28960 21968 28966
rect 21824 28902 21876 28908
rect 21914 28928 21916 28937
rect 21968 28928 21970 28937
rect 21732 28416 21784 28422
rect 21730 28384 21732 28393
rect 21784 28384 21786 28393
rect 21730 28319 21786 28328
rect 21560 26302 21680 26330
rect 21560 25838 21588 26302
rect 21640 26240 21692 26246
rect 21640 26182 21692 26188
rect 21744 26194 21772 28319
rect 21836 28218 21864 28902
rect 21914 28863 21970 28872
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 22020 28098 22048 29650
rect 22204 28422 22232 29718
rect 22284 29096 22336 29102
rect 22284 29038 22336 29044
rect 22296 28762 22324 29038
rect 22284 28756 22336 28762
rect 22284 28698 22336 28704
rect 22480 28626 22508 29990
rect 22572 28694 22600 31078
rect 22664 30122 22692 32456
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22848 30938 22876 32370
rect 22940 32337 22968 32506
rect 22926 32328 22982 32337
rect 22926 32263 22982 32272
rect 23032 31822 23060 33594
rect 23124 32484 23152 33895
rect 23216 33318 23244 33934
rect 23480 33856 23532 33862
rect 23480 33798 23532 33804
rect 23204 33312 23256 33318
rect 23204 33254 23256 33260
rect 23388 32972 23440 32978
rect 23388 32914 23440 32920
rect 23204 32496 23256 32502
rect 23124 32456 23204 32484
rect 23204 32438 23256 32444
rect 23112 32224 23164 32230
rect 23112 32166 23164 32172
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23018 31512 23074 31521
rect 23018 31447 23074 31456
rect 23032 31278 23060 31447
rect 23020 31272 23072 31278
rect 23020 31214 23072 31220
rect 23020 31136 23072 31142
rect 23020 31078 23072 31084
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 23032 30870 23060 31078
rect 23020 30864 23072 30870
rect 23020 30806 23072 30812
rect 22744 30252 22796 30258
rect 22744 30194 22796 30200
rect 22836 30252 22888 30258
rect 22836 30194 22888 30200
rect 22652 30116 22704 30122
rect 22652 30058 22704 30064
rect 22756 29889 22784 30194
rect 22742 29880 22798 29889
rect 22742 29815 22798 29824
rect 22848 29764 22876 30194
rect 22928 30048 22980 30054
rect 22928 29990 22980 29996
rect 22664 29736 22876 29764
rect 22664 29646 22692 29736
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 22664 29306 22692 29582
rect 22652 29300 22704 29306
rect 22652 29242 22704 29248
rect 22744 29300 22796 29306
rect 22744 29242 22796 29248
rect 22560 28688 22612 28694
rect 22560 28630 22612 28636
rect 22664 28626 22692 29242
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22652 28620 22704 28626
rect 22652 28562 22704 28568
rect 22376 28484 22428 28490
rect 22376 28426 22428 28432
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 21836 28070 22048 28098
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 21836 26926 21864 28070
rect 21916 28008 21968 28014
rect 21916 27950 21968 27956
rect 21928 27334 21956 27950
rect 22204 27674 22232 28086
rect 22388 28082 22416 28426
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21824 26920 21876 26926
rect 21824 26862 21876 26868
rect 22192 26920 22244 26926
rect 22192 26862 22244 26868
rect 21836 26314 21864 26862
rect 22008 26852 22060 26858
rect 22008 26794 22060 26800
rect 21914 26344 21970 26353
rect 21824 26308 21876 26314
rect 22020 26314 22048 26794
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 21914 26279 21916 26288
rect 21824 26250 21876 26256
rect 21968 26279 21970 26288
rect 22008 26308 22060 26314
rect 21916 26250 21968 26256
rect 22008 26250 22060 26256
rect 21548 25832 21600 25838
rect 21548 25774 21600 25780
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21560 25294 21588 25434
rect 21652 25362 21680 26182
rect 21744 26166 21956 26194
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21468 25112 21588 25140
rect 21456 24948 21508 24954
rect 21456 24890 21508 24896
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21468 24290 21496 24890
rect 21376 24262 21496 24290
rect 21376 23662 21404 24262
rect 21560 24052 21588 25112
rect 21652 24206 21680 25298
rect 21744 25294 21772 25638
rect 21824 25492 21876 25498
rect 21824 25434 21876 25440
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 21836 24954 21864 25434
rect 21824 24948 21876 24954
rect 21824 24890 21876 24896
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21640 24200 21692 24206
rect 21640 24142 21692 24148
rect 21560 24024 21772 24052
rect 21364 23656 21416 23662
rect 21364 23598 21416 23604
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21652 23322 21680 23462
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21652 23186 21680 23258
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21362 21040 21418 21049
rect 21362 20975 21418 20984
rect 21376 20942 21404 20975
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21284 18834 21312 20538
rect 21364 20528 21416 20534
rect 21364 20470 21416 20476
rect 21376 19854 21404 20470
rect 21468 20466 21496 20878
rect 21560 20534 21588 20878
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21468 20330 21496 20402
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21560 19990 21588 20470
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 18290 21312 18566
rect 21376 18290 21404 19178
rect 21468 18426 21496 19790
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21180 18148 21232 18154
rect 21180 18090 21232 18096
rect 21178 17776 21234 17785
rect 21178 17711 21234 17720
rect 21192 17678 21220 17711
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21100 17134 21128 17478
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20548 15586 20576 15846
rect 20548 15558 20668 15586
rect 20640 15502 20668 15558
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20548 14929 20576 14962
rect 20534 14920 20590 14929
rect 20534 14855 20590 14864
rect 20444 14408 20496 14414
rect 20364 14356 20444 14362
rect 20364 14350 20496 14356
rect 20364 14334 20484 14350
rect 20364 13326 20392 14334
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20548 13394 20576 13806
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20444 13252 20496 13258
rect 20496 13212 20576 13240
rect 20444 13194 20496 13200
rect 20272 13110 20484 13138
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 19996 12430 20208 12458
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 20180 11830 20208 12430
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19904 10606 19932 11698
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10169 19932 10406
rect 19996 10198 20024 11222
rect 20180 11218 20208 11766
rect 20272 11762 20300 12310
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20258 11112 20314 11121
rect 20258 11047 20314 11056
rect 20272 11014 20300 11047
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20074 10704 20130 10713
rect 20074 10639 20130 10648
rect 20088 10266 20116 10639
rect 20364 10554 20392 12582
rect 20180 10526 20392 10554
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19984 10192 20036 10198
rect 19890 10160 19946 10169
rect 19984 10134 20036 10140
rect 19890 10095 19946 10104
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 19720 7478 19748 7754
rect 19708 7472 19760 7478
rect 19708 7414 19760 7420
rect 19904 7206 19932 9454
rect 19892 7200 19944 7206
rect 19996 7188 20024 10134
rect 20074 9616 20130 9625
rect 20074 9551 20130 9560
rect 20088 9042 20116 9551
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20076 7200 20128 7206
rect 19996 7160 20076 7188
rect 19892 7142 19944 7148
rect 20076 7142 20128 7148
rect 19904 7002 19932 7142
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 20088 6934 20116 7142
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 19708 6792 19760 6798
rect 19628 6752 19708 6780
rect 19628 6662 19656 6752
rect 19708 6734 19760 6740
rect 19982 6760 20038 6769
rect 19982 6695 20038 6704
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19628 5710 19656 6394
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19720 5710 19748 6258
rect 19996 5710 20024 6695
rect 19260 5630 19380 5658
rect 19432 5704 19484 5710
rect 19616 5704 19668 5710
rect 19484 5664 19564 5692
rect 19432 5646 19484 5652
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19168 5234 19196 5306
rect 19260 5302 19288 5630
rect 19536 5574 19564 5664
rect 19616 5646 19668 5652
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 18524 4826 18552 5170
rect 19352 5030 19380 5510
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18418 4312 18474 4321
rect 18418 4247 18420 4256
rect 18472 4247 18474 4256
rect 18420 4218 18472 4224
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18616 4049 18644 4082
rect 18602 4040 18658 4049
rect 18602 3975 18604 3984
rect 18656 3975 18658 3984
rect 18604 3946 18656 3952
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18432 3194 18460 3334
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18616 3058 18644 3402
rect 18800 3194 18828 3878
rect 19536 3738 19564 5510
rect 19720 5030 19748 5646
rect 20180 5098 20208 10526
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20272 9042 20300 10406
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20258 8528 20314 8537
rect 20258 8463 20260 8472
rect 20312 8463 20314 8472
rect 20260 8434 20312 8440
rect 20364 8294 20392 8842
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20272 5710 20300 7890
rect 20456 7546 20484 13110
rect 20548 12646 20576 13212
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20548 11762 20576 11834
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20640 11506 20668 15438
rect 20732 14550 20760 17070
rect 21284 16998 21312 18226
rect 21560 18193 21588 18702
rect 21546 18184 21602 18193
rect 21546 18119 21602 18128
rect 21652 17882 21680 21626
rect 21744 18222 21772 24024
rect 21836 20398 21864 24278
rect 21928 24070 21956 26166
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22020 25401 22048 25842
rect 22006 25392 22062 25401
rect 22006 25327 22062 25336
rect 22008 25152 22060 25158
rect 22008 25094 22060 25100
rect 22020 24886 22048 25094
rect 22008 24880 22060 24886
rect 22008 24822 22060 24828
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 22112 23730 22140 26386
rect 22204 26353 22232 26862
rect 22388 26586 22416 28018
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22652 27872 22704 27878
rect 22652 27814 22704 27820
rect 22572 27062 22600 27814
rect 22560 27056 22612 27062
rect 22560 26998 22612 27004
rect 22560 26920 22612 26926
rect 22560 26862 22612 26868
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22190 26344 22246 26353
rect 22190 26279 22246 26288
rect 22572 25906 22600 26862
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22192 25220 22244 25226
rect 22192 25162 22244 25168
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 21928 22098 21956 23054
rect 22112 23050 22140 23530
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22100 23044 22152 23050
rect 22100 22986 22152 22992
rect 22020 22545 22048 22986
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22006 22536 22062 22545
rect 22006 22471 22062 22480
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21928 21146 21956 22034
rect 22112 22030 22140 22578
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 22020 21554 22048 21830
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 21824 20392 21876 20398
rect 21824 20334 21876 20340
rect 22020 20330 22048 21490
rect 22204 21026 22232 25162
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22388 21486 22416 23666
rect 22572 23118 22600 25842
rect 22664 23769 22692 27814
rect 22756 26314 22784 29242
rect 22848 29170 22876 29582
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 22940 29102 22968 29990
rect 23020 29504 23072 29510
rect 23020 29446 23072 29452
rect 22928 29096 22980 29102
rect 22928 29038 22980 29044
rect 22836 28688 22888 28694
rect 22836 28630 22888 28636
rect 22848 28014 22876 28630
rect 23032 28558 23060 29446
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 22926 28112 22982 28121
rect 22926 28047 22928 28056
rect 22980 28047 22982 28056
rect 22928 28018 22980 28024
rect 22836 28008 22888 28014
rect 22836 27950 22888 27956
rect 22848 27849 22876 27950
rect 22928 27940 22980 27946
rect 22928 27882 22980 27888
rect 22834 27840 22890 27849
rect 22834 27775 22890 27784
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22744 26308 22796 26314
rect 22744 26250 22796 26256
rect 22848 25974 22876 27270
rect 22940 26926 22968 27882
rect 22928 26920 22980 26926
rect 22928 26862 22980 26868
rect 22928 26580 22980 26586
rect 22928 26522 22980 26528
rect 22940 26382 22968 26522
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 22836 25968 22888 25974
rect 22836 25910 22888 25916
rect 22848 25498 22876 25910
rect 23032 25838 23060 28494
rect 23124 28082 23152 32166
rect 23216 31346 23244 32438
rect 23400 32434 23428 32914
rect 23492 32570 23520 33798
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23480 32360 23532 32366
rect 23480 32302 23532 32308
rect 23204 31340 23256 31346
rect 23204 31282 23256 31288
rect 23204 31136 23256 31142
rect 23204 31078 23256 31084
rect 23216 30734 23244 31078
rect 23492 30977 23520 32302
rect 23584 31346 23612 34682
rect 23676 34066 23704 36196
rect 23860 35154 23888 36722
rect 24400 36712 24452 36718
rect 24400 36654 24452 36660
rect 24412 36378 24440 36654
rect 24400 36372 24452 36378
rect 24400 36314 24452 36320
rect 24504 35698 24532 38926
rect 25044 36236 25096 36242
rect 25044 36178 25096 36184
rect 23940 35692 23992 35698
rect 23940 35634 23992 35640
rect 24492 35692 24544 35698
rect 24492 35634 24544 35640
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 23848 35148 23900 35154
rect 23848 35090 23900 35096
rect 23848 34740 23900 34746
rect 23848 34682 23900 34688
rect 23860 34474 23888 34682
rect 23952 34610 23980 35634
rect 24124 34672 24176 34678
rect 24124 34614 24176 34620
rect 23940 34604 23992 34610
rect 23940 34546 23992 34552
rect 23848 34468 23900 34474
rect 23848 34410 23900 34416
rect 23664 34060 23716 34066
rect 23664 34002 23716 34008
rect 24136 33998 24164 34614
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 24124 33992 24176 33998
rect 24124 33934 24176 33940
rect 23940 33924 23992 33930
rect 23940 33866 23992 33872
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23676 32978 23704 33254
rect 23664 32972 23716 32978
rect 23664 32914 23716 32920
rect 23846 32872 23902 32881
rect 23846 32807 23902 32816
rect 23664 32768 23716 32774
rect 23664 32710 23716 32716
rect 23676 32609 23704 32710
rect 23662 32600 23718 32609
rect 23662 32535 23718 32544
rect 23676 31754 23704 32535
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23768 31793 23796 32370
rect 23860 32026 23888 32807
rect 23848 32020 23900 32026
rect 23848 31962 23900 31968
rect 23754 31784 23810 31793
rect 23664 31748 23716 31754
rect 23754 31719 23810 31728
rect 23664 31690 23716 31696
rect 23768 31686 23796 31719
rect 23756 31680 23808 31686
rect 23756 31622 23808 31628
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23478 30968 23534 30977
rect 23478 30903 23534 30912
rect 23388 30864 23440 30870
rect 23388 30806 23440 30812
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23204 30592 23256 30598
rect 23204 30534 23256 30540
rect 23216 30326 23244 30534
rect 23204 30320 23256 30326
rect 23256 30280 23336 30308
rect 23204 30262 23256 30268
rect 23204 30048 23256 30054
rect 23204 29990 23256 29996
rect 23216 29034 23244 29990
rect 23308 29646 23336 30280
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23400 29306 23428 30806
rect 23480 30728 23532 30734
rect 23480 30670 23532 30676
rect 23388 29300 23440 29306
rect 23388 29242 23440 29248
rect 23294 29200 23350 29209
rect 23492 29152 23520 30670
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23584 30297 23612 30534
rect 23570 30288 23626 30297
rect 23768 30258 23796 31622
rect 23860 30326 23888 31962
rect 23952 31634 23980 33866
rect 24032 33856 24084 33862
rect 24032 33798 24084 33804
rect 24044 32910 24072 33798
rect 24400 33584 24452 33590
rect 24400 33526 24452 33532
rect 24124 33040 24176 33046
rect 24124 32982 24176 32988
rect 24412 32994 24440 33526
rect 24504 33114 24532 34478
rect 24872 34406 24900 35634
rect 25056 35630 25084 36178
rect 25044 35624 25096 35630
rect 25044 35566 25096 35572
rect 25148 34678 25176 38926
rect 25228 37324 25280 37330
rect 25228 37266 25280 37272
rect 25240 36378 25268 37266
rect 25792 36854 25820 38926
rect 25780 36848 25832 36854
rect 25780 36790 25832 36796
rect 25228 36372 25280 36378
rect 25228 36314 25280 36320
rect 25594 36136 25650 36145
rect 25594 36071 25596 36080
rect 25648 36071 25650 36080
rect 25596 36042 25648 36048
rect 26436 35698 26464 38926
rect 26424 35692 26476 35698
rect 26424 35634 26476 35640
rect 27080 35290 27108 38926
rect 29012 37262 29040 38926
rect 29656 37262 29684 38926
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 29000 37256 29052 37262
rect 29000 37198 29052 37204
rect 29644 37256 29696 37262
rect 29644 37198 29696 37204
rect 29276 37120 29328 37126
rect 29276 37062 29328 37068
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 27068 35284 27120 35290
rect 27068 35226 27120 35232
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 25320 35012 25372 35018
rect 25320 34954 25372 34960
rect 25136 34672 25188 34678
rect 25136 34614 25188 34620
rect 25332 34610 25360 34954
rect 26608 34944 26660 34950
rect 26608 34886 26660 34892
rect 27344 34944 27396 34950
rect 27344 34886 27396 34892
rect 25412 34740 25464 34746
rect 25412 34682 25464 34688
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 24860 34400 24912 34406
rect 24860 34342 24912 34348
rect 24768 34196 24820 34202
rect 24768 34138 24820 34144
rect 24676 33652 24728 33658
rect 24676 33594 24728 33600
rect 24492 33108 24544 33114
rect 24492 33050 24544 33056
rect 24584 33040 24636 33046
rect 24032 32904 24084 32910
rect 24030 32872 24032 32881
rect 24084 32872 24086 32881
rect 24030 32807 24086 32816
rect 24032 32768 24084 32774
rect 24032 32710 24084 32716
rect 24044 32366 24072 32710
rect 24136 32570 24164 32982
rect 24412 32966 24532 32994
rect 24584 32982 24636 32988
rect 24400 32904 24452 32910
rect 24400 32846 24452 32852
rect 24124 32564 24176 32570
rect 24124 32506 24176 32512
rect 24306 32464 24362 32473
rect 24306 32399 24308 32408
rect 24360 32399 24362 32408
rect 24308 32370 24360 32376
rect 24032 32360 24084 32366
rect 24032 32302 24084 32308
rect 24044 31890 24072 32302
rect 24308 32224 24360 32230
rect 24308 32166 24360 32172
rect 24124 31952 24176 31958
rect 24124 31894 24176 31900
rect 24032 31884 24084 31890
rect 24032 31826 24084 31832
rect 24030 31648 24086 31657
rect 23952 31606 24030 31634
rect 24030 31583 24086 31592
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 23848 30320 23900 30326
rect 23848 30262 23900 30268
rect 23570 30223 23626 30232
rect 23756 30252 23808 30258
rect 23756 30194 23808 30200
rect 23768 30161 23796 30194
rect 23952 30190 23980 30670
rect 23940 30184 23992 30190
rect 23754 30152 23810 30161
rect 23940 30126 23992 30132
rect 23754 30087 23810 30096
rect 23952 29850 23980 30126
rect 23940 29844 23992 29850
rect 23940 29786 23992 29792
rect 23664 29572 23716 29578
rect 23664 29514 23716 29520
rect 23350 29144 23520 29152
rect 23294 29135 23296 29144
rect 23348 29124 23520 29144
rect 23296 29106 23348 29112
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 23216 28422 23244 28970
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23308 28098 23336 28970
rect 23388 28960 23440 28966
rect 23388 28902 23440 28908
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 23216 28070 23336 28098
rect 23400 28082 23428 28902
rect 23388 28076 23440 28082
rect 23112 27872 23164 27878
rect 23110 27840 23112 27849
rect 23164 27840 23166 27849
rect 23110 27775 23166 27784
rect 23112 27396 23164 27402
rect 23112 27338 23164 27344
rect 23124 27130 23152 27338
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 23216 26790 23244 28070
rect 23388 28018 23440 28024
rect 23296 28008 23348 28014
rect 23296 27950 23348 27956
rect 23308 27674 23336 27950
rect 23296 27668 23348 27674
rect 23296 27610 23348 27616
rect 23400 27538 23428 28018
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23492 26874 23520 29124
rect 23572 28484 23624 28490
rect 23572 28426 23624 28432
rect 23584 27470 23612 28426
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23400 26846 23520 26874
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 23020 25832 23072 25838
rect 23020 25774 23072 25780
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 23020 25424 23072 25430
rect 23020 25366 23072 25372
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22756 24954 22784 25230
rect 23032 25226 23060 25366
rect 23020 25220 23072 25226
rect 23020 25162 23072 25168
rect 22744 24948 22796 24954
rect 22744 24890 22796 24896
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 22650 23760 22706 23769
rect 22650 23695 22706 23704
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22572 22710 22600 22918
rect 22560 22704 22612 22710
rect 22560 22646 22612 22652
rect 22664 22642 22692 22918
rect 22848 22778 22876 23054
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22480 22234 22508 22374
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22112 20998 22232 21026
rect 22112 20806 22140 20998
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 22204 20602 22232 20810
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21732 18216 21784 18222
rect 21732 18158 21784 18164
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21638 17640 21694 17649
rect 21376 17338 21404 17614
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20812 15088 20864 15094
rect 20810 15056 20812 15065
rect 20864 15056 20866 15065
rect 20810 14991 20866 15000
rect 21008 14958 21036 16730
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 21008 14414 21036 14894
rect 20720 14408 20772 14414
rect 20718 14376 20720 14385
rect 20812 14408 20864 14414
rect 20772 14376 20774 14385
rect 20812 14350 20864 14356
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20718 14311 20774 14320
rect 20824 13190 20852 14350
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20548 11478 20668 11506
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20548 11150 20576 11478
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20640 10742 20668 11018
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20732 10674 20760 11494
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20824 10554 20852 12038
rect 20916 10713 20944 14282
rect 21100 13410 21128 14350
rect 21008 13382 21128 13410
rect 21008 10742 21036 13382
rect 21192 12617 21220 15302
rect 21284 14929 21312 15370
rect 21376 15065 21404 15642
rect 21468 15162 21496 17614
rect 21638 17575 21694 17584
rect 21652 16522 21680 17575
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21744 16266 21772 18158
rect 21836 17898 21864 18906
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 21928 18057 21956 18702
rect 22020 18358 22048 18770
rect 22112 18766 22140 19994
rect 22100 18760 22152 18766
rect 22152 18720 22232 18748
rect 22100 18702 22152 18708
rect 22008 18352 22060 18358
rect 22008 18294 22060 18300
rect 22008 18080 22060 18086
rect 21914 18048 21970 18057
rect 22008 18022 22060 18028
rect 21914 17983 21970 17992
rect 21836 17870 21956 17898
rect 21824 17808 21876 17814
rect 21824 17750 21876 17756
rect 21836 17542 21864 17750
rect 21928 17626 21956 17870
rect 22020 17746 22048 18022
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 21928 17610 22140 17626
rect 21928 17604 22152 17610
rect 21928 17598 22100 17604
rect 22100 17546 22152 17552
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 21560 16238 21772 16266
rect 21560 16046 21588 16238
rect 21640 16176 21692 16182
rect 21638 16144 21640 16153
rect 21692 16144 21694 16153
rect 21638 16079 21694 16088
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 21560 15570 21588 15982
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21362 15056 21418 15065
rect 21362 14991 21418 15000
rect 21270 14920 21326 14929
rect 21270 14855 21326 14864
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21376 14074 21404 14826
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21560 14074 21588 14758
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21652 13938 21680 14486
rect 21836 14006 21864 17478
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 21928 16833 21956 17206
rect 22020 17184 22048 17478
rect 22100 17196 22152 17202
rect 22020 17156 22100 17184
rect 22100 17138 22152 17144
rect 21914 16824 21970 16833
rect 21914 16759 21970 16768
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21928 15638 21956 16050
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 22020 14929 22048 16662
rect 22204 16590 22232 18720
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22296 16436 22324 20742
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22388 17882 22416 20402
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22480 17762 22508 21830
rect 22652 21412 22704 21418
rect 22652 21354 22704 21360
rect 22664 19922 22692 21354
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22558 19680 22614 19689
rect 22558 19615 22614 19624
rect 22572 19514 22600 19615
rect 22650 19544 22706 19553
rect 22560 19508 22612 19514
rect 22650 19479 22706 19488
rect 22560 19450 22612 19456
rect 22558 19408 22614 19417
rect 22664 19378 22692 19479
rect 22558 19343 22614 19352
rect 22652 19372 22704 19378
rect 22112 16408 22324 16436
rect 22388 17734 22508 17762
rect 22112 16046 22140 16408
rect 22284 16108 22336 16114
rect 22284 16050 22336 16056
rect 22100 16040 22152 16046
rect 22192 16040 22244 16046
rect 22100 15982 22152 15988
rect 22190 16008 22192 16017
rect 22244 16008 22246 16017
rect 22190 15943 22246 15952
rect 22098 15328 22154 15337
rect 22098 15263 22154 15272
rect 22006 14920 22062 14929
rect 22006 14855 22062 14864
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21364 13796 21416 13802
rect 21364 13738 21416 13744
rect 21178 12608 21234 12617
rect 21178 12543 21234 12552
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21100 12102 21128 12242
rect 21284 12209 21312 12242
rect 21376 12220 21404 13738
rect 21546 13560 21602 13569
rect 21546 13495 21602 13504
rect 21560 13462 21588 13495
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21456 12232 21508 12238
rect 21270 12200 21326 12209
rect 21376 12192 21456 12220
rect 21456 12174 21508 12180
rect 21270 12135 21326 12144
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20996 10736 21048 10742
rect 20902 10704 20958 10713
rect 20996 10678 21048 10684
rect 21100 10674 21128 10746
rect 20902 10639 20958 10648
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20996 10600 21048 10606
rect 20732 10526 20852 10554
rect 20916 10560 20996 10588
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20548 8498 20576 8910
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20640 7970 20668 8434
rect 20732 8430 20760 10526
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20824 10266 20852 10406
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20916 9722 20944 10560
rect 20996 10542 21048 10548
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21008 10266 21036 10406
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 21192 10062 21220 12038
rect 21284 10810 21312 12135
rect 21454 11792 21510 11801
rect 21454 11727 21510 11736
rect 21548 11756 21600 11762
rect 21468 11626 21496 11727
rect 21548 11698 21600 11704
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21362 10704 21418 10713
rect 21272 10668 21324 10674
rect 21362 10639 21418 10648
rect 21456 10668 21508 10674
rect 21272 10610 21324 10616
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 20824 9489 20852 9522
rect 20810 9480 20866 9489
rect 20916 9450 20944 9522
rect 20810 9415 20866 9424
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20640 7942 20760 7970
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7546 20576 7686
rect 20640 7562 20668 7822
rect 20732 7750 20760 7942
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20536 7540 20588 7546
rect 20640 7534 20760 7562
rect 20536 7482 20588 7488
rect 20456 6798 20484 7482
rect 20732 7410 20760 7534
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20548 6458 20576 6734
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 20640 3738 20668 7346
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20732 7002 20760 7210
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 5914 20760 6054
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20732 4826 20760 5578
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 16500 2310 16528 2366
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17880 2310 17908 2926
rect 18984 2650 19012 3470
rect 19536 3466 19564 3674
rect 20824 3534 20852 6598
rect 20916 6322 20944 9386
rect 21008 9110 21036 9522
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21086 7984 21142 7993
rect 21086 7919 21142 7928
rect 21100 7886 21128 7919
rect 21088 7880 21140 7886
rect 21180 7880 21232 7886
rect 21088 7822 21140 7828
rect 21178 7848 21180 7857
rect 21232 7848 21234 7857
rect 21100 7478 21128 7822
rect 21178 7783 21234 7792
rect 21088 7472 21140 7478
rect 21088 7414 21140 7420
rect 21088 6384 21140 6390
rect 21140 6332 21220 6338
rect 21088 6326 21220 6332
rect 20904 6316 20956 6322
rect 21100 6310 21220 6326
rect 20904 6258 20956 6264
rect 20916 5914 20944 6258
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 21192 5234 21220 6310
rect 21284 5914 21312 10610
rect 21376 8537 21404 10639
rect 21456 10610 21508 10616
rect 21468 9994 21496 10610
rect 21560 10577 21588 11698
rect 21546 10568 21602 10577
rect 21546 10503 21602 10512
rect 21560 10062 21588 10503
rect 21652 10169 21680 13874
rect 22112 12850 22140 15263
rect 22296 12986 22324 16050
rect 22388 13802 22416 17734
rect 22572 17678 22600 19343
rect 22652 19314 22704 19320
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22466 17368 22522 17377
rect 22466 17303 22522 17312
rect 22376 13796 22428 13802
rect 22376 13738 22428 13744
rect 22480 13734 22508 17303
rect 22558 17232 22614 17241
rect 22558 17167 22614 17176
rect 22652 17196 22704 17202
rect 22572 17134 22600 17167
rect 22652 17138 22704 17144
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22560 16992 22612 16998
rect 22664 16946 22692 17138
rect 22612 16940 22692 16946
rect 22560 16934 22692 16940
rect 22572 16918 22692 16934
rect 22572 14482 22600 16918
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22664 16425 22692 16594
rect 22650 16416 22706 16425
rect 22650 16351 22706 16360
rect 22652 15972 22704 15978
rect 22652 15914 22704 15920
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22664 14346 22692 15914
rect 22756 14890 22784 21966
rect 22940 21298 22968 24754
rect 23020 22160 23072 22166
rect 23018 22128 23020 22137
rect 23072 22128 23074 22137
rect 23018 22063 23074 22072
rect 23124 22030 23152 26318
rect 23216 25480 23244 26726
rect 23400 26518 23428 26846
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23296 26512 23348 26518
rect 23294 26480 23296 26489
rect 23388 26512 23440 26518
rect 23348 26480 23350 26489
rect 23388 26454 23440 26460
rect 23294 26415 23350 26424
rect 23296 25492 23348 25498
rect 23216 25452 23296 25480
rect 23296 25434 23348 25440
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23216 22710 23244 24142
rect 23204 22704 23256 22710
rect 23204 22646 23256 22652
rect 23204 22228 23256 22234
rect 23204 22170 23256 22176
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21350 23152 21966
rect 23112 21344 23164 21350
rect 22940 21270 23060 21298
rect 23112 21286 23164 21292
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22848 20466 22876 20742
rect 22940 20466 22968 21082
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 22836 19440 22888 19446
rect 22834 19408 22836 19417
rect 22888 19408 22890 19417
rect 22834 19343 22890 19352
rect 22836 17672 22888 17678
rect 22834 17640 22836 17649
rect 22888 17640 22890 17649
rect 22834 17575 22890 17584
rect 22836 17536 22888 17542
rect 22836 17478 22888 17484
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 22664 14056 22692 14282
rect 22572 14028 22692 14056
rect 22572 13938 22600 14028
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22468 13728 22520 13734
rect 22520 13688 22600 13716
rect 22468 13670 22520 13676
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 21744 12442 21772 12786
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21638 10160 21694 10169
rect 21638 10095 21694 10104
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21362 8528 21418 8537
rect 21362 8463 21418 8472
rect 21468 6730 21496 9930
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21560 8430 21588 8570
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21652 7177 21680 7346
rect 21638 7168 21694 7177
rect 21638 7103 21694 7112
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21546 6896 21602 6905
rect 21546 6831 21602 6840
rect 21456 6724 21508 6730
rect 21456 6666 21508 6672
rect 21468 6458 21496 6666
rect 21560 6662 21588 6831
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21652 6458 21680 6938
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21560 5710 21588 6326
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21652 5710 21680 6054
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21546 5400 21602 5409
rect 21546 5335 21602 5344
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21086 5128 21142 5137
rect 21086 5063 21088 5072
rect 21140 5063 21142 5072
rect 21088 5034 21140 5040
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 20994 4176 21050 4185
rect 21100 4146 21128 4762
rect 20994 4111 20996 4120
rect 21048 4111 21050 4120
rect 21088 4140 21140 4146
rect 20996 4082 21048 4088
rect 21088 4082 21140 4088
rect 21088 3664 21140 3670
rect 21086 3632 21088 3641
rect 21140 3632 21142 3641
rect 21192 3602 21220 5170
rect 21272 4752 21324 4758
rect 21272 4694 21324 4700
rect 21364 4752 21416 4758
rect 21364 4694 21416 4700
rect 21284 3942 21312 4694
rect 21376 4554 21404 4694
rect 21364 4548 21416 4554
rect 21364 4490 21416 4496
rect 21376 4146 21404 4490
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21468 4010 21496 4082
rect 21560 4078 21588 5335
rect 21744 5302 21772 12174
rect 21836 10810 21864 12582
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 21928 7954 21956 12786
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22112 12374 22140 12582
rect 22282 12472 22338 12481
rect 22282 12407 22338 12416
rect 22100 12368 22152 12374
rect 22100 12310 22152 12316
rect 22296 12238 22324 12407
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22296 11830 22324 12038
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22112 8090 22140 11290
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22112 7954 22140 8026
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 21928 7478 21956 7890
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 22008 7404 22060 7410
rect 22204 7392 22232 9522
rect 22282 9480 22338 9489
rect 22282 9415 22284 9424
rect 22336 9415 22338 9424
rect 22284 9386 22336 9392
rect 22388 7410 22416 12582
rect 22480 12442 22508 12650
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22480 12102 22508 12378
rect 22572 12374 22600 13688
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22664 11778 22692 13874
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22756 12238 22784 13466
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22572 11750 22692 11778
rect 22572 10538 22600 11750
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22664 11150 22692 11494
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22560 10532 22612 10538
rect 22560 10474 22612 10480
rect 22664 10266 22692 11086
rect 22756 10606 22784 11086
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22480 9722 22508 10066
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22560 9716 22612 9722
rect 22756 9704 22784 10542
rect 22612 9676 22784 9704
rect 22560 9658 22612 9664
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22480 7410 22508 7686
rect 22060 7364 22232 7392
rect 22376 7404 22428 7410
rect 22008 7346 22060 7352
rect 22376 7346 22428 7352
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22020 6866 22048 7346
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22112 7002 22140 7210
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 21824 6384 21876 6390
rect 21824 6326 21876 6332
rect 21836 5710 21864 6326
rect 22388 6118 22416 7346
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22572 5846 22600 9114
rect 22848 7410 22876 17478
rect 22940 14346 22968 20402
rect 23032 18426 23060 21270
rect 23112 20868 23164 20874
rect 23216 20856 23244 22170
rect 23164 20828 23244 20856
rect 23112 20810 23164 20816
rect 23124 18970 23152 20810
rect 23308 20369 23336 25434
rect 23400 25362 23428 26454
rect 23492 25702 23520 26726
rect 23676 26246 23704 29514
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23768 28150 23796 28358
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23768 27470 23796 28086
rect 23756 27464 23808 27470
rect 23756 27406 23808 27412
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23952 26926 23980 27406
rect 23940 26920 23992 26926
rect 23940 26862 23992 26868
rect 23664 26240 23716 26246
rect 23664 26182 23716 26188
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 23480 25696 23532 25702
rect 23480 25638 23532 25644
rect 23388 25356 23440 25362
rect 23388 25298 23440 25304
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23400 24274 23428 24754
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23400 23322 23428 24210
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23492 22642 23520 25638
rect 23584 24614 23612 25842
rect 23676 25430 23704 25842
rect 23664 25424 23716 25430
rect 23664 25366 23716 25372
rect 23860 24818 23888 25842
rect 23952 25809 23980 25842
rect 23938 25800 23994 25809
rect 23938 25735 23994 25744
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 23756 24744 23808 24750
rect 23676 24704 23756 24732
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23676 24138 23704 24704
rect 23756 24686 23808 24692
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23768 22642 23796 24550
rect 23952 23798 23980 25638
rect 24044 24954 24072 31583
rect 24136 28422 24164 31894
rect 24320 31822 24348 32166
rect 24308 31816 24360 31822
rect 24308 31758 24360 31764
rect 24228 31482 24348 31498
rect 24228 31476 24360 31482
rect 24228 31470 24308 31476
rect 24228 30666 24256 31470
rect 24308 31418 24360 31424
rect 24308 31272 24360 31278
rect 24308 31214 24360 31220
rect 24320 30666 24348 31214
rect 24216 30660 24268 30666
rect 24216 30602 24268 30608
rect 24308 30660 24360 30666
rect 24308 30602 24360 30608
rect 24228 28778 24256 30602
rect 24320 30326 24348 30602
rect 24308 30320 24360 30326
rect 24308 30262 24360 30268
rect 24228 28750 24348 28778
rect 24412 28762 24440 32846
rect 24504 31521 24532 32966
rect 24596 31958 24624 32982
rect 24688 32910 24716 33594
rect 24676 32904 24728 32910
rect 24676 32846 24728 32852
rect 24674 32464 24730 32473
rect 24674 32399 24730 32408
rect 24584 31952 24636 31958
rect 24584 31894 24636 31900
rect 24688 31754 24716 32399
rect 24780 31890 24808 34138
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 24872 33114 24900 33934
rect 25056 33658 25084 34546
rect 25332 34066 25360 34546
rect 25320 34060 25372 34066
rect 25320 34002 25372 34008
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 25320 32972 25372 32978
rect 25320 32914 25372 32920
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 25044 32904 25096 32910
rect 25096 32864 25176 32892
rect 25044 32846 25096 32852
rect 24872 32502 24900 32846
rect 24952 32768 25004 32774
rect 25148 32756 25176 32864
rect 25228 32768 25280 32774
rect 25004 32728 25084 32756
rect 25148 32728 25228 32756
rect 24952 32710 25004 32716
rect 24860 32496 24912 32502
rect 24860 32438 24912 32444
rect 24768 31884 24820 31890
rect 24768 31826 24820 31832
rect 24596 31726 24716 31754
rect 24768 31748 24820 31754
rect 24596 31686 24624 31726
rect 24768 31690 24820 31696
rect 24952 31748 25004 31754
rect 24952 31690 25004 31696
rect 24584 31680 24636 31686
rect 24584 31622 24636 31628
rect 24490 31512 24546 31521
rect 24490 31447 24546 31456
rect 24492 30320 24544 30326
rect 24492 30262 24544 30268
rect 24504 29782 24532 30262
rect 24492 29776 24544 29782
rect 24492 29718 24544 29724
rect 24504 29238 24532 29718
rect 24492 29232 24544 29238
rect 24492 29174 24544 29180
rect 24124 28416 24176 28422
rect 24124 28358 24176 28364
rect 24216 25764 24268 25770
rect 24216 25706 24268 25712
rect 24228 25294 24256 25706
rect 24216 25288 24268 25294
rect 24216 25230 24268 25236
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 24228 24614 24256 25230
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 24032 24404 24084 24410
rect 24032 24346 24084 24352
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23952 22642 23980 23734
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23400 20534 23428 20878
rect 23492 20806 23520 22578
rect 23952 22522 23980 22578
rect 23860 22494 23980 22522
rect 23756 22432 23808 22438
rect 23756 22374 23808 22380
rect 23768 22234 23796 22374
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23756 21956 23808 21962
rect 23756 21898 23808 21904
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23584 20398 23612 21082
rect 23676 20942 23704 21286
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23676 20806 23704 20878
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23572 20392 23624 20398
rect 23294 20360 23350 20369
rect 23676 20369 23704 20402
rect 23572 20334 23624 20340
rect 23662 20360 23718 20369
rect 23294 20295 23350 20304
rect 23662 20295 23718 20304
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23388 19712 23440 19718
rect 23294 19680 23350 19689
rect 23388 19654 23440 19660
rect 23294 19615 23350 19624
rect 23202 19544 23258 19553
rect 23202 19479 23204 19488
rect 23256 19479 23258 19488
rect 23204 19450 23256 19456
rect 23308 19446 23336 19615
rect 23296 19440 23348 19446
rect 23202 19408 23258 19417
rect 23296 19382 23348 19388
rect 23202 19343 23258 19352
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23032 17814 23060 18362
rect 23110 18184 23166 18193
rect 23110 18119 23166 18128
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 23124 17678 23152 18119
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23032 17377 23060 17614
rect 23018 17368 23074 17377
rect 23018 17303 23074 17312
rect 23124 16538 23152 17614
rect 23216 16726 23244 19343
rect 23400 19310 23428 19654
rect 23296 19304 23348 19310
rect 23294 19272 23296 19281
rect 23388 19304 23440 19310
rect 23348 19272 23350 19281
rect 23388 19246 23440 19252
rect 23294 19207 23350 19216
rect 23294 18864 23350 18873
rect 23294 18799 23350 18808
rect 23308 18766 23336 18799
rect 23492 18766 23520 19722
rect 23768 19334 23796 21898
rect 23860 21026 23888 22494
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23952 21146 23980 22374
rect 24044 21622 24072 24346
rect 24228 24070 24256 24550
rect 24320 24206 24348 28750
rect 24400 28756 24452 28762
rect 24400 28698 24452 28704
rect 24412 28642 24440 28698
rect 24596 28694 24624 31622
rect 24780 31396 24808 31690
rect 24964 31657 24992 31690
rect 24950 31648 25006 31657
rect 24950 31583 25006 31592
rect 24780 31368 24900 31396
rect 24872 30734 24900 31368
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 24860 30728 24912 30734
rect 24780 30676 24860 30682
rect 24780 30670 24912 30676
rect 24780 30654 24900 30670
rect 24780 30598 24808 30654
rect 24768 30592 24820 30598
rect 24860 30592 24912 30598
rect 24768 30534 24820 30540
rect 24858 30560 24860 30569
rect 24912 30560 24914 30569
rect 24858 30495 24914 30504
rect 24872 30394 24900 30495
rect 24860 30388 24912 30394
rect 24860 30330 24912 30336
rect 24964 29306 24992 31214
rect 25056 30852 25084 32728
rect 25228 32710 25280 32716
rect 25332 32570 25360 32914
rect 25424 32910 25452 34682
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 26148 34536 26200 34542
rect 26148 34478 26200 34484
rect 25504 34060 25556 34066
rect 25504 34002 25556 34008
rect 25516 33454 25544 34002
rect 26160 33930 26188 34478
rect 25780 33924 25832 33930
rect 25780 33866 25832 33872
rect 26148 33924 26200 33930
rect 26148 33866 26200 33872
rect 25792 33658 25820 33866
rect 25780 33652 25832 33658
rect 25780 33594 25832 33600
rect 26056 33516 26108 33522
rect 26056 33458 26108 33464
rect 25504 33448 25556 33454
rect 25504 33390 25556 33396
rect 25964 33448 26016 33454
rect 25964 33390 26016 33396
rect 25516 32910 25544 33390
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 25504 32904 25556 32910
rect 25504 32846 25556 32852
rect 25780 32904 25832 32910
rect 25780 32846 25832 32852
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25136 32224 25188 32230
rect 25136 32166 25188 32172
rect 25148 31958 25176 32166
rect 25136 31952 25188 31958
rect 25136 31894 25188 31900
rect 25332 31822 25360 32506
rect 25594 32328 25650 32337
rect 25594 32263 25650 32272
rect 25608 32026 25636 32263
rect 25688 32224 25740 32230
rect 25688 32166 25740 32172
rect 25504 32020 25556 32026
rect 25504 31962 25556 31968
rect 25596 32020 25648 32026
rect 25596 31962 25648 31968
rect 25320 31816 25372 31822
rect 25372 31776 25452 31804
rect 25320 31758 25372 31764
rect 25228 31680 25280 31686
rect 25228 31622 25280 31628
rect 25318 31648 25374 31657
rect 25240 31210 25268 31622
rect 25318 31583 25374 31592
rect 25332 31414 25360 31583
rect 25320 31408 25372 31414
rect 25320 31350 25372 31356
rect 25424 31278 25452 31776
rect 25412 31272 25464 31278
rect 25412 31214 25464 31220
rect 25228 31204 25280 31210
rect 25228 31146 25280 31152
rect 25056 30824 25176 30852
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 24952 29300 25004 29306
rect 24952 29242 25004 29248
rect 24584 28688 24636 28694
rect 24412 28626 24532 28642
rect 24584 28630 24636 28636
rect 24768 28688 24820 28694
rect 24768 28630 24820 28636
rect 24412 28620 24544 28626
rect 24412 28614 24492 28620
rect 24492 28562 24544 28568
rect 24596 28370 24624 28630
rect 24780 28490 24808 28630
rect 25056 28558 25084 30670
rect 25148 28694 25176 30824
rect 25424 30598 25452 31214
rect 25412 30592 25464 30598
rect 25412 30534 25464 30540
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25240 29481 25268 29514
rect 25226 29472 25282 29481
rect 25226 29407 25282 29416
rect 25136 28688 25188 28694
rect 25136 28630 25188 28636
rect 24860 28552 24912 28558
rect 24952 28552 25004 28558
rect 24860 28494 24912 28500
rect 24950 28520 24952 28529
rect 25044 28552 25096 28558
rect 25004 28520 25006 28529
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24412 28342 24624 28370
rect 24676 28416 24728 28422
rect 24676 28358 24728 28364
rect 24412 24857 24440 28342
rect 24584 28212 24636 28218
rect 24584 28154 24636 28160
rect 24490 26888 24546 26897
rect 24490 26823 24546 26832
rect 24504 26790 24532 26823
rect 24492 26784 24544 26790
rect 24492 26726 24544 26732
rect 24398 24848 24454 24857
rect 24398 24783 24454 24792
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 24216 24064 24268 24070
rect 24216 24006 24268 24012
rect 24228 23118 24256 24006
rect 24216 23112 24268 23118
rect 24216 23054 24268 23060
rect 24124 23044 24176 23050
rect 24124 22986 24176 22992
rect 24136 22642 24164 22986
rect 24228 22642 24256 23054
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24032 21616 24084 21622
rect 24032 21558 24084 21564
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23860 20998 23980 21026
rect 23584 19306 23796 19334
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 23124 16510 23244 16538
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23018 16008 23074 16017
rect 23018 15943 23074 15952
rect 23032 15910 23060 15943
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 23124 15638 23152 16390
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23216 15502 23244 16510
rect 23020 15496 23072 15502
rect 23204 15496 23256 15502
rect 23020 15438 23072 15444
rect 23202 15464 23204 15473
rect 23256 15464 23258 15473
rect 23032 15162 23060 15438
rect 23202 15399 23258 15408
rect 23020 15156 23072 15162
rect 23020 15098 23072 15104
rect 23032 14618 23060 15098
rect 23020 14612 23072 14618
rect 23020 14554 23072 14560
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 23216 13938 23244 14418
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 22940 13308 22968 13738
rect 22940 13280 23060 13308
rect 23032 12918 23060 13280
rect 23020 12912 23072 12918
rect 23020 12854 23072 12860
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 22940 10826 22968 12786
rect 23032 12306 23060 12854
rect 23216 12646 23244 13874
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 23216 12481 23244 12582
rect 23202 12472 23258 12481
rect 23202 12407 23258 12416
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23032 11898 23060 12038
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 23216 11830 23244 12038
rect 23204 11824 23256 11830
rect 23204 11766 23256 11772
rect 23308 11354 23336 18566
rect 23492 18358 23520 18702
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23400 16658 23428 17138
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23584 16266 23612 19306
rect 23664 18692 23716 18698
rect 23664 18634 23716 18640
rect 23676 18290 23704 18634
rect 23952 18465 23980 20998
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 23938 18456 23994 18465
rect 23938 18391 23994 18400
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23676 17882 23704 18226
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 23768 17678 23796 18226
rect 23952 18057 23980 18226
rect 23938 18048 23994 18057
rect 23938 17983 23994 17992
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 24044 16794 24072 20878
rect 24136 20534 24164 22578
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24216 21616 24268 21622
rect 24216 21558 24268 21564
rect 24228 20856 24256 21558
rect 24320 20924 24348 22510
rect 24412 22409 24440 22578
rect 24398 22400 24454 22409
rect 24398 22335 24454 22344
rect 24504 21690 24532 26726
rect 24596 25906 24624 28154
rect 24688 28014 24716 28358
rect 24768 28076 24820 28082
rect 24768 28018 24820 28024
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24780 26994 24808 28018
rect 24872 27713 24900 28494
rect 25148 28529 25176 28630
rect 25044 28494 25096 28500
rect 25134 28520 25190 28529
rect 24950 28455 25006 28464
rect 25056 28150 25084 28494
rect 25134 28455 25190 28464
rect 25410 28248 25466 28257
rect 25136 28212 25188 28218
rect 25410 28183 25466 28192
rect 25136 28154 25188 28160
rect 25044 28144 25096 28150
rect 25044 28086 25096 28092
rect 24858 27704 24914 27713
rect 24858 27639 24914 27648
rect 25148 27538 25176 28154
rect 25136 27532 25188 27538
rect 25136 27474 25188 27480
rect 24952 27124 25004 27130
rect 24952 27066 25004 27072
rect 25044 27124 25096 27130
rect 25044 27066 25096 27072
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24780 26858 24808 26930
rect 24768 26852 24820 26858
rect 24768 26794 24820 26800
rect 24964 26586 24992 27066
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 24964 25974 24992 26522
rect 25056 26450 25084 27066
rect 25148 27062 25176 27474
rect 25136 27056 25188 27062
rect 25136 26998 25188 27004
rect 25044 26444 25096 26450
rect 25044 26386 25096 26392
rect 24952 25968 25004 25974
rect 24952 25910 25004 25916
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24872 25498 24900 25842
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 25056 25430 25084 26386
rect 25424 26382 25452 28183
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 25228 25968 25280 25974
rect 25228 25910 25280 25916
rect 25044 25424 25096 25430
rect 25044 25366 25096 25372
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24584 22228 24636 22234
rect 24584 22170 24636 22176
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24504 21078 24532 21422
rect 24596 21078 24624 22170
rect 24492 21072 24544 21078
rect 24492 21014 24544 21020
rect 24584 21072 24636 21078
rect 24584 21014 24636 21020
rect 24492 20936 24544 20942
rect 24320 20896 24492 20924
rect 24492 20878 24544 20884
rect 24228 20828 24348 20856
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24122 19408 24178 19417
rect 24122 19343 24124 19352
rect 24176 19343 24178 19352
rect 24124 19314 24176 19320
rect 24228 18698 24256 20402
rect 24320 20398 24348 20828
rect 24308 20392 24360 20398
rect 24308 20334 24360 20340
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24412 19174 24440 19314
rect 24308 19168 24360 19174
rect 24308 19110 24360 19116
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24320 18970 24348 19110
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24216 18692 24268 18698
rect 24216 18634 24268 18640
rect 24228 18358 24256 18634
rect 24216 18352 24268 18358
rect 24216 18294 24268 18300
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 23584 16238 23888 16266
rect 23664 16176 23716 16182
rect 23664 16118 23716 16124
rect 23480 16040 23532 16046
rect 23478 16008 23480 16017
rect 23532 16008 23534 16017
rect 23478 15943 23534 15952
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23400 13802 23428 14350
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23492 12918 23520 14962
rect 23584 14414 23612 15030
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23572 12640 23624 12646
rect 23570 12608 23572 12617
rect 23624 12608 23626 12617
rect 23570 12543 23626 12552
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23032 11150 23060 11290
rect 23400 11150 23428 12310
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23492 11354 23520 11834
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23112 11076 23164 11082
rect 23112 11018 23164 11024
rect 22940 10798 23060 10826
rect 22928 10736 22980 10742
rect 22926 10704 22928 10713
rect 22980 10704 22982 10713
rect 22926 10639 22982 10648
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 9178 22968 9862
rect 23032 9654 23060 10798
rect 23124 10674 23152 11018
rect 23584 11014 23612 12174
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 23110 10296 23166 10305
rect 23110 10231 23166 10240
rect 23204 10260 23256 10266
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 23032 7834 23060 9590
rect 23124 9042 23152 10231
rect 23204 10202 23256 10208
rect 23216 9382 23244 10202
rect 23478 10160 23534 10169
rect 23478 10095 23534 10104
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23296 9376 23348 9382
rect 23400 9353 23428 9522
rect 23296 9318 23348 9324
rect 23386 9344 23442 9353
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23308 8974 23336 9318
rect 23386 9279 23442 9288
rect 23400 9178 23428 9279
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23112 8832 23164 8838
rect 23112 8774 23164 8780
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 23124 8362 23152 8774
rect 23308 8498 23336 8774
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 23112 8356 23164 8362
rect 23112 8298 23164 8304
rect 23124 8090 23152 8298
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23216 7868 23244 8366
rect 23296 8288 23348 8294
rect 23400 8276 23428 8910
rect 23492 8786 23520 10095
rect 23676 9738 23704 16118
rect 23756 14408 23808 14414
rect 23756 14350 23808 14356
rect 23584 9710 23704 9738
rect 23584 8906 23612 9710
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23676 8974 23704 9522
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23572 8900 23624 8906
rect 23572 8842 23624 8848
rect 23492 8758 23612 8786
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23348 8248 23428 8276
rect 23296 8230 23348 8236
rect 23308 8090 23336 8230
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23492 7886 23520 8570
rect 23584 8537 23612 8758
rect 23570 8528 23626 8537
rect 23570 8463 23626 8472
rect 23584 8430 23612 8463
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23480 7880 23532 7886
rect 23216 7840 23480 7868
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22560 5840 22612 5846
rect 22560 5782 22612 5788
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 22006 5400 22062 5409
rect 22006 5335 22008 5344
rect 22060 5335 22062 5344
rect 22008 5306 22060 5312
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 21640 5092 21692 5098
rect 21640 5034 21692 5040
rect 21652 4622 21680 5034
rect 21744 4758 21772 5238
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22204 4826 22232 5170
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21272 3936 21324 3942
rect 21272 3878 21324 3884
rect 21086 3567 21142 3576
rect 21180 3596 21232 3602
rect 21100 3534 21128 3567
rect 21180 3538 21232 3544
rect 21284 3534 21312 3878
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 20442 3224 20498 3233
rect 20442 3159 20498 3168
rect 20456 3126 20484 3159
rect 20444 3120 20496 3126
rect 20444 3062 20496 3068
rect 21468 3058 21496 3538
rect 21836 3534 21864 4558
rect 22192 4072 22244 4078
rect 22190 4040 22192 4049
rect 22244 4040 22246 4049
rect 22190 3975 22246 3984
rect 21916 3936 21968 3942
rect 21968 3896 22048 3924
rect 21916 3878 21968 3884
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19076 2514 19104 2790
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 19996 800 20024 2994
rect 21836 2922 21864 3470
rect 21914 3224 21970 3233
rect 21914 3159 21970 3168
rect 21824 2916 21876 2922
rect 21824 2858 21876 2864
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 20732 2446 20760 2790
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20640 800 20668 2246
rect 21284 800 21312 2790
rect 21928 2774 21956 3159
rect 22020 2802 22048 3896
rect 22204 3670 22232 3975
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22112 3194 22140 3334
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22204 3126 22232 3606
rect 22296 3466 22324 4558
rect 22480 3942 22508 5170
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22572 3602 22600 4966
rect 22664 4690 22692 7142
rect 22834 6896 22890 6905
rect 22834 6831 22890 6840
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 22756 5914 22784 6190
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 22848 5710 22876 6831
rect 22940 6730 22968 7822
rect 23032 7806 23152 7834
rect 23480 7822 23532 7828
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 23032 7410 23060 7686
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 23124 6322 23152 7806
rect 23492 7206 23520 7822
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 23124 4826 23152 6258
rect 23584 5710 23612 8026
rect 23676 7274 23704 8910
rect 23768 8634 23796 14350
rect 23860 12209 23888 16238
rect 23952 16114 23980 16526
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 23952 12442 23980 16050
rect 24044 15026 24072 16050
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 23846 12200 23902 12209
rect 23846 12135 23902 12144
rect 23940 12164 23992 12170
rect 23860 10810 23888 12135
rect 23940 12106 23992 12112
rect 23952 12073 23980 12106
rect 23938 12064 23994 12073
rect 23938 11999 23994 12008
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 23860 10470 23888 10542
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 9994 23888 10406
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23860 9722 23888 9930
rect 23848 9716 23900 9722
rect 23848 9658 23900 9664
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23860 8430 23888 9658
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23768 7954 23796 8366
rect 23756 7948 23808 7954
rect 23756 7890 23808 7896
rect 23664 7268 23716 7274
rect 23664 7210 23716 7216
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23768 5710 23796 6394
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23952 5574 23980 11999
rect 24030 11928 24086 11937
rect 24030 11863 24086 11872
rect 24044 11762 24072 11863
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 24030 9480 24086 9489
rect 24030 9415 24086 9424
rect 24044 6390 24072 9415
rect 24136 6866 24164 18226
rect 24216 16720 24268 16726
rect 24216 16662 24268 16668
rect 24228 16182 24256 16662
rect 24320 16182 24348 18702
rect 24412 18086 24440 19110
rect 24400 18080 24452 18086
rect 24400 18022 24452 18028
rect 24504 17814 24532 20878
rect 24596 18426 24624 21014
rect 24688 19514 24716 24686
rect 24872 24256 24900 25094
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24780 24228 24900 24256
rect 24780 23746 24808 24228
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24872 23866 24900 24074
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24780 23718 24900 23746
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24780 20602 24808 20878
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24768 20392 24820 20398
rect 24768 20334 24820 20340
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24780 19446 24808 20334
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24676 18760 24728 18766
rect 24728 18720 24808 18748
rect 24676 18702 24728 18708
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24674 18320 24730 18329
rect 24674 18255 24730 18264
rect 24582 18184 24638 18193
rect 24688 18154 24716 18255
rect 24582 18119 24638 18128
rect 24676 18148 24728 18154
rect 24492 17808 24544 17814
rect 24492 17750 24544 17756
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24216 16176 24268 16182
rect 24216 16118 24268 16124
rect 24308 16176 24360 16182
rect 24308 16118 24360 16124
rect 24216 14952 24268 14958
rect 24214 14920 24216 14929
rect 24268 14920 24270 14929
rect 24214 14855 24270 14864
rect 24214 13968 24270 13977
rect 24214 13903 24216 13912
rect 24268 13903 24270 13912
rect 24412 13920 24440 17138
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24504 14550 24532 16526
rect 24596 16114 24624 18119
rect 24676 18090 24728 18096
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24688 16522 24716 17818
rect 24676 16516 24728 16522
rect 24676 16458 24728 16464
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24688 15162 24716 16458
rect 24780 16114 24808 18720
rect 24872 18222 24900 23718
rect 24964 21010 24992 24754
rect 25044 24676 25096 24682
rect 25044 24618 25096 24624
rect 25056 23662 25084 24618
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25148 24206 25176 24550
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 25148 23798 25176 24142
rect 25240 24138 25268 25910
rect 25320 25900 25372 25906
rect 25320 25842 25372 25848
rect 25332 25362 25360 25842
rect 25410 25392 25466 25401
rect 25320 25356 25372 25362
rect 25410 25327 25466 25336
rect 25320 25298 25372 25304
rect 25228 24132 25280 24138
rect 25228 24074 25280 24080
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25044 23656 25096 23662
rect 25240 23644 25268 24074
rect 25044 23598 25096 23604
rect 25148 23616 25268 23644
rect 25148 22166 25176 23616
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 25136 22160 25188 22166
rect 25136 22102 25188 22108
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24964 20602 24992 20946
rect 25148 20602 25176 21422
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25240 19378 25268 23258
rect 25332 23254 25360 25298
rect 25424 25294 25452 25327
rect 25412 25288 25464 25294
rect 25412 25230 25464 25236
rect 25410 23488 25466 23497
rect 25410 23423 25466 23432
rect 25320 23248 25372 23254
rect 25320 23190 25372 23196
rect 25424 22778 25452 23423
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 25424 22681 25452 22714
rect 25410 22672 25466 22681
rect 25410 22607 25466 22616
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25318 21040 25374 21049
rect 25318 20975 25374 20984
rect 25332 20874 25360 20975
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25134 18864 25190 18873
rect 25134 18799 25190 18808
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24964 17882 24992 18566
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24780 14822 24808 16050
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24492 14544 24544 14550
rect 24492 14486 24544 14492
rect 24492 13932 24544 13938
rect 24412 13892 24492 13920
rect 24216 13874 24268 13880
rect 24492 13874 24544 13880
rect 24504 13530 24532 13874
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24320 12238 24348 12582
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24412 12102 24440 12922
rect 24596 12442 24624 14758
rect 24688 14618 24716 14758
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24872 13977 24900 16526
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24964 16114 24992 16186
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24964 15434 24992 16050
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 24858 13968 24914 13977
rect 24858 13903 24914 13912
rect 24952 13932 25004 13938
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24872 12170 24900 13903
rect 24952 13874 25004 13880
rect 24964 12238 24992 13874
rect 25056 12866 25084 18158
rect 25148 17898 25176 18799
rect 25240 18766 25268 19314
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25148 17870 25268 17898
rect 25136 17808 25188 17814
rect 25136 17750 25188 17756
rect 25148 17202 25176 17750
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25240 16794 25268 17870
rect 25332 17202 25360 20810
rect 25424 18329 25452 22510
rect 25516 22250 25544 31962
rect 25608 31278 25636 31962
rect 25700 31822 25728 32166
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 25792 31686 25820 32846
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 25688 31680 25740 31686
rect 25688 31622 25740 31628
rect 25780 31680 25832 31686
rect 25780 31622 25832 31628
rect 25700 31521 25728 31622
rect 25686 31512 25742 31521
rect 25884 31482 25912 31758
rect 25686 31447 25742 31456
rect 25872 31476 25924 31482
rect 25872 31418 25924 31424
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 25596 31272 25648 31278
rect 25596 31214 25648 31220
rect 25596 31136 25648 31142
rect 25596 31078 25648 31084
rect 25608 29345 25636 31078
rect 25884 30938 25912 31282
rect 25872 30932 25924 30938
rect 25872 30874 25924 30880
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25688 29504 25740 29510
rect 25688 29446 25740 29452
rect 25594 29336 25650 29345
rect 25594 29271 25650 29280
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 25608 28762 25636 29038
rect 25596 28756 25648 28762
rect 25596 28698 25648 28704
rect 25700 28626 25728 29446
rect 25792 28801 25820 29582
rect 25778 28792 25834 28801
rect 25778 28727 25834 28736
rect 25792 28694 25820 28727
rect 25780 28688 25832 28694
rect 25780 28630 25832 28636
rect 25688 28620 25740 28626
rect 25688 28562 25740 28568
rect 25870 27976 25926 27985
rect 25870 27911 25872 27920
rect 25924 27911 25926 27920
rect 25872 27882 25924 27888
rect 25884 27674 25912 27882
rect 25872 27668 25924 27674
rect 25872 27610 25924 27616
rect 25870 27568 25926 27577
rect 25870 27503 25926 27512
rect 25884 27470 25912 27503
rect 25872 27464 25924 27470
rect 25872 27406 25924 27412
rect 25976 26874 26004 33390
rect 26068 32570 26096 33458
rect 26160 32774 26188 33866
rect 26436 33454 26464 34546
rect 26620 33930 26648 34886
rect 27356 34610 27384 34886
rect 27436 34740 27488 34746
rect 27436 34682 27488 34688
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 27344 34060 27396 34066
rect 27448 34048 27476 34682
rect 27396 34020 27476 34048
rect 27344 34002 27396 34008
rect 26608 33924 26660 33930
rect 26608 33866 26660 33872
rect 26884 33924 26936 33930
rect 26884 33866 26936 33872
rect 26700 33652 26752 33658
rect 26700 33594 26752 33600
rect 26424 33448 26476 33454
rect 26424 33390 26476 33396
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26608 33312 26660 33318
rect 26608 33254 26660 33260
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 26160 32230 26188 32710
rect 26252 32570 26280 33254
rect 26422 32736 26478 32745
rect 26422 32671 26478 32680
rect 26240 32564 26292 32570
rect 26240 32506 26292 32512
rect 26252 32366 26280 32506
rect 26436 32502 26464 32671
rect 26516 32564 26568 32570
rect 26516 32506 26568 32512
rect 26424 32496 26476 32502
rect 26424 32438 26476 32444
rect 26436 32366 26464 32438
rect 26528 32366 26556 32506
rect 26620 32434 26648 33254
rect 26712 32842 26740 33594
rect 26896 33386 26924 33866
rect 27448 33522 27476 34020
rect 27436 33516 27488 33522
rect 27436 33458 27488 33464
rect 27160 33448 27212 33454
rect 27160 33390 27212 33396
rect 26884 33380 26936 33386
rect 26884 33322 26936 33328
rect 26700 32836 26752 32842
rect 26700 32778 26752 32784
rect 26698 32464 26754 32473
rect 26608 32428 26660 32434
rect 26698 32399 26754 32408
rect 26608 32370 26660 32376
rect 26240 32360 26292 32366
rect 26240 32302 26292 32308
rect 26424 32360 26476 32366
rect 26424 32302 26476 32308
rect 26516 32360 26568 32366
rect 26516 32302 26568 32308
rect 26148 32224 26200 32230
rect 26424 32224 26476 32230
rect 26148 32166 26200 32172
rect 26252 32172 26424 32178
rect 26252 32166 26476 32172
rect 26252 32150 26464 32166
rect 26148 31884 26200 31890
rect 26252 31872 26280 32150
rect 26422 32056 26478 32065
rect 26422 31991 26478 32000
rect 26200 31844 26280 31872
rect 26148 31826 26200 31832
rect 26436 31822 26464 31991
rect 26424 31816 26476 31822
rect 26712 31793 26740 32399
rect 26792 32224 26844 32230
rect 26792 32166 26844 32172
rect 26424 31758 26476 31764
rect 26698 31784 26754 31793
rect 26148 31748 26200 31754
rect 26068 31708 26148 31736
rect 26068 27441 26096 31708
rect 26698 31719 26754 31728
rect 26148 31690 26200 31696
rect 26516 31680 26568 31686
rect 26238 31648 26294 31657
rect 26516 31622 26568 31628
rect 26238 31583 26294 31592
rect 26252 31346 26280 31583
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 26252 31113 26280 31282
rect 26528 31278 26556 31622
rect 26608 31408 26660 31414
rect 26608 31350 26660 31356
rect 26700 31408 26752 31414
rect 26700 31350 26752 31356
rect 26424 31272 26476 31278
rect 26424 31214 26476 31220
rect 26516 31272 26568 31278
rect 26516 31214 26568 31220
rect 26332 31136 26384 31142
rect 26238 31104 26294 31113
rect 26332 31078 26384 31084
rect 26238 31039 26294 31048
rect 26344 30784 26372 31078
rect 26436 30852 26464 31214
rect 26516 31136 26568 31142
rect 26620 31113 26648 31350
rect 26516 31078 26568 31084
rect 26606 31104 26662 31113
rect 26528 30920 26556 31078
rect 26606 31039 26662 31048
rect 26528 30892 26648 30920
rect 26436 30824 26556 30852
rect 26620 30841 26648 30892
rect 26344 30756 26464 30784
rect 26436 30666 26464 30756
rect 26332 30660 26384 30666
rect 26332 30602 26384 30608
rect 26424 30660 26476 30666
rect 26424 30602 26476 30608
rect 26148 30592 26200 30598
rect 26148 30534 26200 30540
rect 26160 30258 26188 30534
rect 26238 30424 26294 30433
rect 26238 30359 26294 30368
rect 26148 30252 26200 30258
rect 26148 30194 26200 30200
rect 26252 30190 26280 30359
rect 26240 30184 26292 30190
rect 26240 30126 26292 30132
rect 26344 29850 26372 30602
rect 26332 29844 26384 29850
rect 26332 29786 26384 29792
rect 26148 29776 26200 29782
rect 26200 29736 26280 29764
rect 26148 29718 26200 29724
rect 26252 29617 26280 29736
rect 26238 29608 26294 29617
rect 26148 29572 26200 29578
rect 26238 29543 26294 29552
rect 26148 29514 26200 29520
rect 26160 29170 26188 29514
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26054 27432 26110 27441
rect 26054 27367 26110 27376
rect 26056 27328 26108 27334
rect 26056 27270 26108 27276
rect 26068 26994 26096 27270
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 25976 26846 26096 26874
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 25596 26512 25648 26518
rect 25594 26480 25596 26489
rect 25648 26480 25650 26489
rect 25594 26415 25650 26424
rect 25778 26480 25834 26489
rect 25778 26415 25780 26424
rect 25832 26415 25834 26424
rect 25780 26386 25832 26392
rect 25884 26382 25912 26522
rect 25872 26376 25924 26382
rect 25872 26318 25924 26324
rect 25780 26308 25832 26314
rect 25780 26250 25832 26256
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25608 23050 25636 23666
rect 25596 23044 25648 23050
rect 25596 22986 25648 22992
rect 25608 22778 25636 22986
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25700 22642 25728 24890
rect 25792 24206 25820 26250
rect 25884 24954 25912 26318
rect 25872 24948 25924 24954
rect 25872 24890 25924 24896
rect 25870 24848 25926 24857
rect 25976 24818 26004 26726
rect 26068 26058 26096 26846
rect 26160 26228 26188 29106
rect 26252 28082 26280 29543
rect 26528 29186 26556 30824
rect 26606 30832 26662 30841
rect 26606 30767 26662 30776
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26620 30433 26648 30670
rect 26606 30424 26662 30433
rect 26606 30359 26662 30368
rect 26606 30288 26662 30297
rect 26606 30223 26608 30232
rect 26660 30223 26662 30232
rect 26608 30194 26660 30200
rect 26608 29572 26660 29578
rect 26608 29514 26660 29520
rect 26620 29306 26648 29514
rect 26712 29492 26740 31350
rect 26804 29646 26832 32166
rect 26896 31498 26924 33322
rect 27172 32774 27200 33390
rect 27540 32910 27568 35022
rect 27804 35012 27856 35018
rect 27804 34954 27856 34960
rect 27620 34468 27672 34474
rect 27620 34410 27672 34416
rect 27632 34134 27660 34410
rect 27620 34128 27672 34134
rect 27620 34070 27672 34076
rect 27712 33448 27764 33454
rect 27712 33390 27764 33396
rect 27724 32978 27752 33390
rect 27712 32972 27764 32978
rect 27712 32914 27764 32920
rect 27528 32904 27580 32910
rect 27250 32872 27306 32881
rect 27528 32846 27580 32852
rect 27250 32807 27306 32816
rect 27160 32768 27212 32774
rect 27160 32710 27212 32716
rect 26976 32360 27028 32366
rect 26976 32302 27028 32308
rect 26988 31657 27016 32302
rect 27172 31822 27200 32710
rect 27264 31822 27292 32807
rect 27528 32496 27580 32502
rect 27712 32496 27764 32502
rect 27528 32438 27580 32444
rect 27632 32456 27712 32484
rect 27344 32020 27396 32026
rect 27344 31962 27396 31968
rect 27356 31890 27384 31962
rect 27344 31884 27396 31890
rect 27344 31826 27396 31832
rect 27068 31816 27120 31822
rect 27066 31784 27068 31793
rect 27160 31816 27212 31822
rect 27120 31784 27122 31793
rect 27160 31758 27212 31764
rect 27252 31816 27304 31822
rect 27436 31816 27488 31822
rect 27252 31758 27304 31764
rect 27356 31764 27436 31770
rect 27356 31758 27488 31764
rect 27066 31719 27122 31728
rect 26974 31648 27030 31657
rect 27030 31606 27108 31634
rect 26974 31583 27030 31592
rect 26896 31470 27016 31498
rect 26884 31340 26936 31346
rect 26884 31282 26936 31288
rect 26896 30394 26924 31282
rect 26884 30388 26936 30394
rect 26884 30330 26936 30336
rect 26884 30048 26936 30054
rect 26884 29990 26936 29996
rect 26896 29646 26924 29990
rect 26988 29714 27016 31470
rect 27080 30734 27108 31606
rect 27264 31521 27292 31758
rect 27356 31742 27476 31758
rect 27250 31512 27306 31521
rect 27250 31447 27306 31456
rect 27356 31396 27384 31742
rect 27540 31686 27568 32438
rect 27632 31958 27660 32456
rect 27712 32438 27764 32444
rect 27712 32360 27764 32366
rect 27712 32302 27764 32308
rect 27724 31958 27752 32302
rect 27816 32230 27844 34954
rect 29000 34672 29052 34678
rect 29000 34614 29052 34620
rect 27988 34536 28040 34542
rect 27988 34478 28040 34484
rect 28000 33862 28028 34478
rect 28172 34400 28224 34406
rect 28172 34342 28224 34348
rect 28264 34400 28316 34406
rect 28264 34342 28316 34348
rect 28184 34066 28212 34342
rect 28172 34060 28224 34066
rect 28172 34002 28224 34008
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 28000 33590 28028 33798
rect 27988 33584 28040 33590
rect 27988 33526 28040 33532
rect 27894 33008 27950 33017
rect 27894 32943 27950 32952
rect 27908 32910 27936 32943
rect 27896 32904 27948 32910
rect 27896 32846 27948 32852
rect 28080 32904 28132 32910
rect 28080 32846 28132 32852
rect 28092 32570 28120 32846
rect 28184 32609 28212 34002
rect 28276 33046 28304 34342
rect 28908 33924 28960 33930
rect 28908 33866 28960 33872
rect 28540 33856 28592 33862
rect 28540 33798 28592 33804
rect 28264 33040 28316 33046
rect 28264 32982 28316 32988
rect 28356 33040 28408 33046
rect 28356 32982 28408 32988
rect 28368 32745 28396 32982
rect 28552 32910 28580 33798
rect 28920 33017 28948 33866
rect 29012 33522 29040 34614
rect 29184 33924 29236 33930
rect 29184 33866 29236 33872
rect 29000 33516 29052 33522
rect 29000 33458 29052 33464
rect 29196 33454 29224 33866
rect 29184 33448 29236 33454
rect 29184 33390 29236 33396
rect 28906 33008 28962 33017
rect 29288 32978 29316 37062
rect 29748 35894 29776 37062
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 29748 35866 30144 35894
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 29368 34196 29420 34202
rect 29368 34138 29420 34144
rect 29380 33318 29408 34138
rect 29460 34128 29512 34134
rect 29460 34070 29512 34076
rect 29472 33522 29500 34070
rect 29920 33924 29972 33930
rect 29920 33866 29972 33872
rect 29932 33590 29960 33866
rect 29920 33584 29972 33590
rect 29920 33526 29972 33532
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 29644 33448 29696 33454
rect 29644 33390 29696 33396
rect 29368 33312 29420 33318
rect 29368 33254 29420 33260
rect 29656 33114 29684 33390
rect 29644 33108 29696 33114
rect 29644 33050 29696 33056
rect 28906 32943 28962 32952
rect 29184 32972 29236 32978
rect 29184 32914 29236 32920
rect 29276 32972 29328 32978
rect 29328 32932 29408 32960
rect 29276 32914 29328 32920
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28816 32904 28868 32910
rect 29000 32904 29052 32910
rect 28816 32846 28868 32852
rect 28920 32864 29000 32892
rect 28632 32836 28684 32842
rect 28632 32778 28684 32784
rect 28644 32745 28672 32778
rect 28354 32736 28410 32745
rect 28354 32671 28410 32680
rect 28630 32736 28686 32745
rect 28630 32671 28686 32680
rect 28170 32600 28226 32609
rect 28080 32564 28132 32570
rect 28170 32535 28226 32544
rect 28080 32506 28132 32512
rect 28172 32496 28224 32502
rect 28170 32464 28172 32473
rect 28224 32464 28226 32473
rect 27988 32428 28040 32434
rect 28170 32399 28226 32408
rect 27988 32370 28040 32376
rect 27804 32224 27856 32230
rect 27804 32166 27856 32172
rect 27620 31952 27672 31958
rect 27620 31894 27672 31900
rect 27712 31952 27764 31958
rect 27712 31894 27764 31900
rect 27620 31816 27672 31822
rect 27618 31784 27620 31793
rect 27672 31784 27674 31793
rect 27618 31719 27674 31728
rect 27528 31680 27580 31686
rect 27434 31648 27490 31657
rect 27528 31622 27580 31628
rect 27434 31583 27490 31592
rect 27172 31368 27384 31396
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 27068 30388 27120 30394
rect 27068 30330 27120 30336
rect 26976 29708 27028 29714
rect 26976 29650 27028 29656
rect 27080 29646 27108 30330
rect 27172 29850 27200 31368
rect 27356 31142 27384 31368
rect 27448 31142 27476 31583
rect 27540 31346 27568 31622
rect 27724 31346 27752 31894
rect 27528 31340 27580 31346
rect 27528 31282 27580 31288
rect 27712 31340 27764 31346
rect 27712 31282 27764 31288
rect 27344 31136 27396 31142
rect 27344 31078 27396 31084
rect 27436 31136 27488 31142
rect 27436 31078 27488 31084
rect 27540 30920 27568 31282
rect 27620 31204 27672 31210
rect 27620 31146 27672 31152
rect 27632 30938 27660 31146
rect 27448 30892 27568 30920
rect 27620 30932 27672 30938
rect 27342 30832 27398 30841
rect 27342 30767 27398 30776
rect 27250 30288 27306 30297
rect 27356 30258 27384 30767
rect 27448 30734 27476 30892
rect 27620 30874 27672 30880
rect 27632 30841 27660 30874
rect 27618 30832 27674 30841
rect 27528 30796 27580 30802
rect 27618 30767 27674 30776
rect 27528 30738 27580 30744
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27434 30560 27490 30569
rect 27434 30495 27490 30504
rect 27448 30394 27476 30495
rect 27436 30388 27488 30394
rect 27436 30330 27488 30336
rect 27250 30223 27306 30232
rect 27344 30252 27396 30258
rect 27160 29844 27212 29850
rect 27160 29786 27212 29792
rect 26792 29640 26844 29646
rect 26792 29582 26844 29588
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 27068 29640 27120 29646
rect 27068 29582 27120 29588
rect 26712 29464 26832 29492
rect 26804 29306 26832 29464
rect 26608 29300 26660 29306
rect 26608 29242 26660 29248
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26528 29170 26740 29186
rect 26528 29164 26752 29170
rect 26528 29158 26700 29164
rect 26700 29106 26752 29112
rect 26608 29096 26660 29102
rect 26608 29038 26660 29044
rect 26516 28960 26568 28966
rect 26436 28908 26516 28914
rect 26436 28902 26568 28908
rect 26436 28886 26556 28902
rect 26332 28484 26384 28490
rect 26332 28426 26384 28432
rect 26240 28076 26292 28082
rect 26240 28018 26292 28024
rect 26252 27878 26280 28018
rect 26344 28014 26372 28426
rect 26436 28150 26464 28886
rect 26620 28558 26648 29038
rect 26700 28756 26752 28762
rect 26700 28698 26752 28704
rect 26712 28626 26740 28698
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26516 28552 26568 28558
rect 26516 28494 26568 28500
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26528 28218 26556 28494
rect 26516 28212 26568 28218
rect 26516 28154 26568 28160
rect 26424 28144 26476 28150
rect 26424 28086 26476 28092
rect 26332 28008 26384 28014
rect 26332 27950 26384 27956
rect 26240 27872 26292 27878
rect 26240 27814 26292 27820
rect 26252 27538 26280 27814
rect 26344 27606 26372 27950
rect 26332 27600 26384 27606
rect 26332 27542 26384 27548
rect 26240 27532 26292 27538
rect 26240 27474 26292 27480
rect 26344 27418 26372 27542
rect 26252 27390 26372 27418
rect 26252 26994 26280 27390
rect 26436 27305 26464 28086
rect 26620 27690 26648 28494
rect 26528 27662 26648 27690
rect 26712 27674 26740 28562
rect 26700 27668 26752 27674
rect 26422 27296 26478 27305
rect 26422 27231 26478 27240
rect 26240 26988 26292 26994
rect 26240 26930 26292 26936
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 26238 26480 26294 26489
rect 26238 26415 26294 26424
rect 26252 26382 26280 26415
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26436 26246 26464 26930
rect 26424 26240 26476 26246
rect 26160 26200 26372 26228
rect 26068 26030 26188 26058
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 26068 25226 26096 25842
rect 26056 25220 26108 25226
rect 26056 25162 26108 25168
rect 25870 24783 25872 24792
rect 25924 24783 25926 24792
rect 25964 24812 26016 24818
rect 25872 24754 25924 24760
rect 25964 24754 26016 24760
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 25780 24200 25832 24206
rect 25780 24142 25832 24148
rect 25780 23656 25832 23662
rect 25780 23598 25832 23604
rect 25792 23118 25820 23598
rect 25884 23254 25912 24754
rect 26068 24410 26096 24754
rect 26056 24404 26108 24410
rect 26056 24346 26108 24352
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 25872 23248 25924 23254
rect 25872 23190 25924 23196
rect 25780 23112 25832 23118
rect 25780 23054 25832 23060
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 25608 22409 25636 22578
rect 25688 22500 25740 22506
rect 25688 22442 25740 22448
rect 25594 22400 25650 22409
rect 25594 22335 25650 22344
rect 25516 22222 25636 22250
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25516 20942 25544 21490
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25608 19281 25636 22222
rect 25700 20466 25728 22442
rect 25792 21894 25820 23054
rect 25884 22574 25912 23054
rect 25872 22568 25924 22574
rect 25872 22510 25924 22516
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 25792 20602 25820 20742
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25792 20466 25820 20538
rect 25976 20466 26004 24142
rect 26056 23520 26108 23526
rect 26056 23462 26108 23468
rect 26068 22098 26096 23462
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 26056 21412 26108 21418
rect 26056 21354 26108 21360
rect 26068 20874 26096 21354
rect 26056 20868 26108 20874
rect 26056 20810 26108 20816
rect 26160 20777 26188 26030
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26252 24410 26280 24618
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 26240 24132 26292 24138
rect 26240 24074 26292 24080
rect 26252 23526 26280 24074
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26344 22098 26372 26200
rect 26424 26182 26476 26188
rect 26436 25498 26464 26182
rect 26424 25492 26476 25498
rect 26424 25434 26476 25440
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 26436 24206 26464 24754
rect 26528 24410 26556 27662
rect 26700 27610 26752 27616
rect 26608 27532 26660 27538
rect 26608 27474 26660 27480
rect 26620 27334 26648 27474
rect 26608 27328 26660 27334
rect 26608 27270 26660 27276
rect 26804 26790 26832 29242
rect 26884 29096 26936 29102
rect 26884 29038 26936 29044
rect 26896 28966 26924 29038
rect 26884 28960 26936 28966
rect 26884 28902 26936 28908
rect 26974 28928 27030 28937
rect 26974 28863 27030 28872
rect 26882 28248 26938 28257
rect 26882 28183 26938 28192
rect 26896 28150 26924 28183
rect 26884 28144 26936 28150
rect 26884 28086 26936 28092
rect 26988 27985 27016 28863
rect 27080 28762 27108 29582
rect 27264 28994 27292 30223
rect 27344 30194 27396 30200
rect 27356 29646 27384 30194
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 27342 29472 27398 29481
rect 27342 29407 27398 29416
rect 27172 28966 27292 28994
rect 27068 28756 27120 28762
rect 27068 28698 27120 28704
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 26974 27976 27030 27985
rect 26974 27911 26976 27920
rect 27028 27911 27030 27920
rect 26976 27882 27028 27888
rect 27080 27878 27108 28018
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 26974 27568 27030 27577
rect 26974 27503 27030 27512
rect 26884 27328 26936 27334
rect 26884 27270 26936 27276
rect 26896 27169 26924 27270
rect 26882 27160 26938 27169
rect 26882 27095 26938 27104
rect 26792 26784 26844 26790
rect 26792 26726 26844 26732
rect 26700 26580 26752 26586
rect 26700 26522 26752 26528
rect 26608 26444 26660 26450
rect 26608 26386 26660 26392
rect 26620 25906 26648 26386
rect 26712 26382 26740 26522
rect 26700 26376 26752 26382
rect 26700 26318 26752 26324
rect 26792 26240 26844 26246
rect 26792 26182 26844 26188
rect 26608 25900 26660 25906
rect 26608 25842 26660 25848
rect 26608 24812 26660 24818
rect 26608 24754 26660 24760
rect 26620 24410 26648 24754
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26608 24404 26660 24410
rect 26608 24346 26660 24352
rect 26608 24268 26660 24274
rect 26608 24210 26660 24216
rect 26424 24200 26476 24206
rect 26476 24160 26556 24188
rect 26424 24142 26476 24148
rect 26528 24070 26556 24160
rect 26424 24064 26476 24070
rect 26424 24006 26476 24012
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 26332 22092 26384 22098
rect 26332 22034 26384 22040
rect 26240 22024 26292 22030
rect 26238 21992 26240 22001
rect 26292 21992 26294 22001
rect 26294 21950 26372 21978
rect 26238 21927 26294 21936
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26146 20768 26202 20777
rect 26146 20703 26202 20712
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 25594 19272 25650 19281
rect 25594 19207 25650 19216
rect 25594 18728 25650 18737
rect 25594 18663 25596 18672
rect 25648 18663 25650 18672
rect 25596 18634 25648 18640
rect 25504 18624 25556 18630
rect 25504 18566 25556 18572
rect 25410 18320 25466 18329
rect 25410 18255 25412 18264
rect 25464 18255 25466 18264
rect 25412 18226 25464 18232
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 25228 16788 25280 16794
rect 25228 16730 25280 16736
rect 25332 16726 25360 17138
rect 25320 16720 25372 16726
rect 25320 16662 25372 16668
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 25148 15570 25176 16594
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25240 16114 25268 16526
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25136 15564 25188 15570
rect 25136 15506 25188 15512
rect 25240 14958 25268 16050
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25056 12838 25176 12866
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25056 12238 25084 12718
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 24860 12164 24912 12170
rect 24860 12106 24912 12112
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24228 10810 24256 10950
rect 24216 10804 24268 10810
rect 24216 10746 24268 10752
rect 24320 9489 24348 11290
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24400 11076 24452 11082
rect 24400 11018 24452 11024
rect 24412 10470 24440 11018
rect 24780 10742 24808 11154
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24400 10464 24452 10470
rect 24400 10406 24452 10412
rect 24412 10266 24440 10406
rect 24490 10296 24546 10305
rect 24400 10260 24452 10266
rect 24490 10231 24492 10240
rect 24400 10202 24452 10208
rect 24544 10231 24546 10240
rect 24492 10202 24544 10208
rect 24400 9988 24452 9994
rect 24400 9930 24452 9936
rect 24306 9480 24362 9489
rect 24306 9415 24362 9424
rect 24412 9217 24440 9930
rect 24398 9208 24454 9217
rect 24398 9143 24454 9152
rect 24306 8936 24362 8945
rect 24306 8871 24362 8880
rect 24320 8022 24348 8871
rect 24412 8090 24440 9143
rect 24400 8084 24452 8090
rect 24400 8026 24452 8032
rect 24308 8016 24360 8022
rect 24308 7958 24360 7964
rect 24596 7954 24624 10610
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24780 8634 24808 10474
rect 24872 10062 24900 11018
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24216 6928 24268 6934
rect 24216 6870 24268 6876
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 24032 6384 24084 6390
rect 24032 6326 24084 6332
rect 24124 6316 24176 6322
rect 24228 6304 24256 6870
rect 24688 6458 24716 7822
rect 24964 7750 24992 12174
rect 25056 11830 25084 12174
rect 25044 11824 25096 11830
rect 25044 11766 25096 11772
rect 25148 10810 25176 12838
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 25042 10432 25098 10441
rect 25042 10367 25098 10376
rect 25056 10266 25084 10367
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 25056 9110 25084 10202
rect 25240 9654 25268 14758
rect 25332 13870 25360 15846
rect 25424 14550 25452 18022
rect 25516 17785 25544 18566
rect 25608 18290 25636 18634
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25608 18034 25636 18226
rect 25700 18154 25728 20402
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 25964 19848 26016 19854
rect 25962 19816 25964 19825
rect 26016 19816 26018 19825
rect 25962 19751 26018 19760
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25792 18426 25820 19110
rect 26068 18834 26096 19994
rect 26056 18828 26108 18834
rect 26056 18770 26108 18776
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25884 18630 25912 18702
rect 26068 18698 26096 18770
rect 26056 18692 26108 18698
rect 26056 18634 26108 18640
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25884 18170 25912 18566
rect 26068 18290 26096 18634
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26160 18193 26188 18226
rect 26146 18184 26202 18193
rect 25688 18148 25740 18154
rect 25884 18142 26096 18170
rect 25688 18090 25740 18096
rect 25608 18006 25912 18034
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 25502 17776 25558 17785
rect 25502 17711 25558 17720
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25516 15094 25544 17138
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25504 15088 25556 15094
rect 25504 15030 25556 15036
rect 25608 15042 25636 16730
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 25700 16250 25728 16526
rect 25688 16244 25740 16250
rect 25688 16186 25740 16192
rect 25412 14544 25464 14550
rect 25412 14486 25464 14492
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 25424 13734 25452 14486
rect 25516 14414 25544 15030
rect 25608 15014 25728 15042
rect 25596 14952 25648 14958
rect 25594 14920 25596 14929
rect 25648 14920 25650 14929
rect 25594 14855 25650 14864
rect 25504 14408 25556 14414
rect 25504 14350 25556 14356
rect 25596 14340 25648 14346
rect 25596 14282 25648 14288
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25608 12170 25636 14282
rect 25700 13802 25728 15014
rect 25792 14958 25820 17818
rect 25780 14952 25832 14958
rect 25780 14894 25832 14900
rect 25884 14804 25912 18006
rect 25964 17060 26016 17066
rect 25964 17002 26016 17008
rect 25792 14776 25912 14804
rect 25792 14385 25820 14776
rect 25976 14550 26004 17002
rect 26068 16114 26096 18142
rect 26146 18119 26202 18128
rect 26252 16794 26280 21830
rect 26344 21690 26372 21950
rect 26436 21894 26464 24006
rect 26528 23730 26556 24006
rect 26516 23724 26568 23730
rect 26516 23666 26568 23672
rect 26620 23594 26648 24210
rect 26608 23588 26660 23594
rect 26608 23530 26660 23536
rect 26516 23248 26568 23254
rect 26516 23190 26568 23196
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26332 21684 26384 21690
rect 26332 21626 26384 21632
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 26344 20466 26372 21082
rect 26528 20641 26556 23190
rect 26514 20632 26570 20641
rect 26514 20567 26570 20576
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26344 17270 26372 20402
rect 26436 19990 26464 20402
rect 26528 20330 26556 20402
rect 26516 20324 26568 20330
rect 26516 20266 26568 20272
rect 26424 19984 26476 19990
rect 26424 19926 26476 19932
rect 26528 19922 26556 20266
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26528 19334 26556 19858
rect 26436 19306 26556 19334
rect 26332 17264 26384 17270
rect 26332 17206 26384 17212
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26332 16788 26384 16794
rect 26332 16730 26384 16736
rect 26344 16522 26372 16730
rect 26332 16516 26384 16522
rect 26332 16458 26384 16464
rect 26344 16182 26372 16458
rect 26332 16176 26384 16182
rect 26332 16118 26384 16124
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26160 14618 26188 15982
rect 26240 15632 26292 15638
rect 26240 15574 26292 15580
rect 26252 15026 26280 15574
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 25964 14544 26016 14550
rect 25964 14486 26016 14492
rect 25872 14408 25924 14414
rect 25778 14376 25834 14385
rect 25872 14350 25924 14356
rect 25778 14311 25834 14320
rect 25688 13796 25740 13802
rect 25688 13738 25740 13744
rect 25688 12300 25740 12306
rect 25688 12242 25740 12248
rect 25596 12164 25648 12170
rect 25596 12106 25648 12112
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 25332 11694 25360 12038
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25332 11082 25360 11630
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25318 10704 25374 10713
rect 25318 10639 25374 10648
rect 25332 10062 25360 10639
rect 25516 10266 25544 11494
rect 25608 10441 25636 12106
rect 25700 11121 25728 12242
rect 25686 11112 25742 11121
rect 25686 11047 25742 11056
rect 25792 10810 25820 14311
rect 25884 14074 25912 14350
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 25976 12442 26004 14486
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 14074 26188 14214
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26054 12472 26110 12481
rect 25964 12436 26016 12442
rect 26054 12407 26110 12416
rect 25964 12378 26016 12384
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25594 10432 25650 10441
rect 25594 10367 25650 10376
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 25424 9761 25452 9998
rect 25410 9752 25466 9761
rect 25410 9687 25466 9696
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25044 9104 25096 9110
rect 25044 9046 25096 9052
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 25332 7886 25360 8774
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25424 8498 25452 8570
rect 25412 8492 25464 8498
rect 25792 8480 25820 10202
rect 25884 9382 25912 12174
rect 25964 12164 26016 12170
rect 25964 12106 26016 12112
rect 25976 10062 26004 12106
rect 26068 10130 26096 12407
rect 26252 10470 26280 14962
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26240 10464 26292 10470
rect 26240 10406 26292 10412
rect 26238 10160 26294 10169
rect 26056 10124 26108 10130
rect 26238 10095 26294 10104
rect 26056 10066 26108 10072
rect 26252 10062 26280 10095
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 26056 9988 26108 9994
rect 26056 9930 26108 9936
rect 26068 9586 26096 9930
rect 26344 9722 26372 13806
rect 26436 13734 26464 19306
rect 26620 19145 26648 23530
rect 26804 23474 26832 26182
rect 26896 24138 26924 27095
rect 26988 26450 27016 27503
rect 27080 27470 27108 27814
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 26976 26444 27028 26450
rect 26976 26386 27028 26392
rect 27080 26330 27108 27406
rect 27172 27169 27200 28966
rect 27250 28792 27306 28801
rect 27356 28778 27384 29407
rect 27306 28750 27384 28778
rect 27250 28727 27306 28736
rect 27448 28676 27476 29990
rect 27540 29714 27568 30738
rect 27620 30728 27672 30734
rect 27618 30696 27620 30705
rect 27672 30696 27674 30705
rect 27724 30666 27752 31282
rect 27618 30631 27674 30640
rect 27712 30660 27764 30666
rect 27712 30602 27764 30608
rect 27620 30592 27672 30598
rect 27620 30534 27672 30540
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27528 29572 27580 29578
rect 27528 29514 27580 29520
rect 27540 29170 27568 29514
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27356 28648 27476 28676
rect 27356 28490 27384 28648
rect 27632 28642 27660 30534
rect 27712 30388 27764 30394
rect 27712 30330 27764 30336
rect 27724 30297 27752 30330
rect 27710 30288 27766 30297
rect 27710 30223 27766 30232
rect 27816 29889 27844 32166
rect 27896 31476 27948 31482
rect 27896 31418 27948 31424
rect 27908 31210 27936 31418
rect 27896 31204 27948 31210
rect 27896 31146 27948 31152
rect 27908 30734 27936 31146
rect 27896 30728 27948 30734
rect 28000 30705 28028 32370
rect 28356 32360 28408 32366
rect 28262 32328 28318 32337
rect 28356 32302 28408 32308
rect 28262 32263 28318 32272
rect 28172 32224 28224 32230
rect 28172 32166 28224 32172
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 28092 31385 28120 31758
rect 28078 31376 28134 31385
rect 28078 31311 28134 31320
rect 28080 31204 28132 31210
rect 28080 31146 28132 31152
rect 28092 31113 28120 31146
rect 28078 31104 28134 31113
rect 28078 31039 28134 31048
rect 28092 30938 28120 31039
rect 28080 30932 28132 30938
rect 28080 30874 28132 30880
rect 28080 30728 28132 30734
rect 27896 30670 27948 30676
rect 27986 30696 28042 30705
rect 28080 30670 28132 30676
rect 27986 30631 28042 30640
rect 28000 30394 28028 30631
rect 27988 30388 28040 30394
rect 27988 30330 28040 30336
rect 27896 30116 27948 30122
rect 27896 30058 27948 30064
rect 27802 29880 27858 29889
rect 27802 29815 27858 29824
rect 27710 29744 27766 29753
rect 27710 29679 27766 29688
rect 27724 29646 27752 29679
rect 27712 29640 27764 29646
rect 27712 29582 27764 29588
rect 27710 29472 27766 29481
rect 27710 29407 27766 29416
rect 27724 29034 27752 29407
rect 27804 29164 27856 29170
rect 27804 29106 27856 29112
rect 27712 29028 27764 29034
rect 27712 28970 27764 28976
rect 27712 28756 27764 28762
rect 27712 28698 27764 28704
rect 27540 28626 27660 28642
rect 27528 28620 27660 28626
rect 27580 28614 27660 28620
rect 27528 28562 27580 28568
rect 27252 28484 27304 28490
rect 27252 28426 27304 28432
rect 27344 28484 27396 28490
rect 27344 28426 27396 28432
rect 27264 27674 27292 28426
rect 27356 28218 27384 28426
rect 27540 28370 27568 28562
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27471 28342 27568 28370
rect 27471 28234 27499 28342
rect 27344 28212 27396 28218
rect 27344 28154 27396 28160
rect 27448 28206 27499 28234
rect 27632 28218 27660 28494
rect 27724 28218 27752 28698
rect 27528 28212 27580 28218
rect 27344 27872 27396 27878
rect 27344 27814 27396 27820
rect 27356 27713 27384 27814
rect 27342 27704 27398 27713
rect 27252 27668 27304 27674
rect 27342 27639 27398 27648
rect 27252 27610 27304 27616
rect 27356 27538 27384 27639
rect 27344 27532 27396 27538
rect 27344 27474 27396 27480
rect 27252 27396 27304 27402
rect 27252 27338 27304 27344
rect 27264 27305 27292 27338
rect 27250 27296 27306 27305
rect 27250 27231 27306 27240
rect 27158 27160 27214 27169
rect 27158 27095 27214 27104
rect 27160 27056 27212 27062
rect 27160 26998 27212 27004
rect 27172 26897 27200 26998
rect 27158 26888 27214 26897
rect 27158 26823 27214 26832
rect 27160 26784 27212 26790
rect 27160 26726 27212 26732
rect 26988 26314 27108 26330
rect 26976 26308 27108 26314
rect 27028 26302 27108 26308
rect 26976 26250 27028 26256
rect 27172 26228 27200 26726
rect 27264 26246 27292 27231
rect 27448 26994 27476 28206
rect 27528 28154 27580 28160
rect 27620 28212 27672 28218
rect 27620 28154 27672 28160
rect 27712 28212 27764 28218
rect 27712 28154 27764 28160
rect 27540 27470 27568 28154
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27618 27432 27674 27441
rect 27540 26994 27568 27406
rect 27618 27367 27674 27376
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27528 26988 27580 26994
rect 27528 26930 27580 26936
rect 27632 26926 27660 27367
rect 27816 27334 27844 29106
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27620 26920 27672 26926
rect 27620 26862 27672 26868
rect 27908 26382 27936 30058
rect 28000 29617 28028 30330
rect 28092 30326 28120 30670
rect 28184 30598 28212 32166
rect 28276 31822 28304 32263
rect 28368 31958 28396 32302
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28644 32026 28672 32166
rect 28632 32020 28684 32026
rect 28632 31962 28684 31968
rect 28356 31952 28408 31958
rect 28356 31894 28408 31900
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28276 31657 28304 31758
rect 28262 31648 28318 31657
rect 28262 31583 28318 31592
rect 28262 31376 28318 31385
rect 28262 31311 28318 31320
rect 28276 31210 28304 31311
rect 28264 31204 28316 31210
rect 28264 31146 28316 31152
rect 28172 30592 28224 30598
rect 28172 30534 28224 30540
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 28184 30190 28212 30534
rect 28264 30320 28316 30326
rect 28262 30288 28264 30297
rect 28316 30288 28318 30297
rect 28262 30223 28318 30232
rect 28172 30184 28224 30190
rect 28172 30126 28224 30132
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28080 30116 28132 30122
rect 28080 30058 28132 30064
rect 28092 30025 28120 30058
rect 28078 30016 28134 30025
rect 28078 29951 28134 29960
rect 28078 29880 28134 29889
rect 28078 29815 28134 29824
rect 27986 29608 28042 29617
rect 27986 29543 28042 29552
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 28000 26382 28028 29446
rect 28092 29084 28120 29815
rect 28276 29730 28304 30126
rect 28184 29702 28304 29730
rect 28184 29510 28212 29702
rect 28264 29640 28316 29646
rect 28262 29608 28264 29617
rect 28316 29608 28318 29617
rect 28262 29543 28318 29552
rect 28172 29504 28224 29510
rect 28172 29446 28224 29452
rect 28184 29238 28212 29446
rect 28172 29232 28224 29238
rect 28172 29174 28224 29180
rect 28262 29200 28318 29209
rect 28262 29135 28264 29144
rect 28316 29135 28318 29144
rect 28264 29106 28316 29112
rect 28092 29056 28212 29084
rect 28080 28960 28132 28966
rect 28080 28902 28132 28908
rect 28092 28694 28120 28902
rect 28080 28688 28132 28694
rect 28080 28630 28132 28636
rect 27436 26376 27488 26382
rect 27356 26336 27436 26364
rect 27080 26200 27200 26228
rect 27252 26240 27304 26246
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26884 24132 26936 24138
rect 26884 24074 26936 24080
rect 26896 23594 26924 24074
rect 26884 23588 26936 23594
rect 26884 23530 26936 23536
rect 26804 23446 26924 23474
rect 26792 20800 26844 20806
rect 26792 20742 26844 20748
rect 26804 20534 26832 20742
rect 26792 20528 26844 20534
rect 26792 20470 26844 20476
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26700 19236 26752 19242
rect 26700 19178 26752 19184
rect 26606 19136 26662 19145
rect 26606 19071 26662 19080
rect 26620 18170 26648 19071
rect 26712 18873 26740 19178
rect 26698 18864 26754 18873
rect 26698 18799 26754 18808
rect 26700 18760 26752 18766
rect 26700 18702 26752 18708
rect 26712 18426 26740 18702
rect 26700 18420 26752 18426
rect 26700 18362 26752 18368
rect 26620 18142 26740 18170
rect 26514 16688 26570 16697
rect 26514 16623 26570 16632
rect 26528 16590 26556 16623
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26620 14278 26648 16526
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26424 13728 26476 13734
rect 26476 13688 26556 13716
rect 26424 13670 26476 13676
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26436 12646 26464 13466
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26332 9716 26384 9722
rect 26332 9658 26384 9664
rect 26436 9654 26464 12582
rect 26528 11218 26556 13688
rect 26620 12714 26648 14214
rect 26712 13938 26740 18142
rect 26804 16590 26832 19654
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 26608 12708 26660 12714
rect 26608 12650 26660 12656
rect 26608 12368 26660 12374
rect 26608 12310 26660 12316
rect 26620 11354 26648 12310
rect 26698 11928 26754 11937
rect 26698 11863 26700 11872
rect 26752 11863 26754 11872
rect 26700 11834 26752 11840
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26516 9988 26568 9994
rect 26516 9930 26568 9936
rect 26424 9648 26476 9654
rect 26238 9616 26294 9625
rect 26056 9580 26108 9586
rect 26424 9590 26476 9596
rect 26238 9551 26294 9560
rect 26056 9522 26108 9528
rect 26068 9489 26096 9522
rect 26054 9480 26110 9489
rect 26054 9415 26110 9424
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25884 9178 25912 9318
rect 26146 9208 26202 9217
rect 25872 9172 25924 9178
rect 26146 9143 26202 9152
rect 25872 9114 25924 9120
rect 26160 8498 26188 9143
rect 26252 8514 26280 9551
rect 26148 8492 26200 8498
rect 25792 8452 25912 8480
rect 25412 8434 25464 8440
rect 25688 8424 25740 8430
rect 25740 8384 25820 8412
rect 25688 8366 25740 8372
rect 25792 8294 25820 8384
rect 25688 8288 25740 8294
rect 25502 8256 25558 8265
rect 25688 8230 25740 8236
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25502 8191 25558 8200
rect 25516 7886 25544 8191
rect 25700 8090 25728 8230
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25792 7886 25820 8230
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 25504 7880 25556 7886
rect 25504 7822 25556 7828
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 25228 7812 25280 7818
rect 25228 7754 25280 7760
rect 25412 7812 25464 7818
rect 25412 7754 25464 7760
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24952 7744 25004 7750
rect 24952 7686 25004 7692
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 24872 7290 24900 7686
rect 24964 7546 24992 7686
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 25056 7478 25084 7686
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 25240 7410 25268 7754
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25424 7342 25452 7754
rect 25700 7478 25728 7822
rect 25688 7472 25740 7478
rect 25688 7414 25740 7420
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25412 7336 25464 7342
rect 24950 7304 25006 7313
rect 24872 7262 24950 7290
rect 25412 7278 25464 7284
rect 24950 7239 24952 7248
rect 25004 7239 25006 7248
rect 24952 7210 25004 7216
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 25044 6384 25096 6390
rect 25044 6326 25096 6332
rect 24176 6276 24256 6304
rect 24676 6316 24728 6322
rect 24124 6258 24176 6264
rect 24676 6258 24728 6264
rect 23940 5568 23992 5574
rect 23940 5510 23992 5516
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 22296 3233 22324 3402
rect 22664 3398 22692 4626
rect 23940 4616 23992 4622
rect 23846 4584 23902 4593
rect 23940 4558 23992 4564
rect 23846 4519 23848 4528
rect 23900 4519 23902 4528
rect 23848 4490 23900 4496
rect 23570 4176 23626 4185
rect 23570 4111 23572 4120
rect 23624 4111 23626 4120
rect 23572 4082 23624 4088
rect 23584 3534 23612 4082
rect 23860 3602 23888 4490
rect 23952 4049 23980 4558
rect 23938 4040 23994 4049
rect 23938 3975 23994 3984
rect 23952 3942 23980 3975
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 24044 3738 24072 5170
rect 24136 4146 24164 6258
rect 24688 6118 24716 6258
rect 24584 6112 24636 6118
rect 24584 6054 24636 6060
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24596 5914 24624 6054
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24596 5710 24624 5850
rect 24688 5778 24716 6054
rect 25056 5778 25084 6326
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 25044 5772 25096 5778
rect 25044 5714 25096 5720
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24308 5364 24360 5370
rect 24308 5306 24360 5312
rect 24320 4214 24348 5306
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24412 4214 24440 4762
rect 24308 4208 24360 4214
rect 24308 4150 24360 4156
rect 24400 4208 24452 4214
rect 24400 4150 24452 4156
rect 25332 4146 25360 6938
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 25424 6254 25452 6598
rect 25516 6322 25544 7142
rect 25608 6322 25636 7346
rect 25688 7336 25740 7342
rect 25688 7278 25740 7284
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 25596 6316 25648 6322
rect 25596 6258 25648 6264
rect 25412 6248 25464 6254
rect 25412 6190 25464 6196
rect 25516 5914 25544 6258
rect 25700 6118 25728 7278
rect 25792 6934 25820 7822
rect 25884 7002 25912 8452
rect 26252 8486 26372 8514
rect 26148 8434 26200 8440
rect 26056 8424 26108 8430
rect 26056 8366 26108 8372
rect 26068 8106 26096 8366
rect 26068 8078 26280 8106
rect 26148 8016 26200 8022
rect 26054 7984 26110 7993
rect 26148 7958 26200 7964
rect 26054 7919 26110 7928
rect 26068 7886 26096 7919
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 26160 7410 26188 7958
rect 26252 7546 26280 8078
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 25872 6996 25924 7002
rect 25872 6938 25924 6944
rect 25780 6928 25832 6934
rect 25780 6870 25832 6876
rect 25872 6860 25924 6866
rect 25872 6802 25924 6808
rect 25884 6458 25912 6802
rect 25872 6452 25924 6458
rect 25872 6394 25924 6400
rect 26056 6384 26108 6390
rect 26056 6326 26108 6332
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25504 5908 25556 5914
rect 25504 5850 25556 5856
rect 26068 5681 26096 6326
rect 26160 6186 26188 7346
rect 26344 6866 26372 8486
rect 26436 7002 26464 9590
rect 26528 7886 26556 9930
rect 26620 8634 26648 10406
rect 26712 9194 26740 11698
rect 26804 11354 26832 16526
rect 26896 14482 26924 23446
rect 26988 21962 27016 24346
rect 27080 23050 27108 26200
rect 27252 26182 27304 26188
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 27158 24712 27214 24721
rect 27158 24647 27160 24656
rect 27212 24647 27214 24656
rect 27160 24618 27212 24624
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 27068 23044 27120 23050
rect 27068 22986 27120 22992
rect 27068 22092 27120 22098
rect 27172 22094 27200 24142
rect 27264 23866 27292 24754
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 27172 22066 27292 22094
rect 27068 22034 27120 22040
rect 26976 21956 27028 21962
rect 26976 21898 27028 21904
rect 26988 21146 27016 21898
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 27080 20890 27108 22034
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 26988 20862 27108 20890
rect 26988 17746 27016 20862
rect 27066 20496 27122 20505
rect 27066 20431 27068 20440
rect 27120 20431 27122 20440
rect 27068 20402 27120 20408
rect 27068 18760 27120 18766
rect 27068 18702 27120 18708
rect 27080 18358 27108 18702
rect 27068 18352 27120 18358
rect 27068 18294 27120 18300
rect 26976 17740 27028 17746
rect 26976 17682 27028 17688
rect 27172 17082 27200 21966
rect 27264 21010 27292 22066
rect 27252 21004 27304 21010
rect 27252 20946 27304 20952
rect 27264 20874 27292 20946
rect 27252 20868 27304 20874
rect 27252 20810 27304 20816
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27264 20058 27292 20402
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 27356 18290 27384 26336
rect 27436 26318 27488 26324
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 27988 26376 28040 26382
rect 27988 26318 28040 26324
rect 27620 26308 27672 26314
rect 27620 26250 27672 26256
rect 27632 25906 27660 26250
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 27528 24812 27580 24818
rect 27528 24754 27580 24760
rect 27540 24342 27568 24754
rect 27724 24682 27752 26318
rect 27988 24948 28040 24954
rect 27988 24890 28040 24896
rect 28000 24818 28028 24890
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 27896 24608 27948 24614
rect 27896 24550 27948 24556
rect 27908 24410 27936 24550
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 27528 24336 27580 24342
rect 27528 24278 27580 24284
rect 27816 24274 27844 24346
rect 27804 24268 27856 24274
rect 27804 24210 27856 24216
rect 27528 24200 27580 24206
rect 27526 24168 27528 24177
rect 27580 24168 27582 24177
rect 27526 24103 27582 24112
rect 27620 24132 27672 24138
rect 27620 24074 27672 24080
rect 27632 23322 27660 24074
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27632 22438 27660 23054
rect 28092 22642 28120 28630
rect 28184 24138 28212 29056
rect 28262 28792 28318 28801
rect 28262 28727 28264 28736
rect 28316 28727 28318 28736
rect 28264 28698 28316 28704
rect 28264 28552 28316 28558
rect 28262 28520 28264 28529
rect 28316 28520 28318 28529
rect 28262 28455 28318 28464
rect 28264 28144 28316 28150
rect 28264 28086 28316 28092
rect 28276 27169 28304 28086
rect 28262 27160 28318 27169
rect 28262 27095 28318 27104
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 28276 24818 28304 25094
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28276 24206 28304 24550
rect 28264 24200 28316 24206
rect 28264 24142 28316 24148
rect 28172 24132 28224 24138
rect 28172 24074 28224 24080
rect 28276 23662 28304 24142
rect 28368 23798 28396 31894
rect 28540 31884 28592 31890
rect 28540 31826 28592 31832
rect 28552 31754 28580 31826
rect 28828 31822 28856 32846
rect 28920 31890 28948 32864
rect 29000 32846 29052 32852
rect 29196 32570 29224 32914
rect 29184 32564 29236 32570
rect 29184 32506 29236 32512
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 28908 31884 28960 31890
rect 28908 31826 28960 31832
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28448 31748 28500 31754
rect 28552 31726 28672 31754
rect 28448 31690 28500 31696
rect 28460 30258 28488 31690
rect 28644 31346 28672 31726
rect 28736 31634 28764 31758
rect 28816 31680 28868 31686
rect 28814 31648 28816 31657
rect 28868 31648 28870 31657
rect 28736 31606 28814 31634
rect 28736 31414 28764 31606
rect 28814 31583 28870 31592
rect 28724 31408 28776 31414
rect 28724 31350 28776 31356
rect 28632 31340 28684 31346
rect 28632 31282 28684 31288
rect 28908 31340 28960 31346
rect 28908 31282 28960 31288
rect 28538 30968 28594 30977
rect 28538 30903 28594 30912
rect 28552 30802 28580 30903
rect 28920 30870 28948 31282
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 28908 30864 28960 30870
rect 28722 30832 28778 30841
rect 28540 30796 28592 30802
rect 28908 30806 28960 30812
rect 28722 30767 28778 30776
rect 28540 30738 28592 30744
rect 28448 30252 28500 30258
rect 28448 30194 28500 30200
rect 28460 29850 28488 30194
rect 28552 30054 28580 30738
rect 28736 30734 28764 30767
rect 28724 30728 28776 30734
rect 28724 30670 28776 30676
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28540 30048 28592 30054
rect 28540 29990 28592 29996
rect 28448 29844 28500 29850
rect 28448 29786 28500 29792
rect 28540 29776 28592 29782
rect 28446 29744 28502 29753
rect 28540 29718 28592 29724
rect 28446 29679 28502 29688
rect 28460 29646 28488 29679
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 28448 29028 28500 29034
rect 28448 28970 28500 28976
rect 28460 28937 28488 28970
rect 28552 28966 28580 29718
rect 28540 28960 28592 28966
rect 28446 28928 28502 28937
rect 28540 28902 28592 28908
rect 28446 28863 28502 28872
rect 28446 28792 28502 28801
rect 28446 28727 28502 28736
rect 28460 28422 28488 28727
rect 28448 28416 28500 28422
rect 28448 28358 28500 28364
rect 28460 28082 28488 28358
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28552 28014 28580 28902
rect 28644 28694 28672 30602
rect 28736 30258 28764 30670
rect 28816 30592 28868 30598
rect 28816 30534 28868 30540
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28632 28688 28684 28694
rect 28632 28630 28684 28636
rect 28736 28558 28764 30194
rect 28828 30036 28856 30534
rect 28920 30297 28948 30806
rect 29012 30802 29040 31078
rect 29000 30796 29052 30802
rect 29000 30738 29052 30744
rect 28906 30288 28962 30297
rect 28906 30223 28908 30232
rect 28960 30223 28962 30232
rect 29000 30252 29052 30258
rect 28908 30194 28960 30200
rect 29000 30194 29052 30200
rect 28908 30048 28960 30054
rect 28828 30008 28908 30036
rect 28908 29990 28960 29996
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 28920 29714 28948 29786
rect 29012 29782 29040 30194
rect 29104 29782 29132 32370
rect 29196 31906 29224 32506
rect 29276 32428 29328 32434
rect 29276 32370 29328 32376
rect 29288 32026 29316 32370
rect 29276 32020 29328 32026
rect 29276 31962 29328 31968
rect 29196 31878 29316 31906
rect 29182 31784 29238 31793
rect 29182 31719 29238 31728
rect 29196 31414 29224 31719
rect 29184 31408 29236 31414
rect 29184 31350 29236 31356
rect 29184 30184 29236 30190
rect 29182 30152 29184 30161
rect 29236 30152 29238 30161
rect 29182 30087 29238 30096
rect 29184 29844 29236 29850
rect 29184 29786 29236 29792
rect 29000 29776 29052 29782
rect 29000 29718 29052 29724
rect 29092 29776 29144 29782
rect 29092 29718 29144 29724
rect 28908 29708 28960 29714
rect 28908 29650 28960 29656
rect 28816 29504 28868 29510
rect 28816 29446 28868 29452
rect 28828 28626 28856 29446
rect 29012 29170 29040 29718
rect 29196 29306 29224 29786
rect 29184 29300 29236 29306
rect 29184 29242 29236 29248
rect 29000 29164 29052 29170
rect 29000 29106 29052 29112
rect 28908 28688 28960 28694
rect 28908 28630 28960 28636
rect 28816 28620 28868 28626
rect 28816 28562 28868 28568
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28632 28484 28684 28490
rect 28632 28426 28684 28432
rect 28540 28008 28592 28014
rect 28540 27950 28592 27956
rect 28448 26784 28500 26790
rect 28448 26726 28500 26732
rect 28460 26382 28488 26726
rect 28448 26376 28500 26382
rect 28448 26318 28500 26324
rect 28356 23792 28408 23798
rect 28356 23734 28408 23740
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 28276 23118 28304 23598
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28172 23044 28224 23050
rect 28172 22986 28224 22992
rect 28080 22636 28132 22642
rect 28080 22578 28132 22584
rect 27804 22568 27856 22574
rect 27804 22510 27856 22516
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27632 22098 27660 22374
rect 27620 22092 27672 22098
rect 27620 22034 27672 22040
rect 27632 18766 27660 22034
rect 27816 21962 27844 22510
rect 27804 21956 27856 21962
rect 27804 21898 27856 21904
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27724 21350 27752 21830
rect 27712 21344 27764 21350
rect 27712 21286 27764 21292
rect 27724 20806 27752 21286
rect 27988 20936 28040 20942
rect 27988 20878 28040 20884
rect 27712 20800 27764 20806
rect 28000 20777 28028 20878
rect 27712 20742 27764 20748
rect 27986 20768 28042 20777
rect 27986 20703 28042 20712
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27436 18692 27488 18698
rect 27436 18634 27488 18640
rect 27448 18329 27476 18634
rect 27540 18578 27568 18702
rect 27540 18550 27660 18578
rect 27632 18426 27660 18550
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 27434 18320 27490 18329
rect 27344 18284 27396 18290
rect 27434 18255 27490 18264
rect 27528 18284 27580 18290
rect 27344 18226 27396 18232
rect 27528 18226 27580 18232
rect 27356 17202 27384 18226
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27172 17054 27384 17082
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 26974 16824 27030 16833
rect 26974 16759 27030 16768
rect 26988 16590 27016 16759
rect 27160 16720 27212 16726
rect 27080 16680 27160 16708
rect 26976 16584 27028 16590
rect 26976 16526 27028 16532
rect 27080 15348 27108 16680
rect 27160 16662 27212 16668
rect 26988 15320 27108 15348
rect 26988 15162 27016 15320
rect 26976 15156 27028 15162
rect 26976 15098 27028 15104
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26988 14414 27016 15098
rect 27264 15026 27292 16934
rect 27356 15434 27384 17054
rect 27448 16726 27476 17614
rect 27436 16720 27488 16726
rect 27436 16662 27488 16668
rect 27436 16584 27488 16590
rect 27436 16526 27488 16532
rect 27344 15428 27396 15434
rect 27344 15370 27396 15376
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27250 14920 27306 14929
rect 27448 14906 27476 16526
rect 27250 14855 27306 14864
rect 27356 14878 27476 14906
rect 27160 14544 27212 14550
rect 27160 14486 27212 14492
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26792 11212 26844 11218
rect 26792 11154 26844 11160
rect 26804 9625 26832 11154
rect 26790 9616 26846 9625
rect 26790 9551 26846 9560
rect 26792 9512 26844 9518
rect 26792 9454 26844 9460
rect 26804 9353 26832 9454
rect 26790 9344 26846 9353
rect 26790 9279 26846 9288
rect 26712 9166 26832 9194
rect 26700 8900 26752 8906
rect 26700 8842 26752 8848
rect 26712 8809 26740 8842
rect 26698 8800 26754 8809
rect 26698 8735 26754 8744
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 26528 7206 26556 7822
rect 26620 7818 26648 8570
rect 26698 8528 26754 8537
rect 26698 8463 26700 8472
rect 26752 8463 26754 8472
rect 26700 8434 26752 8440
rect 26804 7993 26832 9166
rect 26896 9081 26924 12174
rect 26988 11880 27016 13126
rect 27080 12306 27108 14282
rect 27172 14006 27200 14486
rect 27264 14414 27292 14855
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 27160 14000 27212 14006
rect 27160 13942 27212 13948
rect 27264 13841 27292 14350
rect 27250 13832 27306 13841
rect 27250 13767 27306 13776
rect 27356 13190 27384 14878
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27448 14618 27476 14758
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27540 14498 27568 18226
rect 27620 17196 27672 17202
rect 27620 17138 27672 17144
rect 27632 17105 27660 17138
rect 27618 17096 27674 17105
rect 27618 17031 27674 17040
rect 27632 16794 27660 17031
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27632 15910 27660 16594
rect 27620 15904 27672 15910
rect 27620 15846 27672 15852
rect 27618 15328 27674 15337
rect 27618 15263 27674 15272
rect 27448 14470 27568 14498
rect 27344 13184 27396 13190
rect 27344 13126 27396 13132
rect 27068 12300 27120 12306
rect 27068 12242 27120 12248
rect 26988 11852 27384 11880
rect 27250 11792 27306 11801
rect 27160 11756 27212 11762
rect 27250 11727 27252 11736
rect 27160 11698 27212 11704
rect 27304 11727 27306 11736
rect 27252 11698 27304 11704
rect 27172 11082 27200 11698
rect 27252 11280 27304 11286
rect 27252 11222 27304 11228
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 26988 10062 27016 10202
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 27068 10056 27120 10062
rect 27068 9998 27120 10004
rect 27080 9722 27108 9998
rect 27068 9716 27120 9722
rect 27068 9658 27120 9664
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 26882 9072 26938 9081
rect 26882 9007 26938 9016
rect 26988 8956 27016 9522
rect 27080 9450 27108 9658
rect 27172 9586 27200 11018
rect 27264 10130 27292 11222
rect 27252 10124 27304 10130
rect 27252 10066 27304 10072
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 27252 9580 27304 9586
rect 27252 9522 27304 9528
rect 27068 9444 27120 9450
rect 27068 9386 27120 9392
rect 27068 8968 27120 8974
rect 26988 8936 27068 8956
rect 27120 8936 27122 8945
rect 26988 8928 27066 8936
rect 27066 8871 27122 8880
rect 26974 8256 27030 8265
rect 26974 8191 27030 8200
rect 26988 8090 27016 8191
rect 26976 8084 27028 8090
rect 26976 8026 27028 8032
rect 26790 7984 26846 7993
rect 26790 7919 26846 7928
rect 26976 7948 27028 7954
rect 26608 7812 26660 7818
rect 26608 7754 26660 7760
rect 26804 7750 26832 7919
rect 26976 7890 27028 7896
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 26988 7342 27016 7890
rect 26976 7336 27028 7342
rect 26976 7278 27028 7284
rect 26516 7200 26568 7206
rect 26516 7142 26568 7148
rect 26424 6996 26476 7002
rect 26424 6938 26476 6944
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26148 6180 26200 6186
rect 26148 6122 26200 6128
rect 26160 5710 26188 6122
rect 26252 6118 26280 6598
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 26148 5704 26200 5710
rect 26054 5672 26110 5681
rect 26148 5646 26200 5652
rect 26054 5607 26110 5616
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24688 3602 24716 3878
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22282 3224 22338 3233
rect 22282 3159 22338 3168
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22560 2848 22612 2854
rect 22020 2774 22140 2802
rect 22560 2790 22612 2796
rect 21836 2746 21956 2774
rect 21836 2446 21864 2746
rect 22112 2514 22140 2774
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 21928 800 21956 2382
rect 22572 800 22600 2790
rect 22664 2446 22692 3334
rect 23584 3126 23612 3470
rect 25424 3466 25452 4762
rect 26068 4146 26096 5607
rect 26344 5574 26372 6802
rect 26528 6118 26556 7142
rect 26884 6724 26936 6730
rect 26884 6666 26936 6672
rect 26792 6180 26844 6186
rect 26792 6122 26844 6128
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 26804 5846 26832 6122
rect 26792 5840 26844 5846
rect 26792 5782 26844 5788
rect 26332 5568 26384 5574
rect 26332 5510 26384 5516
rect 26896 5234 26924 6666
rect 26988 5710 27016 7278
rect 27068 7200 27120 7206
rect 27068 7142 27120 7148
rect 27080 6662 27108 7142
rect 27068 6656 27120 6662
rect 27068 6598 27120 6604
rect 27172 6202 27200 9522
rect 27264 8090 27292 9522
rect 27356 9382 27384 11852
rect 27448 11540 27476 14470
rect 27632 14362 27660 15263
rect 27724 15026 27752 20198
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 27816 19446 27844 19790
rect 27804 19440 27856 19446
rect 27804 19382 27856 19388
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27908 18426 27936 19314
rect 27988 19168 28040 19174
rect 27988 19110 28040 19116
rect 28000 18766 28028 19110
rect 27988 18760 28040 18766
rect 27988 18702 28040 18708
rect 27896 18420 27948 18426
rect 27896 18362 27948 18368
rect 27804 18284 27856 18290
rect 28000 18272 28028 18702
rect 27856 18244 28028 18272
rect 27804 18226 27856 18232
rect 27816 17202 27844 18226
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 27710 14512 27766 14521
rect 27710 14447 27766 14456
rect 27724 14414 27752 14447
rect 27540 14346 27660 14362
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27528 14340 27660 14346
rect 27580 14334 27660 14340
rect 27528 14282 27580 14288
rect 27618 14240 27674 14249
rect 27618 14175 27674 14184
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27540 12374 27568 13806
rect 27632 12442 27660 14175
rect 27816 14006 27844 17138
rect 28000 16454 28028 17138
rect 27988 16448 28040 16454
rect 27988 16390 28040 16396
rect 27894 16144 27950 16153
rect 28092 16114 28120 22578
rect 28184 22545 28212 22986
rect 28170 22536 28226 22545
rect 28170 22471 28226 22480
rect 28172 22024 28224 22030
rect 28172 21966 28224 21972
rect 28184 21894 28212 21966
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 28184 20874 28212 21830
rect 28368 20942 28396 23734
rect 28460 21622 28488 26318
rect 28552 23730 28580 27950
rect 28644 27577 28672 28426
rect 28814 27976 28870 27985
rect 28814 27911 28870 27920
rect 28828 27606 28856 27911
rect 28816 27600 28868 27606
rect 28630 27568 28686 27577
rect 28816 27542 28868 27548
rect 28630 27503 28686 27512
rect 28828 26586 28856 27542
rect 28816 26580 28868 26586
rect 28816 26522 28868 26528
rect 28632 25832 28684 25838
rect 28632 25774 28684 25780
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28540 21956 28592 21962
rect 28540 21898 28592 21904
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 28552 21418 28580 21898
rect 28540 21412 28592 21418
rect 28540 21354 28592 21360
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28264 20868 28316 20874
rect 28264 20810 28316 20816
rect 28184 20602 28212 20810
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28184 19854 28212 20538
rect 28276 20505 28304 20810
rect 28356 20800 28408 20806
rect 28356 20742 28408 20748
rect 28262 20496 28318 20505
rect 28262 20431 28318 20440
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 28184 19174 28212 19790
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 28172 18896 28224 18902
rect 28172 18838 28224 18844
rect 28184 18358 28212 18838
rect 28276 18698 28304 19314
rect 28264 18692 28316 18698
rect 28264 18634 28316 18640
rect 28172 18352 28224 18358
rect 28172 18294 28224 18300
rect 28172 18216 28224 18222
rect 28368 18170 28396 20742
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28224 18164 28396 18170
rect 28172 18158 28396 18164
rect 28184 18142 28396 18158
rect 27894 16079 27896 16088
rect 27948 16079 27950 16088
rect 28080 16108 28132 16114
rect 27896 16050 27948 16056
rect 28080 16050 28132 16056
rect 28080 15360 28132 15366
rect 28080 15302 28132 15308
rect 27896 14408 27948 14414
rect 27896 14350 27948 14356
rect 27908 14074 27936 14350
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 27804 14000 27856 14006
rect 27804 13942 27856 13948
rect 28092 12442 28120 15302
rect 27620 12436 27672 12442
rect 27620 12378 27672 12384
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 27528 12368 27580 12374
rect 27528 12310 27580 12316
rect 27540 12220 27568 12310
rect 28184 12238 28212 18142
rect 28460 16998 28488 20334
rect 28540 19780 28592 19786
rect 28540 19722 28592 19728
rect 28552 19174 28580 19722
rect 28540 19168 28592 19174
rect 28540 19110 28592 19116
rect 28448 16992 28500 16998
rect 28448 16934 28500 16940
rect 28264 16516 28316 16522
rect 28264 16458 28316 16464
rect 28276 16114 28304 16458
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 27620 12232 27672 12238
rect 27540 12192 27620 12220
rect 27540 11898 27568 12192
rect 27988 12232 28040 12238
rect 27620 12174 27672 12180
rect 27908 12192 27988 12220
rect 27710 11928 27766 11937
rect 27528 11892 27580 11898
rect 27710 11863 27766 11872
rect 27528 11834 27580 11840
rect 27724 11762 27752 11863
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27528 11552 27580 11558
rect 27448 11512 27528 11540
rect 27344 9376 27396 9382
rect 27344 9318 27396 9324
rect 27342 9072 27398 9081
rect 27342 9007 27398 9016
rect 27356 8974 27384 9007
rect 27344 8968 27396 8974
rect 27344 8910 27396 8916
rect 27252 8084 27304 8090
rect 27252 8026 27304 8032
rect 27264 7886 27292 8026
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 27448 7546 27476 11512
rect 27528 11494 27580 11500
rect 27632 11354 27660 11698
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27804 11212 27856 11218
rect 27804 11154 27856 11160
rect 27816 10810 27844 11154
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 27620 10600 27672 10606
rect 27620 10542 27672 10548
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 27540 10198 27568 10474
rect 27528 10192 27580 10198
rect 27528 10134 27580 10140
rect 27540 10062 27568 10134
rect 27632 10130 27660 10542
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27724 10062 27752 10746
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27804 9920 27856 9926
rect 27908 9908 27936 12192
rect 27988 12174 28040 12180
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28080 11620 28132 11626
rect 28080 11562 28132 11568
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 28000 10198 28028 11086
rect 28092 10674 28120 11562
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 28080 10464 28132 10470
rect 28080 10406 28132 10412
rect 27988 10192 28040 10198
rect 27988 10134 28040 10140
rect 28092 10062 28120 10406
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 27856 9880 27936 9908
rect 27804 9862 27856 9868
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27436 7540 27488 7546
rect 27436 7482 27488 7488
rect 27540 7206 27568 9454
rect 27620 9444 27672 9450
rect 27620 9386 27672 9392
rect 27632 8906 27660 9386
rect 27816 9042 27844 9862
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27620 8900 27672 8906
rect 27620 8842 27672 8848
rect 27802 7984 27858 7993
rect 27802 7919 27804 7928
rect 27856 7919 27858 7928
rect 27804 7890 27856 7896
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27540 7002 27568 7142
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27816 6769 27844 7890
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 27908 7546 27936 7822
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 27908 7410 27936 7482
rect 28092 7478 28120 9998
rect 28184 9518 28212 11086
rect 28276 9625 28304 16050
rect 28356 14340 28408 14346
rect 28356 14282 28408 14288
rect 28368 12442 28396 14282
rect 28356 12436 28408 12442
rect 28644 12434 28672 25774
rect 28828 24857 28856 26522
rect 28920 24886 28948 28630
rect 29000 27940 29052 27946
rect 29000 27882 29052 27888
rect 29012 27674 29040 27882
rect 29092 27872 29144 27878
rect 29092 27814 29144 27820
rect 29000 27668 29052 27674
rect 29000 27610 29052 27616
rect 29104 27402 29132 27814
rect 29184 27600 29236 27606
rect 29184 27542 29236 27548
rect 29092 27396 29144 27402
rect 29092 27338 29144 27344
rect 29196 25906 29224 27542
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 28908 24880 28960 24886
rect 28814 24848 28870 24857
rect 28908 24822 28960 24828
rect 28814 24783 28870 24792
rect 28816 24744 28868 24750
rect 28722 24712 28778 24721
rect 28816 24686 28868 24692
rect 28722 24647 28778 24656
rect 28736 24614 28764 24647
rect 28724 24608 28776 24614
rect 28724 24550 28776 24556
rect 28722 24440 28778 24449
rect 28828 24410 28856 24686
rect 28722 24375 28778 24384
rect 28816 24404 28868 24410
rect 28736 22642 28764 24375
rect 28816 24346 28868 24352
rect 28816 23724 28868 23730
rect 28816 23666 28868 23672
rect 28828 23497 28856 23666
rect 28920 23526 28948 24822
rect 28908 23520 28960 23526
rect 28814 23488 28870 23497
rect 28908 23462 28960 23468
rect 28814 23423 28870 23432
rect 28724 22636 28776 22642
rect 28724 22578 28776 22584
rect 28816 21548 28868 21554
rect 28816 21490 28868 21496
rect 28828 20398 28856 21490
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28828 20058 28856 20334
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28724 18964 28776 18970
rect 28724 18906 28776 18912
rect 28356 12378 28408 12384
rect 28460 12406 28672 12434
rect 28356 11144 28408 11150
rect 28356 11086 28408 11092
rect 28368 10810 28396 11086
rect 28460 11014 28488 12406
rect 28540 11280 28592 11286
rect 28540 11222 28592 11228
rect 28552 11082 28580 11222
rect 28736 11200 28764 18906
rect 28920 18902 28948 23462
rect 29012 22273 29040 25230
rect 29288 24936 29316 31878
rect 29380 31754 29408 32932
rect 29932 32910 29960 33526
rect 30012 33040 30064 33046
rect 30012 32982 30064 32988
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 30024 32502 30052 32982
rect 29920 32496 29972 32502
rect 29920 32438 29972 32444
rect 30012 32496 30064 32502
rect 30012 32438 30064 32444
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 29828 32428 29880 32434
rect 29828 32370 29880 32376
rect 29460 32360 29512 32366
rect 29512 32320 29592 32348
rect 29460 32302 29512 32308
rect 29460 32224 29512 32230
rect 29460 32166 29512 32172
rect 29368 31748 29420 31754
rect 29368 31690 29420 31696
rect 29380 30734 29408 31690
rect 29368 30728 29420 30734
rect 29368 30670 29420 30676
rect 29366 30288 29422 30297
rect 29366 30223 29368 30232
rect 29420 30223 29422 30232
rect 29368 30194 29420 30200
rect 29368 27872 29420 27878
rect 29368 27814 29420 27820
rect 29380 25838 29408 27814
rect 29472 26382 29500 32166
rect 29564 31793 29592 32320
rect 29656 32230 29684 32370
rect 29736 32292 29788 32298
rect 29736 32234 29788 32240
rect 29644 32224 29696 32230
rect 29644 32166 29696 32172
rect 29550 31784 29606 31793
rect 29550 31719 29606 31728
rect 29748 31736 29776 32234
rect 29840 32026 29868 32370
rect 29932 32230 29960 32438
rect 29920 32224 29972 32230
rect 29920 32166 29972 32172
rect 29918 32056 29974 32065
rect 29828 32020 29880 32026
rect 29918 31991 29974 32000
rect 29828 31962 29880 31968
rect 29828 31748 29880 31754
rect 29748 31708 29828 31736
rect 29552 30592 29604 30598
rect 29552 30534 29604 30540
rect 29564 30258 29592 30534
rect 29552 30252 29604 30258
rect 29552 30194 29604 30200
rect 29644 30048 29696 30054
rect 29644 29990 29696 29996
rect 29552 29164 29604 29170
rect 29552 29106 29604 29112
rect 29564 28762 29592 29106
rect 29552 28756 29604 28762
rect 29552 28698 29604 28704
rect 29552 28484 29604 28490
rect 29552 28426 29604 28432
rect 29460 26376 29512 26382
rect 29460 26318 29512 26324
rect 29368 25832 29420 25838
rect 29420 25780 29500 25786
rect 29368 25774 29500 25780
rect 29380 25758 29500 25774
rect 29368 25696 29420 25702
rect 29366 25664 29368 25673
rect 29420 25664 29422 25673
rect 29366 25599 29422 25608
rect 29104 24908 29316 24936
rect 29368 24948 29420 24954
rect 28998 22264 29054 22273
rect 28998 22199 29054 22208
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 29012 21146 29040 21966
rect 29000 21140 29052 21146
rect 29000 21082 29052 21088
rect 29012 19378 29040 21082
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 28908 18896 28960 18902
rect 28908 18838 28960 18844
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 28920 17882 28948 18566
rect 29012 18290 29040 19314
rect 29104 19310 29132 24908
rect 29368 24890 29420 24896
rect 29276 24744 29328 24750
rect 29276 24686 29328 24692
rect 29288 24206 29316 24686
rect 29276 24200 29328 24206
rect 29276 24142 29328 24148
rect 29288 24070 29316 24142
rect 29276 24064 29328 24070
rect 29276 24006 29328 24012
rect 29184 23724 29236 23730
rect 29184 23666 29236 23672
rect 29196 23322 29224 23666
rect 29276 23520 29328 23526
rect 29276 23462 29328 23468
rect 29184 23316 29236 23322
rect 29184 23258 29236 23264
rect 29184 21548 29236 21554
rect 29184 21490 29236 21496
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 29196 18970 29224 21490
rect 29288 19854 29316 23462
rect 29380 21078 29408 24890
rect 29368 21072 29420 21078
rect 29368 21014 29420 21020
rect 29368 20528 29420 20534
rect 29368 20470 29420 20476
rect 29380 19922 29408 20470
rect 29368 19916 29420 19922
rect 29368 19858 29420 19864
rect 29276 19848 29328 19854
rect 29276 19790 29328 19796
rect 29184 18964 29236 18970
rect 29184 18906 29236 18912
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28828 17134 28856 17614
rect 28816 17128 28868 17134
rect 28816 17070 28868 17076
rect 28828 16794 28856 17070
rect 28816 16788 28868 16794
rect 28816 16730 28868 16736
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28828 13938 28856 14214
rect 28920 13938 28948 17818
rect 29276 17604 29328 17610
rect 29276 17546 29328 17552
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 29092 14340 29144 14346
rect 29092 14282 29144 14288
rect 29104 14006 29132 14282
rect 29092 14000 29144 14006
rect 29092 13942 29144 13948
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 29000 13932 29052 13938
rect 29000 13874 29052 13880
rect 29012 13530 29040 13874
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 28816 13252 28868 13258
rect 28816 13194 28868 13200
rect 28828 12646 28856 13194
rect 28816 12640 28868 12646
rect 28816 12582 28868 12588
rect 28644 11172 28764 11200
rect 28540 11076 28592 11082
rect 28540 11018 28592 11024
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28460 10470 28488 10950
rect 28552 10606 28580 11018
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 28448 10464 28500 10470
rect 28448 10406 28500 10412
rect 28460 10146 28488 10406
rect 28460 10118 28580 10146
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28368 9654 28396 9998
rect 28460 9722 28488 9998
rect 28552 9722 28580 10118
rect 28644 9926 28672 11172
rect 28828 11150 28856 12582
rect 29196 12374 29224 16526
rect 29288 16114 29316 17546
rect 29276 16108 29328 16114
rect 29276 16050 29328 16056
rect 29288 12481 29316 16050
rect 29380 15978 29408 19858
rect 29472 16114 29500 25758
rect 29564 24954 29592 28426
rect 29656 28082 29684 29990
rect 29644 28076 29696 28082
rect 29644 28018 29696 28024
rect 29748 27946 29776 31708
rect 29828 31690 29880 31696
rect 29828 31340 29880 31346
rect 29932 31328 29960 31991
rect 30116 31822 30144 35866
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 31668 34536 31720 34542
rect 31668 34478 31720 34484
rect 30196 33992 30248 33998
rect 30196 33934 30248 33940
rect 30208 32609 30236 33934
rect 31576 33856 31628 33862
rect 31576 33798 31628 33804
rect 31392 33448 31444 33454
rect 31392 33390 31444 33396
rect 31404 33114 31432 33390
rect 31392 33108 31444 33114
rect 31392 33050 31444 33056
rect 31588 32910 31616 33798
rect 31680 33522 31708 34478
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 32496 33992 32548 33998
rect 32496 33934 32548 33940
rect 32312 33652 32364 33658
rect 32312 33594 32364 33600
rect 31668 33516 31720 33522
rect 31668 33458 31720 33464
rect 31680 32978 31708 33458
rect 32220 33312 32272 33318
rect 32324 33266 32352 33594
rect 32404 33448 32456 33454
rect 32404 33390 32456 33396
rect 32272 33260 32352 33266
rect 32220 33254 32352 33260
rect 32232 33238 32352 33254
rect 31668 32972 31720 32978
rect 31668 32914 31720 32920
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 31576 32904 31628 32910
rect 31404 32864 31576 32892
rect 30380 32768 30432 32774
rect 31116 32768 31168 32774
rect 30380 32710 30432 32716
rect 31114 32736 31116 32745
rect 31168 32736 31170 32745
rect 31298 32736 31354 32745
rect 30194 32600 30250 32609
rect 30392 32570 30420 32710
rect 31170 32694 31248 32722
rect 31114 32671 31170 32680
rect 30194 32535 30250 32544
rect 30288 32564 30340 32570
rect 30208 32434 30236 32535
rect 30288 32506 30340 32512
rect 30380 32564 30432 32570
rect 30380 32506 30432 32512
rect 30748 32564 30800 32570
rect 30748 32506 30800 32512
rect 30300 32450 30328 32506
rect 30196 32428 30248 32434
rect 30300 32422 30420 32450
rect 30196 32370 30248 32376
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30104 31816 30156 31822
rect 30104 31758 30156 31764
rect 29880 31300 29960 31328
rect 29828 31282 29880 31288
rect 29840 29850 29868 31282
rect 30024 31142 30052 31758
rect 30116 31210 30144 31758
rect 30208 31521 30236 32370
rect 30392 32201 30420 32422
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30378 32192 30434 32201
rect 30378 32127 30434 32136
rect 30392 32026 30420 32127
rect 30484 32065 30512 32370
rect 30656 32360 30708 32366
rect 30654 32328 30656 32337
rect 30708 32328 30710 32337
rect 30654 32263 30710 32272
rect 30470 32056 30526 32065
rect 30380 32020 30432 32026
rect 30470 31991 30526 32000
rect 30380 31962 30432 31968
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30472 31816 30524 31822
rect 30524 31764 30604 31770
rect 30472 31758 30604 31764
rect 30194 31512 30250 31521
rect 30194 31447 30250 31456
rect 30392 31346 30420 31758
rect 30484 31742 30604 31758
rect 30472 31680 30524 31686
rect 30470 31648 30472 31657
rect 30524 31648 30526 31657
rect 30470 31583 30526 31592
rect 30484 31346 30512 31583
rect 30196 31340 30248 31346
rect 30196 31282 30248 31288
rect 30380 31340 30432 31346
rect 30380 31282 30432 31288
rect 30472 31340 30524 31346
rect 30472 31282 30524 31288
rect 30104 31204 30156 31210
rect 30104 31146 30156 31152
rect 30208 31142 30236 31282
rect 30576 31278 30604 31742
rect 30760 31634 30788 32506
rect 31024 32496 31076 32502
rect 31024 32438 31076 32444
rect 30932 32360 30984 32366
rect 31036 32337 31064 32438
rect 30932 32302 30984 32308
rect 31022 32328 31078 32337
rect 30838 32056 30894 32065
rect 30838 31991 30894 32000
rect 30852 31958 30880 31991
rect 30840 31952 30892 31958
rect 30840 31894 30892 31900
rect 30944 31822 30972 32302
rect 31022 32263 31078 32272
rect 31116 31884 31168 31890
rect 31116 31826 31168 31832
rect 30932 31816 30984 31822
rect 30932 31758 30984 31764
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 30760 31606 30880 31634
rect 30748 31476 30800 31482
rect 30748 31418 30800 31424
rect 30760 31278 30788 31418
rect 30564 31272 30616 31278
rect 30286 31240 30342 31249
rect 30564 31214 30616 31220
rect 30748 31272 30800 31278
rect 30748 31214 30800 31220
rect 30286 31175 30288 31184
rect 30340 31175 30342 31184
rect 30288 31146 30340 31152
rect 30012 31136 30064 31142
rect 30012 31078 30064 31084
rect 30196 31136 30248 31142
rect 30196 31078 30248 31084
rect 30024 30734 30052 31078
rect 30208 30734 30236 31078
rect 30300 30802 30328 31146
rect 30472 30864 30524 30870
rect 30472 30806 30524 30812
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 30196 30728 30248 30734
rect 30196 30670 30248 30676
rect 30012 30320 30064 30326
rect 30012 30262 30064 30268
rect 29828 29844 29880 29850
rect 29828 29786 29880 29792
rect 30024 29073 30052 30262
rect 30208 30258 30236 30670
rect 30196 30252 30248 30258
rect 30196 30194 30248 30200
rect 30484 30122 30512 30806
rect 30760 30666 30788 31214
rect 30748 30660 30800 30666
rect 30748 30602 30800 30608
rect 30852 30569 30880 31606
rect 30838 30560 30894 30569
rect 30838 30495 30894 30504
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 30472 30116 30524 30122
rect 30472 30058 30524 30064
rect 30564 30048 30616 30054
rect 30668 30025 30696 30194
rect 30564 29990 30616 29996
rect 30654 30016 30710 30025
rect 30472 29640 30524 29646
rect 30472 29582 30524 29588
rect 30288 29572 30340 29578
rect 30288 29514 30340 29520
rect 30010 29064 30066 29073
rect 30010 28999 30012 29008
rect 30064 28999 30066 29008
rect 30012 28970 30064 28976
rect 29920 28756 29972 28762
rect 29920 28698 29972 28704
rect 29932 28558 29960 28698
rect 30104 28620 30156 28626
rect 30104 28562 30156 28568
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 29828 28484 29880 28490
rect 29828 28426 29880 28432
rect 29736 27940 29788 27946
rect 29736 27882 29788 27888
rect 29840 27538 29868 28426
rect 30010 28384 30066 28393
rect 30010 28319 30066 28328
rect 30024 28150 30052 28319
rect 30012 28144 30064 28150
rect 29918 28112 29974 28121
rect 30012 28086 30064 28092
rect 29918 28047 29920 28056
rect 29972 28047 29974 28056
rect 29920 28018 29972 28024
rect 30012 28008 30064 28014
rect 30116 27996 30144 28562
rect 30196 28552 30248 28558
rect 30196 28494 30248 28500
rect 30208 28082 30236 28494
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 30064 27968 30144 27996
rect 30012 27950 30064 27956
rect 29828 27532 29880 27538
rect 29828 27474 29880 27480
rect 29644 26376 29696 26382
rect 29920 26376 29972 26382
rect 29644 26318 29696 26324
rect 29748 26336 29920 26364
rect 29656 26042 29684 26318
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 29748 25770 29776 26336
rect 29920 26318 29972 26324
rect 30024 25974 30052 27950
rect 30208 27674 30236 28018
rect 30196 27668 30248 27674
rect 30196 27610 30248 27616
rect 30102 27568 30158 27577
rect 30102 27503 30104 27512
rect 30156 27503 30158 27512
rect 30104 27474 30156 27480
rect 30104 27328 30156 27334
rect 30104 27270 30156 27276
rect 30012 25968 30064 25974
rect 30012 25910 30064 25916
rect 29736 25764 29788 25770
rect 29736 25706 29788 25712
rect 29552 24948 29604 24954
rect 29552 24890 29604 24896
rect 29644 24880 29696 24886
rect 29644 24822 29696 24828
rect 29656 24750 29684 24822
rect 29644 24744 29696 24750
rect 29644 24686 29696 24692
rect 29656 23662 29684 24686
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29748 22094 29776 25706
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 29828 24744 29880 24750
rect 29828 24686 29880 24692
rect 29840 24614 29868 24686
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 29656 22066 29776 22094
rect 29552 21548 29604 21554
rect 29552 21490 29604 21496
rect 29564 21146 29592 21490
rect 29552 21140 29604 21146
rect 29552 21082 29604 21088
rect 29552 20256 29604 20262
rect 29552 20198 29604 20204
rect 29564 20058 29592 20198
rect 29552 20052 29604 20058
rect 29552 19994 29604 20000
rect 29656 19446 29684 22066
rect 29932 21690 29960 25638
rect 30024 25158 30052 25910
rect 30012 25152 30064 25158
rect 30012 25094 30064 25100
rect 30010 24984 30066 24993
rect 30010 24919 30066 24928
rect 30024 24274 30052 24919
rect 30012 24268 30064 24274
rect 30012 24210 30064 24216
rect 30012 21888 30064 21894
rect 30012 21830 30064 21836
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 29644 19440 29696 19446
rect 29644 19382 29696 19388
rect 29656 18766 29684 19382
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29644 18760 29696 18766
rect 29644 18702 29696 18708
rect 29564 17746 29592 18702
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29656 17678 29684 18226
rect 29644 17672 29696 17678
rect 29644 17614 29696 17620
rect 29644 17536 29696 17542
rect 29644 17478 29696 17484
rect 29656 16998 29684 17478
rect 29748 16998 29776 19858
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29840 18766 29868 19246
rect 30024 19174 30052 21830
rect 30116 21554 30144 27270
rect 30196 25696 30248 25702
rect 30194 25664 30196 25673
rect 30248 25664 30250 25673
rect 30194 25599 30250 25608
rect 30300 25514 30328 29514
rect 30378 29472 30434 29481
rect 30378 29407 30434 29416
rect 30392 29238 30420 29407
rect 30380 29232 30432 29238
rect 30380 29174 30432 29180
rect 30484 29102 30512 29582
rect 30472 29096 30524 29102
rect 30472 29038 30524 29044
rect 30576 28082 30604 29990
rect 30654 29951 30710 29960
rect 30852 29696 30880 30495
rect 30760 29668 30880 29696
rect 30760 29617 30788 29668
rect 30746 29608 30802 29617
rect 30746 29543 30748 29552
rect 30800 29543 30802 29552
rect 30840 29572 30892 29578
rect 30748 29514 30800 29520
rect 30840 29514 30892 29520
rect 30748 29232 30800 29238
rect 30748 29174 30800 29180
rect 30656 29164 30708 29170
rect 30656 29106 30708 29112
rect 30668 28966 30696 29106
rect 30656 28960 30708 28966
rect 30656 28902 30708 28908
rect 30564 28076 30616 28082
rect 30564 28018 30616 28024
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30392 27577 30420 27950
rect 30472 27940 30524 27946
rect 30472 27882 30524 27888
rect 30378 27568 30434 27577
rect 30378 27503 30434 27512
rect 30380 26512 30432 26518
rect 30380 26454 30432 26460
rect 30208 25486 30328 25514
rect 30104 21548 30156 21554
rect 30104 21490 30156 21496
rect 30208 19394 30236 25486
rect 30288 24676 30340 24682
rect 30288 24618 30340 24624
rect 30300 24342 30328 24618
rect 30288 24336 30340 24342
rect 30288 24278 30340 24284
rect 30288 22432 30340 22438
rect 30288 22374 30340 22380
rect 30300 22098 30328 22374
rect 30288 22092 30340 22098
rect 30288 22034 30340 22040
rect 30392 21962 30420 26454
rect 30380 21956 30432 21962
rect 30380 21898 30432 21904
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 30300 20466 30328 20742
rect 30288 20460 30340 20466
rect 30288 20402 30340 20408
rect 30116 19366 30236 19394
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 29828 18760 29880 18766
rect 30116 18748 30144 19366
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 30208 18970 30236 19246
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 30300 18850 30328 20402
rect 30484 20262 30512 27882
rect 30576 26042 30604 28018
rect 30656 27532 30708 27538
rect 30656 27474 30708 27480
rect 30564 26036 30616 26042
rect 30564 25978 30616 25984
rect 30668 25786 30696 27474
rect 30760 27334 30788 29174
rect 30852 28966 30880 29514
rect 30944 29510 30972 31758
rect 31036 31482 31064 31758
rect 31024 31476 31076 31482
rect 31024 31418 31076 31424
rect 31128 30297 31156 31826
rect 31114 30288 31170 30297
rect 31114 30223 31116 30232
rect 31168 30223 31170 30232
rect 31116 30194 31168 30200
rect 31022 30016 31078 30025
rect 31022 29951 31078 29960
rect 30932 29504 30984 29510
rect 30932 29446 30984 29452
rect 30944 29238 30972 29446
rect 30932 29232 30984 29238
rect 30932 29174 30984 29180
rect 30840 28960 30892 28966
rect 30840 28902 30892 28908
rect 30852 28422 30880 28902
rect 30840 28416 30892 28422
rect 30840 28358 30892 28364
rect 30748 27328 30800 27334
rect 30748 27270 30800 27276
rect 30852 27146 30880 28358
rect 31036 27985 31064 29951
rect 31116 29504 31168 29510
rect 31116 29446 31168 29452
rect 31022 27976 31078 27985
rect 31022 27911 31078 27920
rect 31036 27674 31064 27911
rect 31024 27668 31076 27674
rect 31024 27610 31076 27616
rect 31128 27606 31156 29446
rect 31220 27606 31248 32694
rect 31298 32671 31354 32680
rect 31312 32570 31340 32671
rect 31300 32564 31352 32570
rect 31300 32506 31352 32512
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 31312 32026 31340 32370
rect 31300 32020 31352 32026
rect 31300 31962 31352 31968
rect 31312 31822 31340 31962
rect 31404 31890 31432 32864
rect 31576 32846 31628 32852
rect 31944 32904 31996 32910
rect 31944 32846 31996 32852
rect 31850 32600 31906 32609
rect 31850 32535 31906 32544
rect 31864 32502 31892 32535
rect 31852 32496 31904 32502
rect 31574 32464 31630 32473
rect 31852 32438 31904 32444
rect 31574 32399 31576 32408
rect 31628 32399 31630 32408
rect 31576 32370 31628 32376
rect 31484 32360 31536 32366
rect 31484 32302 31536 32308
rect 31392 31884 31444 31890
rect 31392 31826 31444 31832
rect 31300 31816 31352 31822
rect 31300 31758 31352 31764
rect 31496 31754 31524 32302
rect 31576 32292 31628 32298
rect 31576 32234 31628 32240
rect 31588 32008 31616 32234
rect 31956 32201 31984 32846
rect 32140 32298 32168 32914
rect 32220 32904 32272 32910
rect 32220 32846 32272 32852
rect 32232 32745 32260 32846
rect 32218 32736 32274 32745
rect 32218 32671 32274 32680
rect 32232 32570 32260 32671
rect 32220 32564 32272 32570
rect 32220 32506 32272 32512
rect 32324 32366 32352 33238
rect 32416 33114 32444 33390
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 32404 32904 32456 32910
rect 32404 32846 32456 32852
rect 32312 32360 32364 32366
rect 32416 32337 32444 32846
rect 32312 32302 32364 32308
rect 32402 32328 32458 32337
rect 32128 32292 32180 32298
rect 32402 32263 32458 32272
rect 32128 32234 32180 32240
rect 31942 32192 31998 32201
rect 31942 32127 31998 32136
rect 32218 32056 32274 32065
rect 31588 31980 31708 32008
rect 32218 31991 32274 32000
rect 32312 32020 32364 32026
rect 31576 31884 31628 31890
rect 31576 31826 31628 31832
rect 31484 31748 31536 31754
rect 31484 31690 31536 31696
rect 31392 31680 31444 31686
rect 31312 31628 31392 31634
rect 31312 31622 31444 31628
rect 31312 31606 31432 31622
rect 31312 31278 31340 31606
rect 31300 31272 31352 31278
rect 31300 31214 31352 31220
rect 31496 30938 31524 31690
rect 31484 30932 31536 30938
rect 31484 30874 31536 30880
rect 31300 30592 31352 30598
rect 31300 30534 31352 30540
rect 31116 27600 31168 27606
rect 31022 27568 31078 27577
rect 30932 27532 30984 27538
rect 31116 27542 31168 27548
rect 31208 27600 31260 27606
rect 31208 27542 31260 27548
rect 31022 27503 31078 27512
rect 30932 27474 30984 27480
rect 30944 27334 30972 27474
rect 31036 27470 31064 27503
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 30932 27328 30984 27334
rect 30932 27270 30984 27276
rect 30576 25758 30696 25786
rect 30760 27118 30880 27146
rect 30576 24052 30604 25758
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30668 24206 30696 24686
rect 30656 24200 30708 24206
rect 30656 24142 30708 24148
rect 30576 24024 30696 24052
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 30576 22982 30604 23734
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30668 22098 30696 24024
rect 30760 23202 30788 27118
rect 30944 26518 30972 27270
rect 31208 26920 31260 26926
rect 31208 26862 31260 26868
rect 30932 26512 30984 26518
rect 30932 26454 30984 26460
rect 31024 25900 31076 25906
rect 31024 25842 31076 25848
rect 30932 24336 30984 24342
rect 30930 24304 30932 24313
rect 30984 24304 30986 24313
rect 30930 24239 30986 24248
rect 31036 24206 31064 25842
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 30932 24132 30984 24138
rect 30932 24074 30984 24080
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30852 23338 30880 24006
rect 30944 23497 30972 24074
rect 31036 23730 31064 24142
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 31116 23724 31168 23730
rect 31116 23666 31168 23672
rect 31128 23526 31156 23666
rect 31116 23520 31168 23526
rect 30930 23488 30986 23497
rect 31116 23462 31168 23468
rect 30930 23423 30986 23432
rect 30852 23310 30972 23338
rect 30760 23174 30880 23202
rect 30852 22574 30880 23174
rect 30840 22568 30892 22574
rect 30840 22510 30892 22516
rect 30748 22500 30800 22506
rect 30748 22442 30800 22448
rect 30656 22092 30708 22098
rect 30656 22034 30708 22040
rect 30760 21962 30788 22442
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30760 21350 30788 21898
rect 30748 21344 30800 21350
rect 30748 21286 30800 21292
rect 30760 20466 30788 21286
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30748 20460 30800 20466
rect 30748 20402 30800 20408
rect 30472 20256 30524 20262
rect 30472 20198 30524 20204
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30392 19417 30420 19450
rect 30378 19408 30434 19417
rect 30378 19343 30434 19352
rect 30472 19236 30524 19242
rect 30472 19178 30524 19184
rect 29828 18702 29880 18708
rect 29932 18720 30144 18748
rect 30208 18822 30328 18850
rect 29840 18086 29868 18702
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29828 17604 29880 17610
rect 29828 17546 29880 17552
rect 29644 16992 29696 16998
rect 29644 16934 29696 16940
rect 29736 16992 29788 16998
rect 29736 16934 29788 16940
rect 29748 16250 29776 16934
rect 29736 16244 29788 16250
rect 29656 16204 29736 16232
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29368 15972 29420 15978
rect 29368 15914 29420 15920
rect 29656 14414 29684 16204
rect 29736 16186 29788 16192
rect 29840 15366 29868 17546
rect 29828 15360 29880 15366
rect 29828 15302 29880 15308
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29828 14000 29880 14006
rect 29828 13942 29880 13948
rect 29460 13796 29512 13802
rect 29460 13738 29512 13744
rect 29472 12986 29500 13738
rect 29644 13388 29696 13394
rect 29644 13330 29696 13336
rect 29656 13258 29684 13330
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29460 12980 29512 12986
rect 29460 12922 29512 12928
rect 29274 12472 29330 12481
rect 29274 12407 29330 12416
rect 29184 12368 29236 12374
rect 29184 12310 29236 12316
rect 29184 12232 29236 12238
rect 29184 12174 29236 12180
rect 29092 12164 29144 12170
rect 29092 12106 29144 12112
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29012 11665 29040 11698
rect 28998 11656 29054 11665
rect 28998 11591 29054 11600
rect 29000 11552 29052 11558
rect 29000 11494 29052 11500
rect 29012 11150 29040 11494
rect 29104 11150 29132 12106
rect 28816 11144 28868 11150
rect 28816 11086 28868 11092
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 28724 11008 28776 11014
rect 28724 10950 28776 10956
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 28736 10674 28764 10950
rect 28816 10804 28868 10810
rect 28816 10746 28868 10752
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28828 10606 28856 10746
rect 28908 10736 28960 10742
rect 28908 10678 28960 10684
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28632 9920 28684 9926
rect 28632 9862 28684 9868
rect 28448 9716 28500 9722
rect 28448 9658 28500 9664
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28356 9648 28408 9654
rect 28262 9616 28318 9625
rect 28356 9590 28408 9596
rect 28262 9551 28318 9560
rect 28172 9512 28224 9518
rect 28172 9454 28224 9460
rect 28080 7472 28132 7478
rect 28080 7414 28132 7420
rect 27896 7404 27948 7410
rect 27896 7346 27948 7352
rect 28170 7168 28226 7177
rect 28170 7103 28226 7112
rect 27802 6760 27858 6769
rect 27620 6724 27672 6730
rect 27802 6695 27858 6704
rect 27620 6666 27672 6672
rect 27252 6656 27304 6662
rect 27252 6598 27304 6604
rect 27344 6656 27396 6662
rect 27632 6610 27660 6666
rect 27344 6598 27396 6604
rect 27264 6390 27292 6598
rect 27252 6384 27304 6390
rect 27252 6326 27304 6332
rect 27356 6322 27384 6598
rect 27540 6582 27660 6610
rect 27540 6361 27568 6582
rect 27526 6352 27582 6361
rect 27344 6316 27396 6322
rect 27526 6287 27582 6296
rect 27344 6258 27396 6264
rect 27172 6174 27384 6202
rect 27252 5840 27304 5846
rect 27252 5782 27304 5788
rect 26976 5704 27028 5710
rect 27264 5692 27292 5782
rect 27028 5664 27292 5692
rect 26976 5646 27028 5652
rect 27356 5574 27384 6174
rect 27344 5568 27396 5574
rect 27344 5510 27396 5516
rect 26884 5228 26936 5234
rect 26884 5170 26936 5176
rect 27356 5030 27384 5510
rect 27436 5228 27488 5234
rect 27436 5170 27488 5176
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 26896 3534 26924 3878
rect 26988 3670 27016 4966
rect 27448 4010 27476 5170
rect 27436 4004 27488 4010
rect 27436 3946 27488 3952
rect 27068 3936 27120 3942
rect 27068 3878 27120 3884
rect 26976 3664 27028 3670
rect 26976 3606 27028 3612
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 25412 3460 25464 3466
rect 25412 3402 25464 3408
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 26160 3058 26188 3470
rect 27080 3398 27108 3878
rect 27448 3738 27476 3946
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 27540 3534 27568 6287
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 28000 5710 28028 5782
rect 27988 5704 28040 5710
rect 27988 5646 28040 5652
rect 28184 5574 28212 7103
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 28276 3602 28304 9551
rect 28368 9110 28396 9590
rect 28356 9104 28408 9110
rect 28356 9046 28408 9052
rect 28736 8945 28764 9998
rect 28828 9994 28856 10542
rect 28920 10044 28948 10678
rect 29012 10674 29040 10950
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 29090 10568 29146 10577
rect 29090 10503 29092 10512
rect 29144 10503 29146 10512
rect 29092 10474 29144 10480
rect 29196 10470 29224 12174
rect 29184 10464 29236 10470
rect 29184 10406 29236 10412
rect 29288 10130 29316 12407
rect 29472 12170 29500 12922
rect 29656 12306 29684 13194
rect 29840 12646 29868 13942
rect 29932 13870 29960 18720
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30116 17678 30144 18566
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 30012 17604 30064 17610
rect 30012 17546 30064 17552
rect 30024 17270 30052 17546
rect 30012 17264 30064 17270
rect 30012 17206 30064 17212
rect 30208 17202 30236 18822
rect 30484 18698 30512 19178
rect 30564 19168 30616 19174
rect 30564 19110 30616 19116
rect 30472 18692 30524 18698
rect 30472 18634 30524 18640
rect 30576 17678 30604 19110
rect 30668 18970 30696 20402
rect 30656 18964 30708 18970
rect 30656 18906 30708 18912
rect 30760 18766 30788 20402
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 30760 18426 30788 18702
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30472 17604 30524 17610
rect 30472 17546 30524 17552
rect 30288 17536 30340 17542
rect 30288 17478 30340 17484
rect 30300 17270 30328 17478
rect 30288 17264 30340 17270
rect 30484 17218 30512 17546
rect 30654 17368 30710 17377
rect 30654 17303 30656 17312
rect 30708 17303 30710 17312
rect 30656 17274 30708 17280
rect 30288 17206 30340 17212
rect 30196 17196 30248 17202
rect 30196 17138 30248 17144
rect 30392 17190 30512 17218
rect 30564 17196 30616 17202
rect 30392 17082 30420 17190
rect 30564 17138 30616 17144
rect 30300 17054 30420 17082
rect 30104 16040 30156 16046
rect 30104 15982 30156 15988
rect 30012 14340 30064 14346
rect 30012 14282 30064 14288
rect 29920 13864 29972 13870
rect 29920 13806 29972 13812
rect 29828 12640 29880 12646
rect 29828 12582 29880 12588
rect 29736 12368 29788 12374
rect 29736 12310 29788 12316
rect 29644 12300 29696 12306
rect 29644 12242 29696 12248
rect 29460 12164 29512 12170
rect 29460 12106 29512 12112
rect 29552 12164 29604 12170
rect 29552 12106 29604 12112
rect 29564 12050 29592 12106
rect 29472 12022 29592 12050
rect 29368 11824 29420 11830
rect 29368 11766 29420 11772
rect 29184 10124 29236 10130
rect 29184 10066 29236 10072
rect 29276 10124 29328 10130
rect 29276 10066 29328 10072
rect 29092 10056 29144 10062
rect 28920 10016 29092 10044
rect 28816 9988 28868 9994
rect 28816 9930 28868 9936
rect 28920 9926 28948 10016
rect 29092 9998 29144 10004
rect 29196 10010 29224 10066
rect 29380 10010 29408 11766
rect 29472 11626 29500 12022
rect 29460 11620 29512 11626
rect 29460 11562 29512 11568
rect 29552 11620 29604 11626
rect 29552 11562 29604 11568
rect 29196 9982 29408 10010
rect 28908 9920 28960 9926
rect 29196 9897 29224 9982
rect 28908 9862 28960 9868
rect 29182 9888 29238 9897
rect 28722 8936 28778 8945
rect 28722 8871 28778 8880
rect 28538 7984 28594 7993
rect 28538 7919 28540 7928
rect 28592 7919 28594 7928
rect 28540 7890 28592 7896
rect 28552 7449 28580 7890
rect 28736 7886 28764 8871
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 28538 7440 28594 7449
rect 28538 7375 28594 7384
rect 28816 6928 28868 6934
rect 28816 6870 28868 6876
rect 28828 6458 28856 6870
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 28632 6316 28684 6322
rect 28632 6258 28684 6264
rect 28356 6112 28408 6118
rect 28356 6054 28408 6060
rect 28368 5642 28396 6054
rect 28356 5636 28408 5642
rect 28356 5578 28408 5584
rect 28644 4146 28672 6258
rect 28920 6254 28948 9862
rect 29182 9823 29238 9832
rect 28998 9752 29054 9761
rect 28998 9687 29054 9696
rect 28908 6248 28960 6254
rect 28908 6190 28960 6196
rect 28920 5778 28948 6190
rect 28908 5772 28960 5778
rect 28908 5714 28960 5720
rect 28632 4140 28684 4146
rect 28632 4082 28684 4088
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 29012 3534 29040 9687
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 29092 9104 29144 9110
rect 29092 9046 29144 9052
rect 29104 8974 29132 9046
rect 29380 8974 29408 9114
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 29472 8838 29500 11562
rect 29564 11150 29592 11562
rect 29748 11506 29776 12310
rect 29840 12170 29868 12582
rect 29828 12164 29880 12170
rect 29828 12106 29880 12112
rect 29656 11478 29776 11506
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29552 11008 29604 11014
rect 29552 10950 29604 10956
rect 29564 10606 29592 10950
rect 29656 10810 29684 11478
rect 29736 11348 29788 11354
rect 29736 11290 29788 11296
rect 29748 11014 29776 11290
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 29748 10674 29776 10950
rect 29828 10736 29880 10742
rect 29828 10678 29880 10684
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29564 9518 29592 10406
rect 29748 9926 29776 10610
rect 29840 10198 29868 10678
rect 29828 10192 29880 10198
rect 29828 10134 29880 10140
rect 29736 9920 29788 9926
rect 29736 9862 29788 9868
rect 29826 9752 29882 9761
rect 29826 9687 29882 9696
rect 29840 9586 29868 9687
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 29460 8832 29512 8838
rect 29460 8774 29512 8780
rect 29104 8566 29132 8774
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29274 8528 29330 8537
rect 29274 8463 29276 8472
rect 29328 8463 29330 8472
rect 29276 8434 29328 8440
rect 29288 7750 29316 8434
rect 29276 7744 29328 7750
rect 29276 7686 29328 7692
rect 29092 6656 29144 6662
rect 29092 6598 29144 6604
rect 29104 4146 29132 6598
rect 29564 5574 29592 9454
rect 29828 8900 29880 8906
rect 29828 8842 29880 8848
rect 29840 8498 29868 8842
rect 29920 8832 29972 8838
rect 29920 8774 29972 8780
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 29840 8090 29868 8434
rect 29828 8084 29880 8090
rect 29828 8026 29880 8032
rect 29828 7812 29880 7818
rect 29932 7800 29960 8774
rect 29880 7772 29960 7800
rect 29828 7754 29880 7760
rect 29840 6798 29868 7754
rect 30024 6882 30052 14282
rect 30116 13258 30144 15982
rect 30196 14272 30248 14278
rect 30196 14214 30248 14220
rect 30104 13252 30156 13258
rect 30104 13194 30156 13200
rect 30208 12442 30236 14214
rect 30300 13530 30328 17054
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30392 15434 30420 16458
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30484 15570 30512 16118
rect 30576 15706 30604 17138
rect 30656 17128 30708 17134
rect 30656 17070 30708 17076
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 30472 15564 30524 15570
rect 30472 15506 30524 15512
rect 30668 15502 30696 17070
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30760 15502 30788 15846
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 30748 15496 30800 15502
rect 30748 15438 30800 15444
rect 30380 15428 30432 15434
rect 30380 15370 30432 15376
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 30380 14884 30432 14890
rect 30380 14826 30432 14832
rect 30392 14346 30420 14826
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 30472 14340 30524 14346
rect 30472 14282 30524 14288
rect 30288 13524 30340 13530
rect 30288 13466 30340 13472
rect 30300 13394 30328 13466
rect 30288 13388 30340 13394
rect 30288 13330 30340 13336
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30196 12436 30248 12442
rect 30196 12378 30248 12384
rect 30102 11792 30158 11801
rect 30300 11762 30328 13194
rect 30484 12238 30512 14282
rect 30576 13530 30604 15302
rect 30668 14346 30696 15438
rect 30748 15360 30800 15366
rect 30748 15302 30800 15308
rect 30656 14340 30708 14346
rect 30656 14282 30708 14288
rect 30656 14068 30708 14074
rect 30656 14010 30708 14016
rect 30668 13841 30696 14010
rect 30654 13832 30710 13841
rect 30654 13767 30710 13776
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30656 13388 30708 13394
rect 30656 13330 30708 13336
rect 30668 13258 30696 13330
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30562 12336 30618 12345
rect 30562 12271 30618 12280
rect 30576 12238 30604 12271
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 30576 11898 30604 12174
rect 30654 12064 30710 12073
rect 30654 11999 30710 12008
rect 30564 11892 30616 11898
rect 30564 11834 30616 11840
rect 30668 11830 30696 11999
rect 30656 11824 30708 11830
rect 30656 11766 30708 11772
rect 30102 11727 30104 11736
rect 30156 11727 30158 11736
rect 30288 11756 30340 11762
rect 30104 11698 30156 11704
rect 30288 11698 30340 11704
rect 30380 11756 30432 11762
rect 30380 11698 30432 11704
rect 30300 11665 30328 11698
rect 30286 11656 30342 11665
rect 30286 11591 30342 11600
rect 30392 10792 30420 11698
rect 30300 10764 30420 10792
rect 30300 10470 30328 10764
rect 30380 10668 30432 10674
rect 30380 10610 30432 10616
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 30194 10296 30250 10305
rect 30194 10231 30250 10240
rect 30208 10130 30236 10231
rect 30196 10124 30248 10130
rect 30196 10066 30248 10072
rect 30104 8832 30156 8838
rect 30104 8774 30156 8780
rect 30116 8566 30144 8774
rect 30104 8560 30156 8566
rect 30104 8502 30156 8508
rect 30104 8288 30156 8294
rect 30104 8230 30156 8236
rect 30116 8090 30144 8230
rect 30104 8084 30156 8090
rect 30104 8026 30156 8032
rect 29932 6866 30052 6882
rect 29920 6860 30052 6866
rect 29972 6854 30052 6860
rect 29920 6802 29972 6808
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 29736 6316 29788 6322
rect 29736 6258 29788 6264
rect 29644 6180 29696 6186
rect 29644 6122 29696 6128
rect 29656 5710 29684 6122
rect 29748 5778 29776 6258
rect 29736 5772 29788 5778
rect 29736 5714 29788 5720
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29840 5234 29868 6734
rect 29932 6254 29960 6802
rect 30116 6390 30144 8026
rect 30104 6384 30156 6390
rect 30104 6326 30156 6332
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 30116 5642 30144 6326
rect 30208 5846 30236 10066
rect 30288 9920 30340 9926
rect 30288 9862 30340 9868
rect 30300 9586 30328 9862
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30392 8498 30420 10610
rect 30564 10600 30616 10606
rect 30564 10542 30616 10548
rect 30472 9988 30524 9994
rect 30472 9930 30524 9936
rect 30484 9586 30512 9930
rect 30472 9580 30524 9586
rect 30472 9522 30524 9528
rect 30484 9110 30512 9522
rect 30472 9104 30524 9110
rect 30472 9046 30524 9052
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30288 8424 30340 8430
rect 30288 8366 30340 8372
rect 30300 8022 30328 8366
rect 30288 8016 30340 8022
rect 30288 7958 30340 7964
rect 30380 8016 30432 8022
rect 30380 7958 30432 7964
rect 30300 6322 30328 7958
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30392 5914 30420 7958
rect 30484 6474 30512 9046
rect 30576 6662 30604 10542
rect 30668 8888 30696 11766
rect 30760 10826 30788 15302
rect 30852 14482 30880 22510
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 30852 14074 30880 14418
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30852 13326 30880 14010
rect 30944 13938 30972 23310
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 31036 19990 31064 22918
rect 31220 21622 31248 26862
rect 31312 24993 31340 30534
rect 31484 30252 31536 30258
rect 31484 30194 31536 30200
rect 31496 29510 31524 30194
rect 31588 30054 31616 31826
rect 31680 30870 31708 31980
rect 31852 31816 31904 31822
rect 31852 31758 31904 31764
rect 31864 31414 31892 31758
rect 31852 31408 31904 31414
rect 31852 31350 31904 31356
rect 31668 30864 31720 30870
rect 31668 30806 31720 30812
rect 31576 30048 31628 30054
rect 31576 29990 31628 29996
rect 31864 29510 31892 31350
rect 32232 31210 32260 31991
rect 32312 31962 32364 31968
rect 32324 31822 32352 31962
rect 32312 31816 32364 31822
rect 32312 31758 32364 31764
rect 32404 31748 32456 31754
rect 32404 31690 32456 31696
rect 32416 31414 32444 31690
rect 32404 31408 32456 31414
rect 32404 31350 32456 31356
rect 32220 31204 32272 31210
rect 32220 31146 32272 31152
rect 32404 30184 32456 30190
rect 32404 30126 32456 30132
rect 32036 29844 32088 29850
rect 32036 29786 32088 29792
rect 31944 29572 31996 29578
rect 31944 29514 31996 29520
rect 31484 29504 31536 29510
rect 31484 29446 31536 29452
rect 31576 29504 31628 29510
rect 31852 29504 31904 29510
rect 31576 29446 31628 29452
rect 31666 29472 31722 29481
rect 31482 29200 31538 29209
rect 31482 29135 31484 29144
rect 31536 29135 31538 29144
rect 31484 29106 31536 29112
rect 31392 28144 31444 28150
rect 31392 28086 31444 28092
rect 31404 27849 31432 28086
rect 31390 27840 31446 27849
rect 31390 27775 31446 27784
rect 31484 27600 31536 27606
rect 31484 27542 31536 27548
rect 31496 27130 31524 27542
rect 31484 27124 31536 27130
rect 31484 27066 31536 27072
rect 31588 26926 31616 29446
rect 31852 29446 31904 29452
rect 31666 29407 31722 29416
rect 31680 29170 31708 29407
rect 31668 29164 31720 29170
rect 31668 29106 31720 29112
rect 31956 29034 31984 29514
rect 31944 29028 31996 29034
rect 31944 28970 31996 28976
rect 31852 28484 31904 28490
rect 31852 28426 31904 28432
rect 31668 28416 31720 28422
rect 31668 28358 31720 28364
rect 31680 27674 31708 28358
rect 31864 28150 31892 28426
rect 31852 28144 31904 28150
rect 31852 28086 31904 28092
rect 31852 27872 31904 27878
rect 31852 27814 31904 27820
rect 31668 27668 31720 27674
rect 31668 27610 31720 27616
rect 31864 27470 31892 27814
rect 31852 27464 31904 27470
rect 31852 27406 31904 27412
rect 31668 26988 31720 26994
rect 31668 26930 31720 26936
rect 31576 26920 31628 26926
rect 31680 26897 31708 26930
rect 31576 26862 31628 26868
rect 31666 26888 31722 26897
rect 31666 26823 31722 26832
rect 31576 26580 31628 26586
rect 31680 26568 31708 26823
rect 31628 26540 31708 26568
rect 31760 26580 31812 26586
rect 31576 26522 31628 26528
rect 31760 26522 31812 26528
rect 31298 24984 31354 24993
rect 31298 24919 31354 24928
rect 31772 24410 31800 26522
rect 31864 26382 31892 27406
rect 31852 26376 31904 26382
rect 31852 26318 31904 26324
rect 31956 26246 31984 28970
rect 32048 28558 32076 29786
rect 32312 29504 32364 29510
rect 32312 29446 32364 29452
rect 32036 28552 32088 28558
rect 32036 28494 32088 28500
rect 32324 28082 32352 29446
rect 32416 28082 32444 30126
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32404 28076 32456 28082
rect 32404 28018 32456 28024
rect 32036 26852 32088 26858
rect 32036 26794 32088 26800
rect 32048 26314 32076 26794
rect 32128 26580 32180 26586
rect 32180 26540 32260 26568
rect 32128 26522 32180 26528
rect 32128 26444 32180 26450
rect 32128 26386 32180 26392
rect 32036 26308 32088 26314
rect 32036 26250 32088 26256
rect 31944 26240 31996 26246
rect 31944 26182 31996 26188
rect 31956 24750 31984 26182
rect 32140 26042 32168 26386
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 32036 25900 32088 25906
rect 32036 25842 32088 25848
rect 32048 25537 32076 25842
rect 32128 25764 32180 25770
rect 32128 25706 32180 25712
rect 32034 25528 32090 25537
rect 32034 25463 32090 25472
rect 32140 25430 32168 25706
rect 32128 25424 32180 25430
rect 32232 25401 32260 26540
rect 32416 26450 32444 28018
rect 32508 26790 32536 33934
rect 32864 33856 32916 33862
rect 32864 33798 32916 33804
rect 32876 33590 32904 33798
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 32864 33584 32916 33590
rect 32864 33526 32916 33532
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 33416 32904 33468 32910
rect 33416 32846 33468 32852
rect 33428 32570 33456 32846
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 33416 32564 33468 32570
rect 33416 32506 33468 32512
rect 32680 32496 32732 32502
rect 32680 32438 32732 32444
rect 34426 32464 34482 32473
rect 32588 32428 32640 32434
rect 32588 32370 32640 32376
rect 32600 32337 32628 32370
rect 32586 32328 32642 32337
rect 32586 32263 32642 32272
rect 32586 32056 32642 32065
rect 32586 31991 32588 32000
rect 32640 31991 32642 32000
rect 32588 31962 32640 31968
rect 32692 31822 32720 32438
rect 32772 32428 32824 32434
rect 34426 32399 34482 32408
rect 32772 32370 32824 32376
rect 32784 31958 32812 32370
rect 32864 32224 32916 32230
rect 32864 32166 32916 32172
rect 32772 31952 32824 31958
rect 32772 31894 32824 31900
rect 32680 31816 32732 31822
rect 32680 31758 32732 31764
rect 32588 31680 32640 31686
rect 32588 31622 32640 31628
rect 32600 31346 32628 31622
rect 32692 31482 32720 31758
rect 32680 31476 32732 31482
rect 32680 31418 32732 31424
rect 32784 31414 32812 31894
rect 32772 31408 32824 31414
rect 32772 31350 32824 31356
rect 32588 31340 32640 31346
rect 32588 31282 32640 31288
rect 32680 31340 32732 31346
rect 32680 31282 32732 31288
rect 32692 29306 32720 31282
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 32692 28626 32720 29242
rect 32680 28620 32732 28626
rect 32680 28562 32732 28568
rect 32680 28076 32732 28082
rect 32680 28018 32732 28024
rect 32692 27062 32720 28018
rect 32680 27056 32732 27062
rect 32680 26998 32732 27004
rect 32496 26784 32548 26790
rect 32496 26726 32548 26732
rect 32508 26466 32536 26726
rect 32404 26444 32456 26450
rect 32508 26438 32628 26466
rect 32404 26386 32456 26392
rect 32404 26240 32456 26246
rect 32404 26182 32456 26188
rect 32312 26036 32364 26042
rect 32312 25978 32364 25984
rect 32324 25945 32352 25978
rect 32310 25936 32366 25945
rect 32310 25871 32366 25880
rect 32128 25366 32180 25372
rect 32218 25392 32274 25401
rect 32036 25356 32088 25362
rect 32218 25327 32274 25336
rect 32324 25344 32352 25871
rect 32416 25770 32444 26182
rect 32600 26042 32628 26438
rect 32680 26444 32732 26450
rect 32680 26386 32732 26392
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 32404 25764 32456 25770
rect 32404 25706 32456 25712
rect 32324 25316 32444 25344
rect 32036 25298 32088 25304
rect 32048 24954 32076 25298
rect 32236 25266 32288 25272
rect 32128 25220 32180 25226
rect 32416 25242 32444 25316
rect 32496 25254 32548 25260
rect 32288 25214 32352 25242
rect 32416 25214 32496 25242
rect 32236 25208 32288 25214
rect 32128 25162 32180 25168
rect 32036 24948 32088 24954
rect 32036 24890 32088 24896
rect 31944 24744 31996 24750
rect 31944 24686 31996 24692
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 31852 24336 31904 24342
rect 31482 24304 31538 24313
rect 31852 24278 31904 24284
rect 31482 24239 31538 24248
rect 31760 24268 31812 24274
rect 31300 24132 31352 24138
rect 31300 24074 31352 24080
rect 31312 23769 31340 24074
rect 31298 23760 31354 23769
rect 31496 23730 31524 24239
rect 31760 24210 31812 24216
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 31588 24070 31616 24142
rect 31576 24064 31628 24070
rect 31576 24006 31628 24012
rect 31298 23695 31354 23704
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31300 23656 31352 23662
rect 31300 23598 31352 23604
rect 31312 22137 31340 23598
rect 31298 22128 31354 22137
rect 31298 22063 31354 22072
rect 31208 21616 31260 21622
rect 31208 21558 31260 21564
rect 31208 21412 31260 21418
rect 31208 21354 31260 21360
rect 31220 21010 31248 21354
rect 31208 21004 31260 21010
rect 31208 20946 31260 20952
rect 31116 20460 31168 20466
rect 31116 20402 31168 20408
rect 31024 19984 31076 19990
rect 31024 19926 31076 19932
rect 31036 16114 31064 19926
rect 31024 16108 31076 16114
rect 31024 16050 31076 16056
rect 31024 15904 31076 15910
rect 31024 15846 31076 15852
rect 31036 15502 31064 15846
rect 31024 15496 31076 15502
rect 31024 15438 31076 15444
rect 31128 14464 31156 20402
rect 31220 20262 31248 20946
rect 31496 20942 31524 23666
rect 31772 23526 31800 24210
rect 31864 23866 31892 24278
rect 31852 23860 31904 23866
rect 31852 23802 31904 23808
rect 31760 23520 31812 23526
rect 31760 23462 31812 23468
rect 31864 22642 31892 23802
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31668 21072 31720 21078
rect 31668 21014 31720 21020
rect 31680 20942 31708 21014
rect 31956 20942 31984 24686
rect 32140 23866 32168 25162
rect 32218 25120 32274 25129
rect 32218 25055 32274 25064
rect 32128 23860 32180 23866
rect 32128 23802 32180 23808
rect 32128 22160 32180 22166
rect 32128 22102 32180 22108
rect 31484 20936 31536 20942
rect 31484 20878 31536 20884
rect 31668 20936 31720 20942
rect 31668 20878 31720 20884
rect 31944 20936 31996 20942
rect 31944 20878 31996 20884
rect 31300 20800 31352 20806
rect 31300 20742 31352 20748
rect 31312 20466 31340 20742
rect 31300 20460 31352 20466
rect 31300 20402 31352 20408
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 31404 20058 31432 20402
rect 31392 20052 31444 20058
rect 31392 19994 31444 20000
rect 31298 19408 31354 19417
rect 31298 19343 31354 19352
rect 31208 18080 31260 18086
rect 31208 18022 31260 18028
rect 31220 17134 31248 18022
rect 31208 17128 31260 17134
rect 31208 17070 31260 17076
rect 31312 16522 31340 19343
rect 31496 18034 31524 20878
rect 31576 18420 31628 18426
rect 31576 18362 31628 18368
rect 31404 18006 31524 18034
rect 31300 16516 31352 16522
rect 31300 16458 31352 16464
rect 31208 15700 31260 15706
rect 31208 15642 31260 15648
rect 31220 15502 31248 15642
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31404 14890 31432 18006
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 31496 17202 31524 17818
rect 31484 17196 31536 17202
rect 31484 17138 31536 17144
rect 31496 16182 31524 17138
rect 31588 17082 31616 18362
rect 31680 17882 31708 20878
rect 32036 20868 32088 20874
rect 32036 20810 32088 20816
rect 31852 18420 31904 18426
rect 31852 18362 31904 18368
rect 31668 17876 31720 17882
rect 31668 17818 31720 17824
rect 31668 17740 31720 17746
rect 31668 17682 31720 17688
rect 31680 17202 31708 17682
rect 31864 17202 31892 18362
rect 31944 18148 31996 18154
rect 31944 18090 31996 18096
rect 31668 17196 31720 17202
rect 31668 17138 31720 17144
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 31864 17082 31892 17138
rect 31588 17054 31892 17082
rect 31956 17066 31984 18090
rect 32048 17338 32076 20810
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 32036 17128 32088 17134
rect 32036 17070 32088 17076
rect 31944 17060 31996 17066
rect 31484 16176 31536 16182
rect 31484 16118 31536 16124
rect 31772 16114 31800 17054
rect 31944 17002 31996 17008
rect 32048 16402 32076 17070
rect 32140 16538 32168 22102
rect 32232 17202 32260 25055
rect 32324 17202 32352 25214
rect 32496 25196 32548 25202
rect 32600 24954 32628 25842
rect 32588 24948 32640 24954
rect 32588 24890 32640 24896
rect 32404 23860 32456 23866
rect 32404 23802 32456 23808
rect 32416 17354 32444 23802
rect 32600 23322 32628 24890
rect 32588 23316 32640 23322
rect 32588 23258 32640 23264
rect 32692 22930 32720 26386
rect 32876 25974 32904 32166
rect 33324 31340 33376 31346
rect 33324 31282 33376 31288
rect 33048 31136 33100 31142
rect 33048 31078 33100 31084
rect 33140 31136 33192 31142
rect 33140 31078 33192 31084
rect 33060 30258 33088 31078
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 32956 29640 33008 29646
rect 32956 29582 33008 29588
rect 32968 27878 32996 29582
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 32864 25968 32916 25974
rect 32864 25910 32916 25916
rect 32770 25528 32826 25537
rect 32770 25463 32826 25472
rect 32784 25294 32812 25463
rect 32772 25288 32824 25294
rect 32772 25230 32824 25236
rect 32864 23656 32916 23662
rect 32864 23598 32916 23604
rect 32772 23520 32824 23526
rect 32772 23462 32824 23468
rect 32600 22902 32720 22930
rect 32600 22778 32628 22902
rect 32588 22772 32640 22778
rect 32588 22714 32640 22720
rect 32680 22772 32732 22778
rect 32680 22714 32732 22720
rect 32600 20534 32628 22714
rect 32692 22166 32720 22714
rect 32784 22642 32812 23462
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 32680 22160 32732 22166
rect 32680 22102 32732 22108
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32784 21146 32812 21490
rect 32772 21140 32824 21146
rect 32772 21082 32824 21088
rect 32588 20528 32640 20534
rect 32588 20470 32640 20476
rect 32784 19378 32812 21082
rect 32876 19394 32904 23598
rect 32968 20754 32996 27814
rect 33152 26994 33180 31078
rect 33336 30258 33364 31282
rect 34058 30424 34114 30433
rect 34058 30359 34114 30368
rect 33324 30252 33376 30258
rect 33324 30194 33376 30200
rect 33416 30252 33468 30258
rect 33416 30194 33468 30200
rect 33232 30116 33284 30122
rect 33232 30058 33284 30064
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 33140 26308 33192 26314
rect 33140 26250 33192 26256
rect 33048 25492 33100 25498
rect 33048 25434 33100 25440
rect 33060 23662 33088 25434
rect 33048 23656 33100 23662
rect 33048 23598 33100 23604
rect 33152 23526 33180 26250
rect 33140 23520 33192 23526
rect 33140 23462 33192 23468
rect 33048 22704 33100 22710
rect 33048 22646 33100 22652
rect 33060 20942 33088 22646
rect 33152 21078 33180 23462
rect 33244 22094 33272 30058
rect 33336 28914 33364 30194
rect 33428 29073 33456 30194
rect 33600 30048 33652 30054
rect 33600 29990 33652 29996
rect 33414 29064 33470 29073
rect 33414 28999 33470 29008
rect 33336 28886 33456 28914
rect 33324 28688 33376 28694
rect 33324 28630 33376 28636
rect 33336 28150 33364 28630
rect 33324 28144 33376 28150
rect 33324 28086 33376 28092
rect 33336 26314 33364 28086
rect 33324 26308 33376 26314
rect 33324 26250 33376 26256
rect 33324 25900 33376 25906
rect 33324 25842 33376 25848
rect 33336 25498 33364 25842
rect 33324 25492 33376 25498
rect 33324 25434 33376 25440
rect 33428 24138 33456 28886
rect 33508 27328 33560 27334
rect 33508 27270 33560 27276
rect 33520 26042 33548 27270
rect 33508 26036 33560 26042
rect 33508 25978 33560 25984
rect 33520 25702 33548 25978
rect 33508 25696 33560 25702
rect 33508 25638 33560 25644
rect 33612 25498 33640 29990
rect 33784 29164 33836 29170
rect 33784 29106 33836 29112
rect 33796 28558 33824 29106
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33968 26988 34020 26994
rect 33968 26930 34020 26936
rect 33980 26382 34008 26930
rect 33968 26376 34020 26382
rect 33968 26318 34020 26324
rect 33784 26240 33836 26246
rect 33784 26182 33836 26188
rect 33600 25492 33652 25498
rect 33600 25434 33652 25440
rect 33416 24132 33468 24138
rect 33416 24074 33468 24080
rect 33612 22094 33640 25434
rect 33796 25294 33824 26182
rect 33980 25906 34008 26318
rect 34072 25906 34100 30359
rect 34440 30274 34468 32399
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 36268 30728 36320 30734
rect 36268 30670 36320 30676
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 34164 30258 34468 30274
rect 34164 30252 34480 30258
rect 34164 30246 34428 30252
rect 34164 26382 34192 30246
rect 34428 30194 34480 30200
rect 34336 30184 34388 30190
rect 34336 30126 34388 30132
rect 34348 28994 34376 30126
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 36176 29232 36228 29238
rect 36176 29174 36228 29180
rect 35808 29164 35860 29170
rect 35808 29106 35860 29112
rect 34520 29096 34572 29102
rect 34520 29038 34572 29044
rect 34796 29096 34848 29102
rect 35820 29073 35848 29106
rect 34796 29038 34848 29044
rect 35806 29064 35862 29073
rect 34348 28966 34468 28994
rect 34440 28694 34468 28966
rect 34428 28688 34480 28694
rect 34428 28630 34480 28636
rect 34440 27062 34468 28630
rect 34428 27056 34480 27062
rect 34428 26998 34480 27004
rect 34152 26376 34204 26382
rect 34152 26318 34204 26324
rect 33968 25900 34020 25906
rect 33968 25842 34020 25848
rect 34060 25900 34112 25906
rect 34060 25842 34112 25848
rect 33876 25832 33928 25838
rect 33876 25774 33928 25780
rect 33692 25288 33744 25294
rect 33692 25230 33744 25236
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33704 24614 33732 25230
rect 33692 24608 33744 24614
rect 33692 24550 33744 24556
rect 33692 22432 33744 22438
rect 33692 22374 33744 22380
rect 33244 22066 33364 22094
rect 33336 22030 33364 22066
rect 33520 22066 33640 22094
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 33140 21072 33192 21078
rect 33140 21014 33192 21020
rect 33048 20936 33100 20942
rect 33048 20878 33100 20884
rect 32968 20726 33180 20754
rect 32772 19372 32824 19378
rect 32876 19366 33088 19394
rect 32772 19314 32824 19320
rect 32864 19304 32916 19310
rect 32864 19246 32916 19252
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 32876 18834 32904 19246
rect 32864 18828 32916 18834
rect 32864 18770 32916 18776
rect 32968 18408 32996 19246
rect 32876 18380 32996 18408
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32784 17678 32812 18226
rect 32772 17672 32824 17678
rect 32772 17614 32824 17620
rect 32416 17326 32628 17354
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 32312 17196 32364 17202
rect 32312 17138 32364 17144
rect 32496 17196 32548 17202
rect 32496 17138 32548 17144
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 32324 16658 32352 16934
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32140 16510 32444 16538
rect 32048 16374 32260 16402
rect 32036 16244 32088 16250
rect 32036 16186 32088 16192
rect 31760 16108 31812 16114
rect 31760 16050 31812 16056
rect 31484 16040 31536 16046
rect 31484 15982 31536 15988
rect 31576 16040 31628 16046
rect 31576 15982 31628 15988
rect 31392 14884 31444 14890
rect 31392 14826 31444 14832
rect 31128 14436 31340 14464
rect 31208 14340 31260 14346
rect 31208 14282 31260 14288
rect 31220 14006 31248 14282
rect 31208 14000 31260 14006
rect 31208 13942 31260 13948
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30932 13796 30984 13802
rect 30932 13738 30984 13744
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30840 12242 30892 12248
rect 30840 12184 30892 12190
rect 30852 11257 30880 12184
rect 30944 11937 30972 13738
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31024 13252 31076 13258
rect 31024 13194 31076 13200
rect 31036 12238 31064 13194
rect 31024 12232 31076 12238
rect 31024 12174 31076 12180
rect 30930 11928 30986 11937
rect 31036 11898 31064 12174
rect 30930 11863 30986 11872
rect 31024 11892 31076 11898
rect 30838 11248 30894 11257
rect 30838 11183 30894 11192
rect 30760 10798 30880 10826
rect 30748 10736 30800 10742
rect 30748 10678 30800 10684
rect 30760 9178 30788 10678
rect 30852 9353 30880 10798
rect 30944 9450 30972 11863
rect 31024 11834 31076 11840
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 31036 11529 31064 11698
rect 31022 11520 31078 11529
rect 31022 11455 31078 11464
rect 31128 10742 31156 13670
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31116 10736 31168 10742
rect 31116 10678 31168 10684
rect 31220 10418 31248 12038
rect 31312 11286 31340 14436
rect 31404 14346 31432 14826
rect 31392 14340 31444 14346
rect 31392 14282 31444 14288
rect 31496 13734 31524 15982
rect 31588 15609 31616 15982
rect 31668 15972 31720 15978
rect 31668 15914 31720 15920
rect 31574 15600 31630 15609
rect 31574 15535 31576 15544
rect 31628 15535 31630 15544
rect 31576 15506 31628 15512
rect 31484 13728 31536 13734
rect 31484 13670 31536 13676
rect 31392 13524 31444 13530
rect 31392 13466 31444 13472
rect 31404 11762 31432 13466
rect 31588 13394 31616 15506
rect 31680 15502 31708 15914
rect 31772 15570 31800 16050
rect 31760 15564 31812 15570
rect 31760 15506 31812 15512
rect 31668 15496 31720 15502
rect 31668 15438 31720 15444
rect 31680 14414 31708 15438
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31772 15026 31800 15302
rect 31852 15088 31904 15094
rect 31852 15030 31904 15036
rect 31760 15020 31812 15026
rect 31760 14962 31812 14968
rect 31668 14408 31720 14414
rect 31668 14350 31720 14356
rect 31680 14056 31708 14350
rect 31680 14028 31800 14056
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31576 13388 31628 13394
rect 31576 13330 31628 13336
rect 31484 13184 31536 13190
rect 31484 13126 31536 13132
rect 31496 12102 31524 13126
rect 31574 13016 31630 13025
rect 31574 12951 31630 12960
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31588 11937 31616 12951
rect 31680 12442 31708 13874
rect 31772 13870 31800 14028
rect 31760 13864 31812 13870
rect 31760 13806 31812 13812
rect 31772 13258 31800 13806
rect 31864 13462 31892 15030
rect 31852 13456 31904 13462
rect 31852 13398 31904 13404
rect 31760 13252 31812 13258
rect 31760 13194 31812 13200
rect 31668 12436 31720 12442
rect 31864 12424 31892 13398
rect 32048 12434 32076 16186
rect 32126 15192 32182 15201
rect 32126 15127 32128 15136
rect 32180 15127 32182 15136
rect 32128 15098 32180 15104
rect 31668 12378 31720 12384
rect 31772 12396 31892 12424
rect 31956 12406 32076 12434
rect 31574 11928 31630 11937
rect 31772 11898 31800 12396
rect 31956 12322 31984 12406
rect 31864 12294 31984 12322
rect 31760 11892 31812 11898
rect 31574 11863 31630 11872
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31588 11642 31616 11863
rect 31496 11614 31616 11642
rect 31680 11852 31760 11880
rect 31390 11520 31446 11529
rect 31390 11455 31446 11464
rect 31300 11280 31352 11286
rect 31300 11222 31352 11228
rect 31312 10577 31340 11222
rect 31404 11150 31432 11455
rect 31392 11144 31444 11150
rect 31392 11086 31444 11092
rect 31298 10568 31354 10577
rect 31298 10503 31354 10512
rect 31390 10432 31446 10441
rect 31220 10390 31340 10418
rect 31206 10296 31262 10305
rect 31206 10231 31208 10240
rect 31260 10231 31262 10240
rect 31208 10202 31260 10208
rect 31312 10198 31340 10390
rect 31390 10367 31446 10376
rect 31300 10192 31352 10198
rect 31300 10134 31352 10140
rect 31024 10056 31076 10062
rect 31024 9998 31076 10004
rect 31036 9722 31064 9998
rect 31024 9716 31076 9722
rect 31024 9658 31076 9664
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 30932 9444 30984 9450
rect 30932 9386 30984 9392
rect 30838 9344 30894 9353
rect 30838 9279 30894 9288
rect 30748 9172 30800 9178
rect 30748 9114 30800 9120
rect 30668 8860 30788 8888
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30668 7274 30696 7686
rect 30656 7268 30708 7274
rect 30656 7210 30708 7216
rect 30564 6656 30616 6662
rect 30564 6598 30616 6604
rect 30484 6446 30696 6474
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30576 5914 30604 6258
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30196 5840 30248 5846
rect 30196 5782 30248 5788
rect 30576 5710 30604 5850
rect 30668 5846 30696 6446
rect 30760 6254 30788 8860
rect 30852 8401 30880 9279
rect 30932 8560 30984 8566
rect 30930 8528 30932 8537
rect 30984 8528 30986 8537
rect 30930 8463 30986 8472
rect 30838 8392 30894 8401
rect 30838 8327 30894 8336
rect 30840 7948 30892 7954
rect 30840 7890 30892 7896
rect 30852 7410 30880 7890
rect 30932 7880 30984 7886
rect 30932 7822 30984 7828
rect 30944 7546 30972 7822
rect 31036 7818 31064 9522
rect 31024 7812 31076 7818
rect 31024 7754 31076 7760
rect 31312 7546 31340 10134
rect 31404 10130 31432 10367
rect 31392 10124 31444 10130
rect 31392 10066 31444 10072
rect 31404 9926 31432 10066
rect 31392 9920 31444 9926
rect 31392 9862 31444 9868
rect 31392 9580 31444 9586
rect 31392 9522 31444 9528
rect 31404 9489 31432 9522
rect 31390 9480 31446 9489
rect 31390 9415 31446 9424
rect 31404 9382 31432 9415
rect 31392 9376 31444 9382
rect 31392 9318 31444 9324
rect 31496 9178 31524 11614
rect 31680 11506 31708 11852
rect 31760 11834 31812 11840
rect 31588 11478 31708 11506
rect 31588 11082 31616 11478
rect 31666 11384 31722 11393
rect 31666 11319 31722 11328
rect 31760 11348 31812 11354
rect 31680 11286 31708 11319
rect 31760 11290 31812 11296
rect 31668 11280 31720 11286
rect 31668 11222 31720 11228
rect 31576 11076 31628 11082
rect 31576 11018 31628 11024
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 31680 10810 31708 11018
rect 31772 10996 31800 11290
rect 31864 11257 31892 12294
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 31944 12164 31996 12170
rect 31944 12106 31996 12112
rect 31850 11248 31906 11257
rect 31956 11218 31984 12106
rect 32034 11656 32090 11665
rect 32034 11591 32090 11600
rect 31850 11183 31906 11192
rect 31944 11212 31996 11218
rect 31944 11154 31996 11160
rect 32048 11150 32076 11591
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 31852 11008 31904 11014
rect 31772 10968 31852 10996
rect 31668 10804 31720 10810
rect 31668 10746 31720 10752
rect 31668 10668 31720 10674
rect 31668 10610 31720 10616
rect 31576 10600 31628 10606
rect 31576 10542 31628 10548
rect 31588 10198 31616 10542
rect 31680 10266 31708 10610
rect 31772 10538 31800 10968
rect 31852 10950 31904 10956
rect 32034 10976 32090 10985
rect 32034 10911 32090 10920
rect 31760 10532 31812 10538
rect 31760 10474 31812 10480
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 31576 10192 31628 10198
rect 31576 10134 31628 10140
rect 31588 9586 31616 10134
rect 31576 9580 31628 9586
rect 31576 9522 31628 9528
rect 31680 9489 31708 10202
rect 31944 10124 31996 10130
rect 31944 10066 31996 10072
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31772 9518 31800 9998
rect 31852 9648 31904 9654
rect 31852 9590 31904 9596
rect 31760 9512 31812 9518
rect 31666 9480 31722 9489
rect 31760 9454 31812 9460
rect 31666 9415 31722 9424
rect 31484 9172 31536 9178
rect 31484 9114 31536 9120
rect 31864 8498 31892 9590
rect 31956 9110 31984 10066
rect 31944 9104 31996 9110
rect 31944 9046 31996 9052
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 31852 8492 31904 8498
rect 31852 8434 31904 8440
rect 31852 7812 31904 7818
rect 31956 7800 31984 8910
rect 32048 8906 32076 10911
rect 32140 10062 32168 12174
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32232 9722 32260 16374
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32324 14346 32352 14962
rect 32312 14340 32364 14346
rect 32312 14282 32364 14288
rect 32324 13326 32352 14282
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 32416 12434 32444 16510
rect 32508 14074 32536 17138
rect 32600 16250 32628 17326
rect 32588 16244 32640 16250
rect 32588 16186 32640 16192
rect 32784 16130 32812 17614
rect 32600 16102 32812 16130
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 32508 13870 32536 14010
rect 32496 13864 32548 13870
rect 32496 13806 32548 13812
rect 32494 13424 32550 13433
rect 32494 13359 32496 13368
rect 32548 13359 32550 13368
rect 32496 13330 32548 13336
rect 32416 12406 32536 12434
rect 32312 12300 32364 12306
rect 32312 12242 32364 12248
rect 32324 11642 32352 12242
rect 32404 11688 32456 11694
rect 32324 11636 32404 11642
rect 32324 11630 32456 11636
rect 32324 11614 32444 11630
rect 32324 11150 32352 11614
rect 32402 11520 32458 11529
rect 32402 11455 32458 11464
rect 32416 11286 32444 11455
rect 32404 11280 32456 11286
rect 32404 11222 32456 11228
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32220 9716 32272 9722
rect 32220 9658 32272 9664
rect 32324 9602 32352 11086
rect 32402 10976 32458 10985
rect 32402 10911 32458 10920
rect 32416 10810 32444 10911
rect 32404 10804 32456 10810
rect 32404 10746 32456 10752
rect 32404 10668 32456 10674
rect 32404 10610 32456 10616
rect 32416 10130 32444 10610
rect 32508 10146 32536 12406
rect 32600 11354 32628 16102
rect 32772 15700 32824 15706
rect 32772 15642 32824 15648
rect 32784 15162 32812 15642
rect 32876 15638 32904 18380
rect 32956 18284 33008 18290
rect 32956 18226 33008 18232
rect 32968 18193 32996 18226
rect 32954 18184 33010 18193
rect 32954 18119 33010 18128
rect 32956 17332 33008 17338
rect 32956 17274 33008 17280
rect 32968 15638 32996 17274
rect 32864 15632 32916 15638
rect 32864 15574 32916 15580
rect 32956 15632 33008 15638
rect 32956 15574 33008 15580
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 32772 15156 32824 15162
rect 32772 15098 32824 15104
rect 32680 15088 32732 15094
rect 32680 15030 32732 15036
rect 32692 12850 32720 15030
rect 32784 13938 32812 15098
rect 32968 15026 32996 15438
rect 32956 15020 33008 15026
rect 32956 14962 33008 14968
rect 32772 13932 32824 13938
rect 32772 13874 32824 13880
rect 32968 13326 32996 14962
rect 32956 13320 33008 13326
rect 32956 13262 33008 13268
rect 32772 13252 32824 13258
rect 32772 13194 32824 13200
rect 32864 13252 32916 13258
rect 32864 13194 32916 13200
rect 32680 12844 32732 12850
rect 32680 12786 32732 12792
rect 32680 12640 32732 12646
rect 32680 12582 32732 12588
rect 32692 12209 32720 12582
rect 32678 12200 32734 12209
rect 32678 12135 32734 12144
rect 32784 11898 32812 13194
rect 32876 12986 32904 13194
rect 32864 12980 32916 12986
rect 32864 12922 32916 12928
rect 32864 12844 32916 12850
rect 32864 12786 32916 12792
rect 32876 12306 32904 12786
rect 32864 12300 32916 12306
rect 32864 12242 32916 12248
rect 32968 12050 32996 13262
rect 33060 12238 33088 19366
rect 33152 15570 33180 20726
rect 33232 18760 33284 18766
rect 33232 18702 33284 18708
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 33140 15428 33192 15434
rect 33140 15370 33192 15376
rect 33048 12232 33100 12238
rect 33048 12174 33100 12180
rect 32876 12022 32996 12050
rect 32876 11898 32904 12022
rect 32954 11928 33010 11937
rect 32772 11892 32824 11898
rect 32772 11834 32824 11840
rect 32864 11892 32916 11898
rect 32954 11863 33010 11872
rect 32864 11834 32916 11840
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 32404 10124 32456 10130
rect 32508 10118 32628 10146
rect 32404 10066 32456 10072
rect 32494 10024 32550 10033
rect 32494 9959 32496 9968
rect 32548 9959 32550 9968
rect 32496 9930 32548 9936
rect 32140 9574 32352 9602
rect 32404 9580 32456 9586
rect 32036 8900 32088 8906
rect 32036 8842 32088 8848
rect 31904 7772 31984 7800
rect 31852 7754 31904 7760
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 31300 7540 31352 7546
rect 31300 7482 31352 7488
rect 31864 7410 31892 7754
rect 30840 7404 30892 7410
rect 30840 7346 30892 7352
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31852 7404 31904 7410
rect 31852 7346 31904 7352
rect 30840 7200 30892 7206
rect 30840 7142 30892 7148
rect 30852 6322 30880 7142
rect 31404 6730 31432 7346
rect 31668 7268 31720 7274
rect 31668 7210 31720 7216
rect 31484 7200 31536 7206
rect 31484 7142 31536 7148
rect 31392 6724 31444 6730
rect 31392 6666 31444 6672
rect 30932 6452 30984 6458
rect 30932 6394 30984 6400
rect 30944 6322 30972 6394
rect 31404 6322 31432 6666
rect 30840 6316 30892 6322
rect 30840 6258 30892 6264
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 31392 6316 31444 6322
rect 31392 6258 31444 6264
rect 30748 6248 30800 6254
rect 30748 6190 30800 6196
rect 30852 5846 30880 6258
rect 30656 5840 30708 5846
rect 30656 5782 30708 5788
rect 30840 5840 30892 5846
rect 30840 5782 30892 5788
rect 30564 5704 30616 5710
rect 30564 5646 30616 5652
rect 30104 5636 30156 5642
rect 30104 5578 30156 5584
rect 30668 5234 30696 5782
rect 30944 5778 30972 6258
rect 31496 6186 31524 7142
rect 31680 6662 31708 7210
rect 31668 6656 31720 6662
rect 31668 6598 31720 6604
rect 31680 6390 31708 6598
rect 31668 6384 31720 6390
rect 31668 6326 31720 6332
rect 31484 6180 31536 6186
rect 31484 6122 31536 6128
rect 31496 5846 31524 6122
rect 31942 5944 31998 5953
rect 31942 5879 31944 5888
rect 31996 5879 31998 5888
rect 31944 5850 31996 5856
rect 31484 5840 31536 5846
rect 31484 5782 31536 5788
rect 32140 5778 32168 9574
rect 32404 9522 32456 9528
rect 32416 8974 32444 9522
rect 32494 9480 32550 9489
rect 32494 9415 32550 9424
rect 32404 8968 32456 8974
rect 32404 8910 32456 8916
rect 32310 8392 32366 8401
rect 32310 8327 32366 8336
rect 32220 8016 32272 8022
rect 32220 7958 32272 7964
rect 32232 6254 32260 7958
rect 32324 6390 32352 8327
rect 32508 7206 32536 9415
rect 32600 9382 32628 10118
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 32692 9178 32720 11698
rect 32772 11280 32824 11286
rect 32772 11222 32824 11228
rect 32784 10742 32812 11222
rect 32876 11150 32904 11834
rect 32968 11830 32996 11863
rect 32956 11824 33008 11830
rect 32956 11766 33008 11772
rect 33048 11552 33100 11558
rect 33048 11494 33100 11500
rect 33060 11354 33088 11494
rect 33152 11354 33180 15370
rect 33244 14074 33272 18702
rect 33336 18630 33364 21966
rect 33324 18624 33376 18630
rect 33324 18566 33376 18572
rect 33336 18290 33364 18566
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 33416 16244 33468 16250
rect 33416 16186 33468 16192
rect 33324 14272 33376 14278
rect 33324 14214 33376 14220
rect 33232 14068 33284 14074
rect 33232 14010 33284 14016
rect 33336 14006 33364 14214
rect 33324 14000 33376 14006
rect 33324 13942 33376 13948
rect 33232 13864 33284 13870
rect 33232 13806 33284 13812
rect 33244 13530 33272 13806
rect 33232 13524 33284 13530
rect 33232 13466 33284 13472
rect 33428 12434 33456 16186
rect 33520 14482 33548 22066
rect 33704 20058 33732 22374
rect 33692 20052 33744 20058
rect 33692 19994 33744 20000
rect 33704 18970 33732 19994
rect 33692 18964 33744 18970
rect 33692 18906 33744 18912
rect 33600 18896 33652 18902
rect 33796 18850 33824 25230
rect 33888 20602 33916 25774
rect 33968 25152 34020 25158
rect 33968 25094 34020 25100
rect 33980 24993 34008 25094
rect 33966 24984 34022 24993
rect 33966 24919 34022 24928
rect 33968 23316 34020 23322
rect 33968 23258 34020 23264
rect 33876 20596 33928 20602
rect 33876 20538 33928 20544
rect 33980 20346 34008 23258
rect 33652 18844 33824 18850
rect 33600 18838 33824 18844
rect 33612 18822 33824 18838
rect 33888 20318 34008 20346
rect 33612 18358 33640 18822
rect 33692 18692 33744 18698
rect 33692 18634 33744 18640
rect 33704 18358 33732 18634
rect 33600 18352 33652 18358
rect 33600 18294 33652 18300
rect 33692 18352 33744 18358
rect 33692 18294 33744 18300
rect 33784 18284 33836 18290
rect 33784 18226 33836 18232
rect 33600 16516 33652 16522
rect 33600 16458 33652 16464
rect 33508 14476 33560 14482
rect 33508 14418 33560 14424
rect 33508 14340 33560 14346
rect 33508 14282 33560 14288
rect 33520 12442 33548 14282
rect 33612 13326 33640 16458
rect 33796 14890 33824 18226
rect 33888 16590 33916 20318
rect 33968 20256 34020 20262
rect 33968 20198 34020 20204
rect 33980 19922 34008 20198
rect 33968 19916 34020 19922
rect 33968 19858 34020 19864
rect 33968 19780 34020 19786
rect 33968 19722 34020 19728
rect 33980 19514 34008 19722
rect 33968 19508 34020 19514
rect 33968 19450 34020 19456
rect 33876 16584 33928 16590
rect 33876 16526 33928 16532
rect 33784 14884 33836 14890
rect 33784 14826 33836 14832
rect 33692 14340 33744 14346
rect 33796 14328 33824 14826
rect 33744 14300 33824 14328
rect 33692 14282 33744 14288
rect 33784 14068 33836 14074
rect 33784 14010 33836 14016
rect 33690 13832 33746 13841
rect 33690 13767 33746 13776
rect 33704 13734 33732 13767
rect 33692 13728 33744 13734
rect 33692 13670 33744 13676
rect 33600 13320 33652 13326
rect 33600 13262 33652 13268
rect 33244 12406 33456 12434
rect 33508 12436 33560 12442
rect 33048 11348 33100 11354
rect 33048 11290 33100 11296
rect 33140 11348 33192 11354
rect 33140 11290 33192 11296
rect 32864 11144 32916 11150
rect 32916 11092 33088 11098
rect 32864 11086 33088 11092
rect 32876 11082 33088 11086
rect 32876 11076 33100 11082
rect 32876 11070 33048 11076
rect 33048 11018 33100 11024
rect 32772 10736 32824 10742
rect 32772 10678 32824 10684
rect 32784 10062 32812 10678
rect 32864 10668 32916 10674
rect 32864 10610 32916 10616
rect 32876 10266 32904 10610
rect 32864 10260 32916 10266
rect 32864 10202 32916 10208
rect 32772 10056 32824 10062
rect 32772 9998 32824 10004
rect 32784 9382 32812 9998
rect 33140 9920 33192 9926
rect 33140 9862 33192 9868
rect 33152 9761 33180 9862
rect 33138 9752 33194 9761
rect 33138 9687 33194 9696
rect 33048 9580 33100 9586
rect 33048 9522 33100 9528
rect 32772 9376 32824 9382
rect 32772 9318 32824 9324
rect 32680 9172 32732 9178
rect 32680 9114 32732 9120
rect 32784 8430 32812 9318
rect 32954 8664 33010 8673
rect 33060 8634 33088 9522
rect 33244 8838 33272 12406
rect 33508 12378 33560 12384
rect 33692 12300 33744 12306
rect 33692 12242 33744 12248
rect 33508 10600 33560 10606
rect 33508 10542 33560 10548
rect 33416 10464 33468 10470
rect 33416 10406 33468 10412
rect 33324 9988 33376 9994
rect 33324 9930 33376 9936
rect 33232 8832 33284 8838
rect 33232 8774 33284 8780
rect 32954 8599 33010 8608
rect 33048 8628 33100 8634
rect 32864 8492 32916 8498
rect 32864 8434 32916 8440
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 32876 7886 32904 8434
rect 32968 8430 32996 8599
rect 33048 8570 33100 8576
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 32864 7880 32916 7886
rect 32864 7822 32916 7828
rect 32876 7410 32904 7822
rect 33046 7576 33102 7585
rect 33046 7511 33102 7520
rect 33060 7478 33088 7511
rect 33048 7472 33100 7478
rect 33048 7414 33100 7420
rect 32864 7404 32916 7410
rect 32864 7346 32916 7352
rect 32496 7200 32548 7206
rect 32496 7142 32548 7148
rect 32508 6866 32536 7142
rect 32876 7002 32904 7346
rect 32864 6996 32916 7002
rect 32864 6938 32916 6944
rect 32496 6860 32548 6866
rect 32496 6802 32548 6808
rect 32876 6798 32904 6938
rect 32864 6792 32916 6798
rect 32864 6734 32916 6740
rect 33336 6458 33364 9930
rect 33428 7886 33456 10406
rect 33520 9625 33548 10542
rect 33704 9654 33732 12242
rect 33796 9654 33824 14010
rect 33888 12434 33916 16526
rect 33980 15706 34008 19450
rect 34072 16794 34100 25842
rect 34164 24886 34192 26318
rect 34428 25968 34480 25974
rect 34428 25910 34480 25916
rect 34440 25498 34468 25910
rect 34428 25492 34480 25498
rect 34428 25434 34480 25440
rect 34152 24880 34204 24886
rect 34152 24822 34204 24828
rect 34336 24812 34388 24818
rect 34336 24754 34388 24760
rect 34348 24614 34376 24754
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 34336 24608 34388 24614
rect 34336 24550 34388 24556
rect 34164 23798 34192 24550
rect 34152 23792 34204 23798
rect 34152 23734 34204 23740
rect 34164 19854 34192 23734
rect 34428 23724 34480 23730
rect 34428 23666 34480 23672
rect 34244 21888 34296 21894
rect 34244 21830 34296 21836
rect 34152 19848 34204 19854
rect 34152 19790 34204 19796
rect 34152 19712 34204 19718
rect 34152 19654 34204 19660
rect 34060 16788 34112 16794
rect 34060 16730 34112 16736
rect 33968 15700 34020 15706
rect 33968 15642 34020 15648
rect 34060 14816 34112 14822
rect 34060 14758 34112 14764
rect 34072 14414 34100 14758
rect 34060 14408 34112 14414
rect 34060 14350 34112 14356
rect 33968 13932 34020 13938
rect 34072 13920 34100 14350
rect 34164 13938 34192 19654
rect 34256 15638 34284 21830
rect 34440 19378 34468 23666
rect 34532 20777 34560 29038
rect 34808 28626 34836 29038
rect 35624 29028 35676 29034
rect 35806 28999 35862 29008
rect 35624 28970 35676 28976
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34888 28756 34940 28762
rect 34888 28698 34940 28704
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 34704 28484 34756 28490
rect 34704 28426 34756 28432
rect 34612 28416 34664 28422
rect 34612 28358 34664 28364
rect 34624 27606 34652 28358
rect 34612 27600 34664 27606
rect 34612 27542 34664 27548
rect 34716 26994 34744 28426
rect 34900 27962 34928 28698
rect 35636 28490 35664 28970
rect 35808 28960 35860 28966
rect 35808 28902 35860 28908
rect 35624 28484 35676 28490
rect 35624 28426 35676 28432
rect 35820 28404 35848 28902
rect 35820 28376 36032 28404
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 34808 27934 34928 27962
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 34612 26852 34664 26858
rect 34612 26794 34664 26800
rect 34624 25158 34652 26794
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 34612 25152 34664 25158
rect 34612 25094 34664 25100
rect 34612 23724 34664 23730
rect 34716 23712 34744 25978
rect 34664 23684 34744 23712
rect 34612 23666 34664 23672
rect 34808 23662 34836 27934
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35348 26784 35400 26790
rect 35348 26726 35400 26732
rect 35440 26784 35492 26790
rect 35440 26726 35492 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 24834 35388 26726
rect 35452 25702 35480 26726
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35440 25696 35492 25702
rect 35440 25638 35492 25644
rect 35440 25288 35492 25294
rect 35440 25230 35492 25236
rect 35268 24818 35388 24834
rect 35256 24812 35388 24818
rect 35308 24806 35388 24812
rect 35256 24754 35308 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 23656 34848 23662
rect 35452 23610 35480 25230
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 36004 24954 36032 28376
rect 36084 25832 36136 25838
rect 36084 25774 36136 25780
rect 36096 25226 36124 25774
rect 36084 25220 36136 25226
rect 36084 25162 36136 25168
rect 35992 24948 36044 24954
rect 35992 24890 36044 24896
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 35900 24608 35952 24614
rect 36004 24585 36032 24754
rect 35900 24550 35952 24556
rect 35990 24576 36046 24585
rect 35912 24426 35940 24550
rect 35990 24511 36046 24520
rect 35912 24398 36032 24426
rect 36188 24410 36216 29174
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 34796 23598 34848 23604
rect 34612 23588 34664 23594
rect 34612 23530 34664 23536
rect 35360 23582 35480 23610
rect 34624 22574 34652 23530
rect 34796 23520 34848 23526
rect 34796 23462 34848 23468
rect 34808 22642 34836 23462
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 34796 22636 34848 22642
rect 34796 22578 34848 22584
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 34612 20800 34664 20806
rect 34518 20768 34574 20777
rect 34612 20742 34664 20748
rect 34518 20703 34574 20712
rect 34624 20398 34652 20742
rect 34612 20392 34664 20398
rect 34612 20334 34664 20340
rect 34520 20256 34572 20262
rect 34520 20198 34572 20204
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34336 18352 34388 18358
rect 34336 18294 34388 18300
rect 34348 17882 34376 18294
rect 34532 17882 34560 20198
rect 34612 18080 34664 18086
rect 34612 18022 34664 18028
rect 34336 17876 34388 17882
rect 34336 17818 34388 17824
rect 34520 17876 34572 17882
rect 34520 17818 34572 17824
rect 34624 17354 34652 18022
rect 34532 17326 34652 17354
rect 34244 15632 34296 15638
rect 34532 15586 34560 17326
rect 34716 17184 34744 22578
rect 34796 22432 34848 22438
rect 34796 22374 34848 22380
rect 34808 22030 34836 22374
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35360 22250 35388 23582
rect 35440 23520 35492 23526
rect 35440 23462 35492 23468
rect 35268 22222 35388 22250
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 35268 21457 35296 22222
rect 35348 22160 35400 22166
rect 35348 22102 35400 22108
rect 35254 21448 35310 21457
rect 35254 21383 35310 21392
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 20324 34848 20330
rect 34796 20266 34848 20272
rect 34244 15574 34296 15580
rect 34348 15558 34560 15586
rect 34624 17156 34744 17184
rect 34624 15586 34652 17156
rect 34704 17060 34756 17066
rect 34704 17002 34756 17008
rect 34716 15706 34744 17002
rect 34808 16153 34836 20266
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35256 19916 35308 19922
rect 35256 19858 35308 19864
rect 35268 19281 35296 19858
rect 35254 19272 35310 19281
rect 35254 19207 35310 19216
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18766 35388 22102
rect 35348 18760 35400 18766
rect 35268 18708 35348 18714
rect 35268 18702 35400 18708
rect 35268 18686 35388 18702
rect 35268 18426 35296 18686
rect 35348 18624 35400 18630
rect 35348 18566 35400 18572
rect 35256 18420 35308 18426
rect 35256 18362 35308 18368
rect 35360 18358 35388 18566
rect 35348 18352 35400 18358
rect 35348 18294 35400 18300
rect 35452 18290 35480 23462
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 36004 22030 36032 24398
rect 36176 24404 36228 24410
rect 36176 24346 36228 24352
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 36096 23905 36124 24142
rect 36082 23896 36138 23905
rect 36082 23831 36138 23840
rect 36280 22778 36308 30670
rect 36360 28212 36412 28218
rect 36360 28154 36412 28160
rect 36268 22772 36320 22778
rect 36268 22714 36320 22720
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 36096 22545 36124 22578
rect 36082 22536 36138 22545
rect 36082 22471 36138 22480
rect 35992 22024 36044 22030
rect 35992 21966 36044 21972
rect 36084 22024 36136 22030
rect 36084 21966 36136 21972
rect 36096 21865 36124 21966
rect 36082 21856 36138 21865
rect 35594 21788 35902 21797
rect 36082 21791 36138 21800
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 36084 21548 36136 21554
rect 36084 21490 36136 21496
rect 35806 21448 35862 21457
rect 35806 21383 35862 21392
rect 35820 20913 35848 21383
rect 36096 21185 36124 21490
rect 36082 21176 36138 21185
rect 36082 21111 36138 21120
rect 35806 20904 35862 20913
rect 35806 20839 35862 20848
rect 35820 20788 35848 20839
rect 35820 20760 36032 20788
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35532 20460 35584 20466
rect 35532 20402 35584 20408
rect 35544 19922 35572 20402
rect 35532 19916 35584 19922
rect 35532 19858 35584 19864
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35256 16652 35308 16658
rect 35256 16594 35308 16600
rect 35268 16561 35296 16594
rect 35254 16552 35310 16561
rect 35254 16487 35310 16496
rect 34794 16144 34850 16153
rect 34794 16079 34850 16088
rect 34796 15904 34848 15910
rect 34796 15846 34848 15852
rect 34808 15706 34836 15846
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 15700 34756 15706
rect 34704 15642 34756 15648
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 34624 15570 34744 15586
rect 34612 15564 34744 15570
rect 34244 14544 34296 14550
rect 34244 14486 34296 14492
rect 34020 13892 34100 13920
rect 34152 13932 34204 13938
rect 33968 13874 34020 13880
rect 34152 13874 34204 13880
rect 34060 13456 34112 13462
rect 34060 13398 34112 13404
rect 33888 12406 34008 12434
rect 33876 10192 33928 10198
rect 33876 10134 33928 10140
rect 33888 10062 33916 10134
rect 33876 10056 33928 10062
rect 33876 9998 33928 10004
rect 33692 9648 33744 9654
rect 33506 9616 33562 9625
rect 33692 9590 33744 9596
rect 33784 9648 33836 9654
rect 33784 9590 33836 9596
rect 33506 9551 33508 9560
rect 33560 9551 33562 9560
rect 33508 9522 33560 9528
rect 33520 8634 33548 9522
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33888 8090 33916 9998
rect 33980 9042 34008 12406
rect 34072 12374 34100 13398
rect 34060 12368 34112 12374
rect 34060 12310 34112 12316
rect 34072 12170 34100 12310
rect 34152 12300 34204 12306
rect 34256 12288 34284 14486
rect 34348 14074 34376 15558
rect 34664 15558 34744 15564
rect 34612 15506 34664 15512
rect 34520 15496 34572 15502
rect 34520 15438 34572 15444
rect 34428 15360 34480 15366
rect 34428 15302 34480 15308
rect 34336 14068 34388 14074
rect 34336 14010 34388 14016
rect 34204 12260 34284 12288
rect 34152 12242 34204 12248
rect 34336 12232 34388 12238
rect 34336 12174 34388 12180
rect 34060 12164 34112 12170
rect 34060 12106 34112 12112
rect 34348 11898 34376 12174
rect 34336 11892 34388 11898
rect 34336 11834 34388 11840
rect 34440 10742 34468 15302
rect 34532 14278 34560 15438
rect 34612 15360 34664 15366
rect 34612 15302 34664 15308
rect 34624 14346 34652 15302
rect 34612 14340 34664 14346
rect 34612 14282 34664 14288
rect 34520 14272 34572 14278
rect 34520 14214 34572 14220
rect 34520 14068 34572 14074
rect 34520 14010 34572 14016
rect 34532 13410 34560 14010
rect 34624 13530 34652 14282
rect 34612 13524 34664 13530
rect 34612 13466 34664 13472
rect 34532 13382 34652 13410
rect 34520 13320 34572 13326
rect 34520 13262 34572 13268
rect 34532 11830 34560 13262
rect 34520 11824 34572 11830
rect 34520 11766 34572 11772
rect 34532 11354 34560 11766
rect 34520 11348 34572 11354
rect 34520 11290 34572 11296
rect 34520 11212 34572 11218
rect 34520 11154 34572 11160
rect 34428 10736 34480 10742
rect 34428 10678 34480 10684
rect 34152 10532 34204 10538
rect 34152 10474 34204 10480
rect 34164 9926 34192 10474
rect 34336 10464 34388 10470
rect 34336 10406 34388 10412
rect 34348 10146 34376 10406
rect 34426 10296 34482 10305
rect 34426 10231 34428 10240
rect 34480 10231 34482 10240
rect 34428 10202 34480 10208
rect 34348 10118 34468 10146
rect 34152 9920 34204 9926
rect 34152 9862 34204 9868
rect 34336 9920 34388 9926
rect 34336 9862 34388 9868
rect 34242 9752 34298 9761
rect 34242 9687 34298 9696
rect 34058 9616 34114 9625
rect 34058 9551 34114 9560
rect 33968 9036 34020 9042
rect 33968 8978 34020 8984
rect 33980 8498 34008 8978
rect 33968 8492 34020 8498
rect 33968 8434 34020 8440
rect 33876 8084 33928 8090
rect 33876 8026 33928 8032
rect 33416 7880 33468 7886
rect 33416 7822 33468 7828
rect 33428 6798 33456 7822
rect 33888 6866 33916 8026
rect 33876 6860 33928 6866
rect 33876 6802 33928 6808
rect 33416 6792 33468 6798
rect 33416 6734 33468 6740
rect 33324 6452 33376 6458
rect 33324 6394 33376 6400
rect 32312 6384 32364 6390
rect 32312 6326 32364 6332
rect 33428 6322 33456 6734
rect 33888 6662 33916 6802
rect 33876 6656 33928 6662
rect 33876 6598 33928 6604
rect 33888 6458 33916 6598
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 32864 6316 32916 6322
rect 32864 6258 32916 6264
rect 33416 6316 33468 6322
rect 33416 6258 33468 6264
rect 32220 6248 32272 6254
rect 32220 6190 32272 6196
rect 30932 5772 30984 5778
rect 30932 5714 30984 5720
rect 32128 5772 32180 5778
rect 32128 5714 32180 5720
rect 32232 5710 32260 6190
rect 32876 5710 32904 6258
rect 32220 5704 32272 5710
rect 32220 5646 32272 5652
rect 32864 5704 32916 5710
rect 32864 5646 32916 5652
rect 33428 5642 33456 6258
rect 33888 5710 33916 6394
rect 33876 5704 33928 5710
rect 33876 5646 33928 5652
rect 33416 5636 33468 5642
rect 33416 5578 33468 5584
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 30656 5228 30708 5234
rect 30656 5170 30708 5176
rect 30378 5128 30434 5137
rect 30378 5063 30380 5072
rect 30432 5063 30434 5072
rect 30380 5034 30432 5040
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 27068 3392 27120 3398
rect 27068 3334 27120 3340
rect 34072 3126 34100 9551
rect 34256 9110 34284 9687
rect 34244 9104 34296 9110
rect 34244 9046 34296 9052
rect 34152 8900 34204 8906
rect 34152 8842 34204 8848
rect 34244 8900 34296 8906
rect 34244 8842 34296 8848
rect 34164 8498 34192 8842
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34256 6186 34284 8842
rect 34348 8838 34376 9862
rect 34440 9654 34468 10118
rect 34428 9648 34480 9654
rect 34428 9590 34480 9596
rect 34440 9110 34468 9590
rect 34428 9104 34480 9110
rect 34428 9046 34480 9052
rect 34336 8832 34388 8838
rect 34336 8774 34388 8780
rect 34440 8498 34468 9046
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34440 8242 34468 8434
rect 34532 8430 34560 11154
rect 34624 9042 34652 13382
rect 34716 12442 34744 15558
rect 34808 13734 34836 15642
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35452 14618 35480 18226
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35530 16144 35586 16153
rect 35530 16079 35586 16088
rect 35544 15502 35572 16079
rect 35532 15496 35584 15502
rect 35532 15438 35584 15444
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35256 14612 35308 14618
rect 35256 14554 35308 14560
rect 35440 14612 35492 14618
rect 35440 14554 35492 14560
rect 35070 14512 35126 14521
rect 35070 14447 35126 14456
rect 34980 14272 35032 14278
rect 34980 14214 35032 14220
rect 34992 13734 35020 14214
rect 35084 13938 35112 14447
rect 35072 13932 35124 13938
rect 35072 13874 35124 13880
rect 35268 13870 35296 14554
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 35440 14068 35492 14074
rect 35440 14010 35492 14016
rect 35256 13864 35308 13870
rect 35256 13806 35308 13812
rect 34796 13728 34848 13734
rect 34796 13670 34848 13676
rect 34980 13728 35032 13734
rect 34980 13670 35032 13676
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 13524 34848 13530
rect 34796 13466 34848 13472
rect 35256 13524 35308 13530
rect 35256 13466 35308 13472
rect 34808 12442 34836 13466
rect 35268 12866 35296 13466
rect 35268 12838 35388 12866
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34796 12436 34848 12442
rect 34796 12378 34848 12384
rect 34794 12336 34850 12345
rect 34794 12271 34850 12280
rect 34808 12238 34836 12271
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 34978 12200 35034 12209
rect 34978 12135 34980 12144
rect 35032 12135 35034 12144
rect 34980 12106 35032 12112
rect 34704 11620 34756 11626
rect 34704 11562 34756 11568
rect 34716 11354 34744 11562
rect 34796 11552 34848 11558
rect 34796 11494 34848 11500
rect 34704 11348 34756 11354
rect 34704 11290 34756 11296
rect 34808 11150 34836 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34888 11348 34940 11354
rect 34888 11290 34940 11296
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 34900 10554 34928 11290
rect 34980 11280 35032 11286
rect 34980 11222 35032 11228
rect 35360 11234 35388 12838
rect 35452 11694 35480 14010
rect 36004 13954 36032 20760
rect 36084 16584 36136 16590
rect 36084 16526 36136 16532
rect 35820 13926 36032 13954
rect 35820 13530 35848 13926
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 36096 12209 36124 16526
rect 36082 12200 36138 12209
rect 36082 12135 36138 12144
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 35440 11688 35492 11694
rect 35440 11630 35492 11636
rect 36084 11688 36136 11694
rect 36084 11630 36136 11636
rect 34992 10742 35020 11222
rect 35360 11206 35480 11234
rect 35348 11144 35400 11150
rect 35348 11086 35400 11092
rect 34980 10736 35032 10742
rect 34980 10678 35032 10684
rect 34808 10526 34928 10554
rect 34808 10146 34836 10526
rect 34992 10470 35020 10678
rect 34980 10464 35032 10470
rect 34980 10406 35032 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34808 10118 34928 10146
rect 34704 10056 34756 10062
rect 34704 9998 34756 10004
rect 34716 9722 34744 9998
rect 34796 9988 34848 9994
rect 34796 9930 34848 9936
rect 34704 9716 34756 9722
rect 34704 9658 34756 9664
rect 34808 9568 34836 9930
rect 34900 9674 34928 10118
rect 35164 9988 35216 9994
rect 35164 9930 35216 9936
rect 34900 9646 35112 9674
rect 35176 9654 35204 9930
rect 35360 9897 35388 11086
rect 35452 10130 35480 11206
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 35532 10464 35584 10470
rect 35532 10406 35584 10412
rect 35440 10124 35492 10130
rect 35440 10066 35492 10072
rect 35544 10010 35572 10406
rect 35452 9982 35572 10010
rect 35992 9988 36044 9994
rect 35346 9888 35402 9897
rect 35346 9823 35402 9832
rect 35084 9586 35112 9646
rect 35164 9648 35216 9654
rect 35162 9616 35164 9625
rect 35216 9616 35218 9625
rect 35360 9602 35388 9823
rect 35452 9674 35480 9982
rect 35992 9930 36044 9936
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 35452 9646 35572 9674
rect 35072 9580 35124 9586
rect 34808 9540 35020 9568
rect 34992 9489 35020 9540
rect 35162 9551 35218 9560
rect 35268 9574 35388 9602
rect 35544 9586 35572 9646
rect 35532 9580 35584 9586
rect 35072 9522 35124 9528
rect 34978 9480 35034 9489
rect 35268 9450 35296 9574
rect 35532 9522 35584 9528
rect 35348 9512 35400 9518
rect 35624 9512 35676 9518
rect 35348 9454 35400 9460
rect 35530 9480 35586 9489
rect 34978 9415 35034 9424
rect 35256 9444 35308 9450
rect 35256 9386 35308 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34612 9036 34664 9042
rect 34612 8978 34664 8984
rect 35072 9036 35124 9042
rect 35072 8978 35124 8984
rect 34888 8832 34940 8838
rect 34808 8780 34888 8786
rect 34808 8774 34940 8780
rect 34808 8758 34928 8774
rect 34520 8424 34572 8430
rect 34520 8366 34572 8372
rect 34612 8288 34664 8294
rect 34440 8214 34560 8242
rect 34612 8230 34664 8236
rect 34244 6180 34296 6186
rect 34244 6122 34296 6128
rect 34532 4826 34560 8214
rect 34624 6322 34652 8230
rect 34808 8022 34836 8758
rect 35084 8430 35112 8978
rect 35164 8968 35216 8974
rect 35164 8910 35216 8916
rect 35072 8424 35124 8430
rect 35072 8366 35124 8372
rect 35176 8294 35204 8910
rect 35164 8288 35216 8294
rect 35164 8230 35216 8236
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 8090 35388 9454
rect 35440 9444 35492 9450
rect 35624 9454 35676 9460
rect 35530 9415 35586 9424
rect 35440 9386 35492 9392
rect 35452 8974 35480 9386
rect 35440 8968 35492 8974
rect 35440 8910 35492 8916
rect 35544 8838 35572 9415
rect 35636 8906 35664 9454
rect 35716 9444 35768 9450
rect 35716 9386 35768 9392
rect 35728 9110 35756 9386
rect 35716 9104 35768 9110
rect 35716 9046 35768 9052
rect 35624 8900 35676 8906
rect 35624 8842 35676 8848
rect 35532 8832 35584 8838
rect 35452 8792 35532 8820
rect 35348 8084 35400 8090
rect 35348 8026 35400 8032
rect 34796 8016 34848 8022
rect 34796 7958 34848 7964
rect 34808 6934 34836 7958
rect 35452 7954 35480 8792
rect 35532 8774 35584 8780
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 35440 7948 35492 7954
rect 35440 7890 35492 7896
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6928 34848 6934
rect 34796 6870 34848 6876
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34612 6316 34664 6322
rect 34612 6258 34664 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34520 4820 34572 4826
rect 34520 4762 34572 4768
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36004 3738 36032 9930
rect 36096 8634 36124 11630
rect 36372 9178 36400 28154
rect 36450 27976 36506 27985
rect 36450 27911 36506 27920
rect 36464 21690 36492 27911
rect 36452 21684 36504 21690
rect 36452 21626 36504 21632
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 36084 8628 36136 8634
rect 36084 8570 36136 8576
rect 35992 3732 36044 3738
rect 35992 3674 36044 3680
rect 36084 3528 36136 3534
rect 36082 3496 36084 3505
rect 36136 3496 36138 3505
rect 36082 3431 36138 3440
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 34060 3120 34112 3126
rect 34060 3062 34112 3068
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 23572 2848 23624 2854
rect 23572 2790 23624 2796
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 23584 2514 23612 2790
rect 23676 2514 23704 2790
rect 25148 2650 25176 2926
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 25136 2644 25188 2650
rect 25136 2586 25188 2592
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 18 0 74 800
rect 662 0 718 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 3698 35400 3754 35456
rect 1306 32680 1362 32736
rect 2410 32000 2466 32056
rect 1306 31356 1308 31376
rect 1308 31356 1360 31376
rect 1360 31356 1362 31376
rect 1306 31320 1362 31356
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4342 32836 4398 32872
rect 4342 32816 4344 32836
rect 4344 32816 4396 32836
rect 4396 32816 4398 32836
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4802 32972 4858 33008
rect 4802 32952 4804 32972
rect 4804 32952 4856 32972
rect 4856 32952 4858 32972
rect 5170 32988 5172 33008
rect 5172 32988 5224 33008
rect 5224 32988 5226 33008
rect 5170 32952 5226 32988
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4986 32408 5042 32464
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 3146 30640 3202 30696
rect 1306 29960 1362 30016
rect 1306 29280 1362 29336
rect 1950 29144 2006 29200
rect 1306 28620 1362 28656
rect 1306 28600 1308 28620
rect 1308 28600 1360 28620
rect 1360 28600 1362 28620
rect 1398 27956 1400 27976
rect 1400 27956 1452 27976
rect 1452 27956 1454 27976
rect 1398 27920 1454 27956
rect 3146 24828 3148 24848
rect 3148 24828 3200 24848
rect 3200 24828 3202 24848
rect 3146 24792 3202 24828
rect 2870 23568 2926 23624
rect 2594 16088 2650 16144
rect 2042 12824 2098 12880
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4434 30796 4490 30832
rect 4434 30776 4436 30796
rect 4436 30776 4488 30796
rect 4488 30776 4490 30796
rect 5078 32272 5134 32328
rect 5262 32272 5318 32328
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4526 30640 4582 30696
rect 4986 30660 5042 30696
rect 4986 30640 4988 30660
rect 4988 30640 5040 30660
rect 5040 30640 5042 30660
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 5722 31728 5778 31784
rect 5446 31592 5502 31648
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 5354 29824 5410 29880
rect 6550 33804 6552 33824
rect 6552 33804 6604 33824
rect 6604 33804 6606 33824
rect 6550 33768 6606 33804
rect 6274 32816 6330 32872
rect 6182 32308 6184 32328
rect 6184 32308 6236 32328
rect 6236 32308 6238 32328
rect 6182 32272 6238 32308
rect 6274 31592 6330 31648
rect 5722 31204 5778 31240
rect 5722 31184 5724 31204
rect 5724 31184 5776 31204
rect 5776 31184 5778 31204
rect 5722 30932 5778 30968
rect 5722 30912 5724 30932
rect 5724 30912 5776 30932
rect 5776 30912 5778 30932
rect 5722 29144 5778 29200
rect 5262 28484 5318 28520
rect 5262 28464 5264 28484
rect 5264 28464 5316 28484
rect 5316 28464 5318 28484
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4066 24112 4122 24168
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 5446 24268 5502 24304
rect 5446 24248 5448 24268
rect 5448 24248 5500 24268
rect 5500 24248 5502 24268
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 5354 23740 5356 23760
rect 5356 23740 5408 23760
rect 5408 23740 5410 23760
rect 5354 23704 5410 23740
rect 3790 19760 3846 19816
rect 3882 18808 3938 18864
rect 3330 16532 3332 16552
rect 3332 16532 3384 16552
rect 3384 16532 3386 16552
rect 3330 16496 3386 16532
rect 2226 9968 2282 10024
rect 3698 17584 3754 17640
rect 4250 22924 4252 22944
rect 4252 22924 4304 22944
rect 4304 22924 4306 22944
rect 4250 22888 4306 22924
rect 4434 22752 4490 22808
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 5078 23432 5134 23488
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 5170 23296 5226 23352
rect 5262 23160 5318 23216
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4894 22616 4950 22672
rect 5170 22480 5226 22536
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4618 20884 4620 20904
rect 4620 20884 4672 20904
rect 4672 20884 4674 20904
rect 4618 20848 4674 20884
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3882 16088 3938 16144
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4434 18128 4490 18184
rect 4618 17992 4674 18048
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 5078 20440 5134 20496
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4710 17856 4766 17912
rect 4342 17740 4398 17776
rect 4342 17720 4344 17740
rect 4344 17720 4396 17740
rect 4396 17720 4398 17740
rect 4250 17332 4306 17368
rect 4250 17312 4252 17332
rect 4252 17312 4304 17332
rect 4304 17312 4306 17332
rect 4894 17620 4896 17640
rect 4896 17620 4948 17640
rect 4948 17620 4950 17640
rect 4894 17584 4950 17620
rect 4710 17312 4766 17368
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 5722 25200 5778 25256
rect 5906 27276 5908 27296
rect 5908 27276 5960 27296
rect 5960 27276 5962 27296
rect 5906 27240 5962 27276
rect 6090 25064 6146 25120
rect 6090 24928 6146 24984
rect 6274 28736 6330 28792
rect 5630 22616 5686 22672
rect 5538 22480 5594 22536
rect 5906 23568 5962 23624
rect 6090 23568 6146 23624
rect 5814 22752 5870 22808
rect 5814 22636 5870 22672
rect 5814 22616 5816 22636
rect 5816 22616 5868 22636
rect 5868 22616 5870 22636
rect 6090 22752 6146 22808
rect 5998 22636 6054 22672
rect 5998 22616 6000 22636
rect 6000 22616 6052 22636
rect 6052 22616 6054 22636
rect 5630 20848 5686 20904
rect 5538 19896 5594 19952
rect 5446 17720 5502 17776
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4526 16632 4582 16688
rect 4434 16532 4436 16552
rect 4436 16532 4488 16552
rect 4488 16532 4490 16552
rect 4434 16496 4490 16532
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4618 15136 4674 15192
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 6458 32952 6514 33008
rect 6826 32408 6882 32464
rect 7378 32988 7380 33008
rect 7380 32988 7432 33008
rect 7432 32988 7434 33008
rect 7378 32952 7434 32988
rect 6642 31592 6698 31648
rect 6458 30368 6514 30424
rect 8022 32020 8078 32056
rect 8022 32000 8024 32020
rect 8024 32000 8076 32020
rect 8076 32000 8078 32020
rect 7286 29688 7342 29744
rect 6550 23704 6606 23760
rect 5262 15308 5264 15328
rect 5264 15308 5316 15328
rect 5316 15308 5318 15328
rect 5262 15272 5318 15308
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4618 13776 4674 13832
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4066 12844 4122 12880
rect 4066 12824 4068 12844
rect 4068 12824 4120 12844
rect 4120 12824 4122 12844
rect 3882 12688 3938 12744
rect 6366 22888 6422 22944
rect 6642 23296 6698 23352
rect 6642 22616 6698 22672
rect 7194 27648 7250 27704
rect 7746 27668 7802 27704
rect 7746 27648 7748 27668
rect 7748 27648 7800 27668
rect 7800 27648 7802 27668
rect 8022 27240 8078 27296
rect 7838 25644 7840 25664
rect 7840 25644 7892 25664
rect 7892 25644 7894 25664
rect 7838 25608 7894 25644
rect 7194 23060 7196 23080
rect 7196 23060 7248 23080
rect 7248 23060 7250 23080
rect 7194 23024 7250 23060
rect 7010 20304 7066 20360
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 5446 13232 5502 13288
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4342 12280 4398 12336
rect 4710 12416 4766 12472
rect 3330 10648 3386 10704
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4894 12552 4950 12608
rect 4802 12144 4858 12200
rect 4986 12144 5042 12200
rect 5170 12552 5226 12608
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5262 11872 5318 11928
rect 4894 11756 4950 11792
rect 4894 11736 4896 11756
rect 4896 11736 4948 11756
rect 4948 11736 4950 11756
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4250 10004 4252 10024
rect 4252 10004 4304 10024
rect 4304 10004 4306 10024
rect 4250 9968 4306 10004
rect 3882 9832 3938 9888
rect 3698 9016 3754 9072
rect 5170 11600 5226 11656
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4710 10104 4766 10160
rect 5538 12688 5594 12744
rect 5814 12552 5870 12608
rect 5446 11600 5502 11656
rect 6182 12688 6238 12744
rect 7378 24148 7380 24168
rect 7380 24148 7432 24168
rect 7432 24148 7434 24168
rect 7378 24112 7434 24148
rect 7378 23724 7434 23760
rect 7378 23704 7380 23724
rect 7380 23704 7432 23724
rect 7432 23704 7434 23724
rect 7378 23432 7434 23488
rect 7470 21972 7472 21992
rect 7472 21972 7524 21992
rect 7524 21972 7526 21992
rect 7470 21936 7526 21972
rect 7654 22752 7710 22808
rect 8482 32000 8538 32056
rect 8850 33360 8906 33416
rect 8574 31204 8630 31240
rect 8574 31184 8576 31204
rect 8576 31184 8628 31204
rect 8628 31184 8630 31204
rect 8390 26288 8446 26344
rect 8114 23296 8170 23352
rect 8114 22344 8170 22400
rect 7838 20884 7840 20904
rect 7840 20884 7892 20904
rect 7892 20884 7894 20904
rect 7838 20848 7894 20884
rect 7010 16088 7066 16144
rect 7838 19352 7894 19408
rect 7746 18420 7802 18456
rect 7746 18400 7748 18420
rect 7748 18400 7800 18420
rect 7800 18400 7802 18420
rect 8114 20440 8170 20496
rect 8390 23160 8446 23216
rect 8482 21936 8538 21992
rect 9126 30912 9182 30968
rect 9402 33396 9404 33416
rect 9404 33396 9456 33416
rect 9456 33396 9458 33416
rect 9402 33360 9458 33396
rect 9126 30268 9128 30288
rect 9128 30268 9180 30288
rect 9180 30268 9182 30288
rect 9126 30232 9182 30268
rect 9310 29824 9366 29880
rect 9126 29724 9128 29744
rect 9128 29724 9180 29744
rect 9180 29724 9182 29744
rect 9126 29688 9182 29724
rect 9770 32544 9826 32600
rect 10598 33768 10654 33824
rect 9770 32272 9826 32328
rect 9586 32000 9642 32056
rect 9678 31884 9734 31920
rect 9678 31864 9680 31884
rect 9680 31864 9732 31884
rect 9732 31864 9734 31884
rect 9494 30776 9550 30832
rect 9586 30132 9588 30152
rect 9588 30132 9640 30152
rect 9640 30132 9642 30152
rect 9586 30096 9642 30132
rect 8850 24792 8906 24848
rect 8758 24656 8814 24712
rect 9402 27512 9458 27568
rect 9770 28076 9826 28112
rect 9770 28056 9772 28076
rect 9772 28056 9824 28076
rect 9824 28056 9826 28076
rect 9678 27956 9680 27976
rect 9680 27956 9732 27976
rect 9732 27956 9734 27976
rect 9678 27920 9734 27956
rect 8666 22072 8722 22128
rect 8298 20576 8354 20632
rect 9034 22636 9090 22672
rect 9034 22616 9036 22636
rect 9036 22616 9088 22636
rect 9088 22616 9090 22636
rect 9126 22500 9182 22536
rect 9126 22480 9128 22500
rect 9128 22480 9180 22500
rect 9180 22480 9182 22500
rect 8666 19488 8722 19544
rect 8942 19896 8998 19952
rect 8758 19080 8814 19136
rect 8942 19352 8998 19408
rect 8482 18128 8538 18184
rect 9126 20440 9182 20496
rect 9402 23296 9458 23352
rect 9770 24248 9826 24304
rect 9770 23568 9826 23624
rect 9586 23432 9642 23488
rect 9586 23180 9642 23216
rect 9586 23160 9588 23180
rect 9588 23160 9640 23180
rect 9640 23160 9642 23180
rect 10230 29452 10232 29472
rect 10232 29452 10284 29472
rect 10284 29452 10286 29472
rect 10230 29416 10286 29452
rect 10874 33904 10930 33960
rect 10966 31864 11022 31920
rect 11058 30132 11060 30152
rect 11060 30132 11112 30152
rect 11112 30132 11114 30152
rect 11058 30096 11114 30132
rect 10230 25472 10286 25528
rect 9678 22228 9734 22264
rect 9678 22208 9680 22228
rect 9680 22208 9732 22228
rect 9732 22208 9734 22228
rect 10046 22208 10102 22264
rect 9402 20304 9458 20360
rect 9126 19488 9182 19544
rect 9402 19488 9458 19544
rect 9310 19352 9366 19408
rect 9218 17448 9274 17504
rect 8574 15544 8630 15600
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4986 9580 5042 9616
rect 4986 9560 4988 9580
rect 4988 9560 5040 9580
rect 5040 9560 5042 9580
rect 5814 10684 5816 10704
rect 5816 10684 5868 10704
rect 5868 10684 5870 10704
rect 5814 10648 5870 10684
rect 5446 9580 5502 9616
rect 5446 9560 5448 9580
rect 5448 9560 5500 9580
rect 5500 9560 5502 9580
rect 4894 9152 4950 9208
rect 4894 9036 4950 9072
rect 4894 9016 4896 9036
rect 4896 9016 4948 9036
rect 4948 9016 4950 9036
rect 4710 8880 4766 8936
rect 4434 8336 4490 8392
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4894 8508 4896 8528
rect 4896 8508 4948 8528
rect 4948 8508 4950 8528
rect 4894 8472 4950 8508
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3514 6840 3570 6896
rect 3974 6704 4030 6760
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 5630 9016 5686 9072
rect 4802 7384 4858 7440
rect 6734 12280 6790 12336
rect 6918 12008 6974 12064
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 7194 12724 7196 12744
rect 7196 12724 7248 12744
rect 7248 12724 7250 12744
rect 7194 12688 7250 12724
rect 8758 15272 8814 15328
rect 5998 7284 6000 7304
rect 6000 7284 6052 7304
rect 6052 7284 6054 7304
rect 5998 7248 6054 7284
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 7010 9288 7066 9344
rect 6550 6840 6606 6896
rect 6734 6568 6790 6624
rect 7378 9580 7434 9616
rect 7378 9560 7380 9580
rect 7380 9560 7432 9580
rect 7432 9560 7434 9580
rect 7746 12008 7802 12064
rect 8298 13640 8354 13696
rect 8666 14476 8722 14512
rect 8666 14456 8668 14476
rect 8668 14456 8720 14476
rect 8720 14456 8722 14476
rect 9586 19896 9642 19952
rect 9586 17176 9642 17232
rect 9862 17856 9918 17912
rect 10046 19080 10102 19136
rect 10598 26288 10654 26344
rect 10782 28076 10838 28112
rect 10782 28056 10784 28076
rect 10784 28056 10836 28076
rect 10836 28056 10838 28076
rect 12530 34448 12586 34504
rect 12346 34060 12402 34096
rect 12346 34040 12348 34060
rect 12348 34040 12400 34060
rect 12400 34040 12402 34060
rect 12162 33768 12218 33824
rect 12438 33516 12494 33552
rect 12438 33496 12440 33516
rect 12440 33496 12492 33516
rect 12492 33496 12494 33516
rect 12070 31184 12126 31240
rect 11794 30096 11850 30152
rect 10506 24520 10562 24576
rect 10414 24112 10470 24168
rect 10506 22616 10562 22672
rect 10046 17584 10102 17640
rect 9954 17332 10010 17368
rect 9954 17312 9956 17332
rect 9956 17312 10008 17332
rect 10008 17312 10010 17332
rect 10138 17312 10194 17368
rect 9954 17196 10010 17232
rect 9954 17176 9956 17196
rect 9956 17176 10008 17196
rect 10008 17176 10010 17196
rect 8482 12860 8484 12880
rect 8484 12860 8536 12880
rect 8536 12860 8538 12880
rect 8482 12824 8538 12860
rect 8022 12180 8024 12200
rect 8024 12180 8076 12200
rect 8076 12180 8078 12200
rect 8022 12144 8078 12180
rect 7746 8608 7802 8664
rect 8390 11872 8446 11928
rect 8390 11600 8446 11656
rect 8298 10140 8300 10160
rect 8300 10140 8352 10160
rect 8352 10140 8354 10160
rect 8298 10104 8354 10140
rect 8206 8744 8262 8800
rect 8942 10104 8998 10160
rect 10046 15544 10102 15600
rect 10598 22480 10654 22536
rect 10598 21836 10600 21856
rect 10600 21836 10652 21856
rect 10652 21836 10654 21856
rect 10598 21800 10654 21836
rect 11058 25900 11114 25936
rect 11058 25880 11060 25900
rect 11060 25880 11112 25900
rect 11112 25880 11114 25900
rect 11150 25472 11206 25528
rect 10874 24928 10930 24984
rect 11058 25064 11114 25120
rect 12714 33632 12770 33688
rect 12438 28464 12494 28520
rect 15842 36080 15898 36136
rect 13818 34448 13874 34504
rect 12070 25880 12126 25936
rect 11058 23060 11060 23080
rect 11060 23060 11112 23080
rect 11112 23060 11114 23080
rect 11058 23024 11114 23060
rect 11334 23568 11390 23624
rect 11610 23044 11666 23080
rect 11610 23024 11612 23044
rect 11612 23024 11664 23044
rect 11664 23024 11666 23044
rect 10874 20168 10930 20224
rect 10598 19352 10654 19408
rect 10414 18128 10470 18184
rect 10598 17912 10654 17968
rect 11610 22480 11666 22536
rect 12162 25064 12218 25120
rect 12438 27240 12494 27296
rect 12714 29280 12770 29336
rect 13358 33224 13414 33280
rect 13726 33768 13782 33824
rect 14462 33768 14518 33824
rect 14278 33632 14334 33688
rect 14186 33516 14242 33552
rect 14186 33496 14188 33516
rect 14188 33496 14240 33516
rect 14240 33496 14242 33516
rect 13910 33396 13912 33416
rect 13912 33396 13964 33416
rect 13964 33396 13966 33416
rect 13910 33360 13966 33396
rect 13726 32020 13782 32056
rect 13726 32000 13728 32020
rect 13728 32000 13780 32020
rect 13780 32000 13782 32020
rect 13082 30232 13138 30288
rect 13542 31048 13598 31104
rect 13358 29552 13414 29608
rect 13082 29280 13138 29336
rect 12806 27784 12862 27840
rect 12714 26288 12770 26344
rect 12806 25900 12862 25936
rect 12806 25880 12808 25900
rect 12808 25880 12860 25900
rect 12860 25880 12862 25900
rect 12346 24928 12402 24984
rect 12254 24812 12310 24848
rect 12254 24792 12256 24812
rect 12256 24792 12308 24812
rect 12308 24792 12310 24812
rect 11978 23316 12034 23352
rect 11978 23296 11980 23316
rect 11980 23296 12032 23316
rect 12032 23296 12034 23316
rect 11886 23044 11942 23080
rect 12530 24384 12586 24440
rect 12714 24656 12770 24712
rect 12622 23160 12678 23216
rect 11886 23024 11888 23044
rect 11888 23024 11940 23044
rect 11940 23024 11942 23044
rect 11794 22344 11850 22400
rect 10874 17912 10930 17968
rect 10782 17720 10838 17776
rect 11058 17720 11114 17776
rect 10414 17312 10470 17368
rect 11334 17720 11390 17776
rect 10782 17312 10838 17368
rect 10966 17176 11022 17232
rect 10782 16904 10838 16960
rect 9402 13368 9458 13424
rect 9954 14476 10010 14512
rect 9954 14456 9956 14476
rect 9956 14456 10008 14476
rect 10008 14456 10010 14476
rect 11426 17484 11428 17504
rect 11428 17484 11480 17504
rect 11480 17484 11482 17504
rect 11426 17448 11482 17484
rect 12162 22636 12218 22672
rect 12162 22616 12164 22636
rect 12164 22616 12216 22636
rect 12216 22616 12218 22636
rect 12070 22208 12126 22264
rect 11610 17312 11666 17368
rect 11794 18708 11796 18728
rect 11796 18708 11848 18728
rect 11848 18708 11850 18728
rect 11794 18672 11850 18708
rect 10690 15136 10746 15192
rect 8850 9580 8906 9616
rect 8850 9560 8852 9580
rect 8852 9560 8904 9580
rect 8904 9560 8906 9580
rect 8758 9288 8814 9344
rect 9034 9152 9090 9208
rect 7470 6604 7472 6624
rect 7472 6604 7524 6624
rect 7524 6604 7526 6624
rect 7470 6568 7526 6604
rect 7746 6704 7802 6760
rect 8758 7520 8814 7576
rect 8666 7404 8722 7440
rect 8666 7384 8668 7404
rect 8668 7384 8720 7404
rect 8720 7384 8722 7404
rect 8574 6840 8630 6896
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 9034 7248 9090 7304
rect 9218 6840 9274 6896
rect 9678 8492 9734 8528
rect 9678 8472 9680 8492
rect 9680 8472 9732 8492
rect 9732 8472 9734 8492
rect 10230 13368 10286 13424
rect 10874 12824 10930 12880
rect 10598 11600 10654 11656
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11242 14456 11298 14512
rect 11058 8336 11114 8392
rect 12346 23060 12348 23080
rect 12348 23060 12400 23080
rect 12400 23060 12402 23080
rect 12346 23024 12402 23060
rect 12346 21956 12402 21992
rect 12346 21936 12348 21956
rect 12348 21936 12400 21956
rect 12400 21936 12402 21956
rect 12254 21140 12310 21176
rect 12254 21120 12256 21140
rect 12256 21120 12308 21140
rect 12308 21120 12310 21140
rect 12898 24656 12954 24712
rect 14094 33224 14150 33280
rect 14094 30096 14150 30152
rect 13450 29144 13506 29200
rect 13726 29552 13782 29608
rect 13634 29280 13690 29336
rect 14002 29144 14058 29200
rect 13082 24248 13138 24304
rect 13726 23568 13782 23624
rect 13266 23432 13322 23488
rect 13634 23160 13690 23216
rect 13450 22636 13506 22672
rect 13450 22616 13452 22636
rect 13452 22616 13504 22636
rect 13504 22616 13506 22636
rect 12990 21120 13046 21176
rect 12070 19080 12126 19136
rect 12254 17720 12310 17776
rect 12622 16632 12678 16688
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 11518 6860 11574 6896
rect 11518 6840 11520 6860
rect 11520 6840 11572 6860
rect 11572 6840 11574 6860
rect 11794 7284 11796 7304
rect 11796 7284 11848 7304
rect 11848 7284 11850 7304
rect 11794 7248 11850 7284
rect 12254 7404 12310 7440
rect 12254 7384 12256 7404
rect 12256 7384 12308 7404
rect 12308 7384 12310 7404
rect 12806 16108 12862 16144
rect 12806 16088 12808 16108
rect 12808 16088 12860 16108
rect 12860 16088 12862 16108
rect 12990 18672 13046 18728
rect 13082 17312 13138 17368
rect 15382 35264 15438 35320
rect 14922 34060 14978 34096
rect 14922 34040 14924 34060
rect 14924 34040 14976 34060
rect 14976 34040 14978 34060
rect 15290 33940 15292 33960
rect 15292 33940 15344 33960
rect 15344 33940 15346 33960
rect 15290 33904 15346 33940
rect 15198 33768 15254 33824
rect 14002 23432 14058 23488
rect 14278 26288 14334 26344
rect 14370 22888 14426 22944
rect 15198 33516 15254 33552
rect 15198 33496 15200 33516
rect 15200 33496 15252 33516
rect 15252 33496 15254 33516
rect 15106 31764 15108 31784
rect 15108 31764 15160 31784
rect 15160 31764 15162 31784
rect 15106 31728 15162 31764
rect 16210 34584 16266 34640
rect 15566 33380 15622 33416
rect 15566 33360 15568 33380
rect 15568 33360 15620 33380
rect 15620 33360 15622 33380
rect 15382 31184 15438 31240
rect 14922 29028 14978 29064
rect 14922 29008 14924 29028
rect 14924 29008 14976 29028
rect 14976 29008 14978 29028
rect 14830 26288 14886 26344
rect 14738 26152 14794 26208
rect 14738 23180 14794 23216
rect 14738 23160 14740 23180
rect 14740 23160 14792 23180
rect 14792 23160 14794 23180
rect 14830 22888 14886 22944
rect 14646 22480 14702 22536
rect 14646 20168 14702 20224
rect 14554 19624 14610 19680
rect 13542 17312 13598 17368
rect 13726 17040 13782 17096
rect 12530 9444 12586 9480
rect 12530 9424 12532 9444
rect 12532 9424 12584 9444
rect 12584 9424 12586 9444
rect 11610 6568 11666 6624
rect 11518 6452 11574 6488
rect 11518 6432 11520 6452
rect 11520 6432 11572 6452
rect 11572 6432 11574 6452
rect 11150 3984 11206 4040
rect 12898 5616 12954 5672
rect 15566 31184 15622 31240
rect 15566 30368 15622 30424
rect 15934 31864 15990 31920
rect 16486 34348 16488 34368
rect 16488 34348 16540 34368
rect 16540 34348 16542 34368
rect 16486 34312 16542 34348
rect 16210 30796 16266 30832
rect 16210 30776 16212 30796
rect 16212 30776 16264 30796
rect 16264 30776 16266 30796
rect 16210 30504 16266 30560
rect 15382 29028 15438 29064
rect 15382 29008 15384 29028
rect 15384 29008 15436 29028
rect 15436 29008 15438 29028
rect 15106 24792 15162 24848
rect 15014 21392 15070 21448
rect 15566 28500 15568 28520
rect 15568 28500 15620 28520
rect 15620 28500 15622 28520
rect 15566 28464 15622 28500
rect 15474 28192 15530 28248
rect 15290 23296 15346 23352
rect 15474 23568 15530 23624
rect 15658 23704 15714 23760
rect 15382 22344 15438 22400
rect 15382 22072 15438 22128
rect 15382 21528 15438 21584
rect 14922 18128 14978 18184
rect 15290 17332 15346 17368
rect 15290 17312 15292 17332
rect 15292 17312 15344 17332
rect 15344 17312 15346 17332
rect 15198 15952 15254 16008
rect 15658 22344 15714 22400
rect 15842 22480 15898 22536
rect 15750 21956 15806 21992
rect 15750 21936 15752 21956
rect 15752 21936 15804 21956
rect 15804 21936 15806 21956
rect 17038 34312 17094 34368
rect 16946 34040 17002 34096
rect 17406 36624 17462 36680
rect 18050 34604 18106 34640
rect 18050 34584 18052 34604
rect 18052 34584 18104 34604
rect 18104 34584 18106 34604
rect 18418 36660 18420 36680
rect 18420 36660 18472 36680
rect 18472 36660 18474 36680
rect 18418 36624 18474 36660
rect 19246 36080 19302 36136
rect 18142 33496 18198 33552
rect 16486 30776 16542 30832
rect 16394 30504 16450 30560
rect 18050 33088 18106 33144
rect 19798 36080 19854 36136
rect 18786 34312 18842 34368
rect 20166 34856 20222 34912
rect 22190 36236 22246 36272
rect 22190 36216 22192 36236
rect 22192 36216 22244 36236
rect 22244 36216 22246 36236
rect 18602 32952 18658 33008
rect 16670 29824 16726 29880
rect 16946 29824 17002 29880
rect 16670 28500 16672 28520
rect 16672 28500 16724 28520
rect 16724 28500 16726 28520
rect 16670 28464 16726 28500
rect 16394 27920 16450 27976
rect 16394 26988 16450 27024
rect 16394 26968 16396 26988
rect 16396 26968 16448 26988
rect 16448 26968 16450 26988
rect 16302 24112 16358 24168
rect 16670 26016 16726 26072
rect 16578 24792 16634 24848
rect 16670 24656 16726 24712
rect 16302 23060 16304 23080
rect 16304 23060 16356 23080
rect 16356 23060 16358 23080
rect 16302 23024 16358 23060
rect 16210 20576 16266 20632
rect 16578 22072 16634 22128
rect 17222 29164 17278 29200
rect 17222 29144 17224 29164
rect 17224 29144 17276 29164
rect 17276 29144 17278 29164
rect 16946 26324 16948 26344
rect 16948 26324 17000 26344
rect 17000 26324 17002 26344
rect 16946 26288 17002 26324
rect 16946 24656 17002 24712
rect 16946 24384 17002 24440
rect 17038 23316 17094 23352
rect 17038 23296 17040 23316
rect 17040 23296 17092 23316
rect 17092 23296 17094 23316
rect 16946 23060 16948 23080
rect 16948 23060 17000 23080
rect 17000 23060 17002 23080
rect 16946 23024 17002 23060
rect 17038 22888 17094 22944
rect 16394 21800 16450 21856
rect 16762 21936 16818 21992
rect 15014 13912 15070 13968
rect 15014 13504 15070 13560
rect 14554 11464 14610 11520
rect 14462 10648 14518 10704
rect 13818 9016 13874 9072
rect 13818 7248 13874 7304
rect 13634 6568 13690 6624
rect 13818 6316 13874 6352
rect 13818 6296 13820 6316
rect 13820 6296 13872 6316
rect 13872 6296 13874 6316
rect 13542 5616 13598 5672
rect 14186 7928 14242 7984
rect 15750 19216 15806 19272
rect 15750 16088 15806 16144
rect 16670 20304 16726 20360
rect 17314 26308 17370 26344
rect 17314 26288 17316 26308
rect 17316 26288 17368 26308
rect 17368 26288 17370 26308
rect 17314 26016 17370 26072
rect 17498 26308 17554 26344
rect 17498 26288 17500 26308
rect 17500 26288 17552 26308
rect 17552 26288 17554 26308
rect 17866 30504 17922 30560
rect 18234 29144 18290 29200
rect 17406 23468 17408 23488
rect 17408 23468 17460 23488
rect 17460 23468 17462 23488
rect 17406 23432 17462 23468
rect 17038 20884 17040 20904
rect 17040 20884 17092 20904
rect 17092 20884 17094 20904
rect 17038 20848 17094 20884
rect 16118 17992 16174 18048
rect 15198 6840 15254 6896
rect 16762 20032 16818 20088
rect 17222 20204 17224 20224
rect 17224 20204 17276 20224
rect 17276 20204 17278 20224
rect 17222 20168 17278 20204
rect 18234 28464 18290 28520
rect 18234 26424 18290 26480
rect 17774 23432 17830 23488
rect 17866 23296 17922 23352
rect 17682 22072 17738 22128
rect 17774 21936 17830 21992
rect 17590 20476 17592 20496
rect 17592 20476 17644 20496
rect 17644 20476 17646 20496
rect 17590 20440 17646 20476
rect 16762 19352 16818 19408
rect 16762 18964 16818 19000
rect 16762 18944 16764 18964
rect 16764 18944 16816 18964
rect 16816 18944 16818 18964
rect 16486 11328 16542 11384
rect 17038 19488 17094 19544
rect 16762 12144 16818 12200
rect 16670 11892 16726 11928
rect 16670 11872 16672 11892
rect 16672 11872 16724 11892
rect 16724 11872 16726 11892
rect 16670 11092 16672 11112
rect 16672 11092 16724 11112
rect 16724 11092 16726 11112
rect 16670 11056 16726 11092
rect 16394 8336 16450 8392
rect 16486 7248 16542 7304
rect 17130 16244 17186 16280
rect 17130 16224 17132 16244
rect 17132 16224 17184 16244
rect 17184 16224 17186 16244
rect 17958 20032 18014 20088
rect 17130 12280 17186 12336
rect 18142 23160 18198 23216
rect 18234 22636 18290 22672
rect 18234 22616 18236 22636
rect 18236 22616 18288 22636
rect 18288 22616 18290 22636
rect 20074 32952 20130 33008
rect 20258 32852 20260 32872
rect 20260 32852 20312 32872
rect 20312 32852 20314 32872
rect 18970 29008 19026 29064
rect 18786 28328 18842 28384
rect 18602 26988 18658 27024
rect 18602 26968 18604 26988
rect 18604 26968 18656 26988
rect 18656 26968 18658 26988
rect 18510 26444 18566 26480
rect 18510 26424 18512 26444
rect 18512 26424 18564 26444
rect 18564 26424 18566 26444
rect 18970 27648 19026 27704
rect 19246 28212 19302 28248
rect 19246 28192 19248 28212
rect 19248 28192 19300 28212
rect 19300 28192 19302 28212
rect 19246 24112 19302 24168
rect 19430 28736 19486 28792
rect 19890 32408 19946 32464
rect 19614 30504 19670 30560
rect 19614 29416 19670 29472
rect 19338 23316 19394 23352
rect 19338 23296 19340 23316
rect 19340 23296 19392 23316
rect 19392 23296 19394 23316
rect 19062 23160 19118 23216
rect 18510 22072 18566 22128
rect 18326 20304 18382 20360
rect 18234 19080 18290 19136
rect 18142 18808 18198 18864
rect 17222 11076 17278 11112
rect 17222 11056 17224 11076
rect 17224 11056 17276 11076
rect 17276 11056 17278 11076
rect 15842 4140 15898 4176
rect 15842 4120 15844 4140
rect 15844 4120 15896 4140
rect 15896 4120 15898 4140
rect 17590 12824 17646 12880
rect 18050 17076 18052 17096
rect 18052 17076 18104 17096
rect 18104 17076 18106 17096
rect 18050 17040 18106 17076
rect 17682 12280 17738 12336
rect 18326 12300 18382 12336
rect 18326 12280 18328 12300
rect 18328 12280 18380 12300
rect 18380 12280 18382 12300
rect 17498 11736 17554 11792
rect 17590 11464 17646 11520
rect 17682 11328 17738 11384
rect 17498 11192 17554 11248
rect 17774 10668 17830 10704
rect 17774 10648 17776 10668
rect 17776 10648 17828 10668
rect 17828 10648 17830 10668
rect 17406 10104 17462 10160
rect 17958 10668 18014 10704
rect 17958 10648 17960 10668
rect 17960 10648 18012 10668
rect 18012 10648 18014 10668
rect 17590 9152 17646 9208
rect 17498 5208 17554 5264
rect 16394 3052 16450 3088
rect 16394 3032 16396 3052
rect 16396 3032 16448 3052
rect 16448 3032 16450 3052
rect 18234 8900 18290 8936
rect 18234 8880 18236 8900
rect 18236 8880 18288 8900
rect 18288 8880 18290 8900
rect 17682 6452 17738 6488
rect 17682 6432 17684 6452
rect 17684 6432 17736 6452
rect 17736 6432 17738 6452
rect 18786 23024 18842 23080
rect 18970 23024 19026 23080
rect 19154 22888 19210 22944
rect 19338 21956 19394 21992
rect 19338 21936 19340 21956
rect 19340 21936 19392 21956
rect 19392 21936 19394 21956
rect 19246 21392 19302 21448
rect 19246 20304 19302 20360
rect 19246 19780 19302 19816
rect 19246 19760 19248 19780
rect 19248 19760 19300 19780
rect 19300 19760 19302 19780
rect 18602 18264 18658 18320
rect 18602 12144 18658 12200
rect 18878 13232 18934 13288
rect 18694 10548 18696 10568
rect 18696 10548 18748 10568
rect 18748 10548 18750 10568
rect 18694 10512 18750 10548
rect 18510 9696 18566 9752
rect 18510 6740 18512 6760
rect 18512 6740 18564 6760
rect 18564 6740 18566 6760
rect 18510 6704 18566 6740
rect 19246 15136 19302 15192
rect 19614 23840 19670 23896
rect 20258 32816 20314 32852
rect 19982 27648 20038 27704
rect 20258 26460 20260 26480
rect 20260 26460 20312 26480
rect 20312 26460 20314 26480
rect 20258 26424 20314 26460
rect 19890 23432 19946 23488
rect 19614 22072 19670 22128
rect 19982 23160 20038 23216
rect 19706 18264 19762 18320
rect 21362 35264 21418 35320
rect 23478 36236 23534 36272
rect 23478 36216 23480 36236
rect 23480 36216 23532 36236
rect 23532 36216 23534 36236
rect 22006 33940 22008 33960
rect 22008 33940 22060 33960
rect 22060 33940 22062 33960
rect 22006 33904 22062 33940
rect 21822 32544 21878 32600
rect 22466 32544 22522 32600
rect 22098 32408 22154 32464
rect 22282 32408 22338 32464
rect 23110 33904 23166 33960
rect 21638 32272 21694 32328
rect 20534 25200 20590 25256
rect 20258 21800 20314 21856
rect 19982 19372 20038 19408
rect 19982 19352 19984 19372
rect 19984 19352 20036 19372
rect 20036 19352 20038 19372
rect 19154 13096 19210 13152
rect 19338 14864 19394 14920
rect 19338 13368 19394 13424
rect 19338 13252 19394 13288
rect 19338 13232 19340 13252
rect 19340 13232 19392 13252
rect 19392 13232 19394 13252
rect 19338 12980 19394 13016
rect 19338 12960 19340 12980
rect 19340 12960 19392 12980
rect 19392 12960 19394 12980
rect 19338 12552 19394 12608
rect 18970 9152 19026 9208
rect 19062 8336 19118 8392
rect 19062 7828 19064 7848
rect 19064 7828 19116 7848
rect 19116 7828 19118 7848
rect 19062 7792 19118 7828
rect 19706 13912 19762 13968
rect 20534 24928 20590 24984
rect 21362 30540 21364 30560
rect 21364 30540 21416 30560
rect 21416 30540 21418 30560
rect 21362 30504 21418 30540
rect 20994 29588 20996 29608
rect 20996 29588 21048 29608
rect 21048 29588 21050 29608
rect 20994 29552 21050 29588
rect 21270 29280 21326 29336
rect 20718 26560 20774 26616
rect 21086 28872 21142 28928
rect 21730 29416 21786 29472
rect 21546 29144 21602 29200
rect 21362 28600 21418 28656
rect 21178 26152 21234 26208
rect 20810 24148 20812 24168
rect 20812 24148 20864 24168
rect 20864 24148 20866 24168
rect 20810 24112 20866 24148
rect 19890 13268 19892 13288
rect 19892 13268 19944 13288
rect 19944 13268 19946 13288
rect 19890 13232 19946 13268
rect 19246 8900 19302 8936
rect 19246 8880 19248 8900
rect 19248 8880 19300 8900
rect 19300 8880 19302 8900
rect 18970 7248 19026 7304
rect 18878 6724 18934 6760
rect 18878 6704 18880 6724
rect 18880 6704 18932 6724
rect 18932 6704 18934 6724
rect 19614 10376 19670 10432
rect 20166 13368 20222 13424
rect 20810 20304 20866 20360
rect 21086 20440 21142 20496
rect 21362 25200 21418 25256
rect 22006 30252 22062 30288
rect 22006 30232 22008 30252
rect 22008 30232 22060 30252
rect 22060 30232 22062 30252
rect 22558 31592 22614 31648
rect 21914 28908 21916 28928
rect 21916 28908 21968 28928
rect 21968 28908 21970 28928
rect 21730 28364 21732 28384
rect 21732 28364 21784 28384
rect 21784 28364 21786 28384
rect 21730 28328 21786 28364
rect 21914 28872 21970 28908
rect 22926 32272 22982 32328
rect 23018 31456 23074 31512
rect 22742 29824 22798 29880
rect 21914 26308 21970 26344
rect 21914 26288 21916 26308
rect 21916 26288 21968 26308
rect 21968 26288 21970 26308
rect 21362 20984 21418 21040
rect 21178 17720 21234 17776
rect 20534 14864 20590 14920
rect 20258 11056 20314 11112
rect 20074 10648 20130 10704
rect 19890 10104 19946 10160
rect 20074 9560 20130 9616
rect 19982 6704 20038 6760
rect 18418 4276 18474 4312
rect 18418 4256 18420 4276
rect 18420 4256 18472 4276
rect 18472 4256 18474 4276
rect 18602 4004 18658 4040
rect 18602 3984 18604 4004
rect 18604 3984 18656 4004
rect 18656 3984 18658 4004
rect 20258 8492 20314 8528
rect 20258 8472 20260 8492
rect 20260 8472 20312 8492
rect 20312 8472 20314 8492
rect 21546 18128 21602 18184
rect 22006 25336 22062 25392
rect 22190 26288 22246 26344
rect 22006 22480 22062 22536
rect 22926 28076 22982 28112
rect 22926 28056 22928 28076
rect 22928 28056 22980 28076
rect 22980 28056 22982 28076
rect 22834 27784 22890 27840
rect 23846 32816 23902 32872
rect 23662 32544 23718 32600
rect 23754 31728 23810 31784
rect 23478 30912 23534 30968
rect 23294 29164 23350 29200
rect 23294 29144 23296 29164
rect 23296 29144 23348 29164
rect 23348 29144 23350 29164
rect 23570 30232 23626 30288
rect 25594 36100 25650 36136
rect 25594 36080 25596 36100
rect 25596 36080 25648 36100
rect 25648 36080 25650 36100
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 24030 32852 24032 32872
rect 24032 32852 24084 32872
rect 24084 32852 24086 32872
rect 24030 32816 24086 32852
rect 24306 32428 24362 32464
rect 24306 32408 24308 32428
rect 24308 32408 24360 32428
rect 24360 32408 24362 32428
rect 24030 31592 24086 31648
rect 23754 30096 23810 30152
rect 23110 27820 23112 27840
rect 23112 27820 23164 27840
rect 23164 27820 23166 27840
rect 23110 27784 23166 27820
rect 22650 23704 22706 23760
rect 20810 15036 20812 15056
rect 20812 15036 20864 15056
rect 20864 15036 20866 15056
rect 20810 15000 20866 15036
rect 20718 14356 20720 14376
rect 20720 14356 20772 14376
rect 20772 14356 20774 14376
rect 20718 14320 20774 14356
rect 21638 17584 21694 17640
rect 21914 17992 21970 18048
rect 21638 16124 21640 16144
rect 21640 16124 21692 16144
rect 21692 16124 21694 16144
rect 21638 16088 21694 16124
rect 21362 15000 21418 15056
rect 21270 14864 21326 14920
rect 21914 16768 21970 16824
rect 22558 19624 22614 19680
rect 22650 19488 22706 19544
rect 22558 19352 22614 19408
rect 22190 15988 22192 16008
rect 22192 15988 22244 16008
rect 22244 15988 22246 16008
rect 22190 15952 22246 15988
rect 22098 15272 22154 15328
rect 22006 14864 22062 14920
rect 21178 12552 21234 12608
rect 21546 13504 21602 13560
rect 21270 12144 21326 12200
rect 20902 10648 20958 10704
rect 21454 11736 21510 11792
rect 21362 10648 21418 10704
rect 20810 9424 20866 9480
rect 21086 7928 21142 7984
rect 21178 7828 21180 7848
rect 21180 7828 21232 7848
rect 21232 7828 21234 7848
rect 21178 7792 21234 7828
rect 21546 10512 21602 10568
rect 22466 17312 22522 17368
rect 22558 17176 22614 17232
rect 22650 16360 22706 16416
rect 23018 22108 23020 22128
rect 23020 22108 23072 22128
rect 23072 22108 23074 22128
rect 23018 22072 23074 22108
rect 23294 26460 23296 26480
rect 23296 26460 23348 26480
rect 23348 26460 23350 26480
rect 23294 26424 23350 26460
rect 22834 19388 22836 19408
rect 22836 19388 22888 19408
rect 22888 19388 22890 19408
rect 22834 19352 22890 19388
rect 22834 17620 22836 17640
rect 22836 17620 22888 17640
rect 22888 17620 22890 17640
rect 22834 17584 22890 17620
rect 21638 10104 21694 10160
rect 21362 8472 21418 8528
rect 21638 7112 21694 7168
rect 21546 6840 21602 6896
rect 21546 5344 21602 5400
rect 21086 5092 21142 5128
rect 21086 5072 21088 5092
rect 21088 5072 21140 5092
rect 21140 5072 21142 5092
rect 20994 4140 21050 4176
rect 20994 4120 20996 4140
rect 20996 4120 21048 4140
rect 21048 4120 21050 4140
rect 21086 3612 21088 3632
rect 21088 3612 21140 3632
rect 21140 3612 21142 3632
rect 21086 3576 21142 3612
rect 22282 12416 22338 12472
rect 22282 9444 22338 9480
rect 22282 9424 22284 9444
rect 22284 9424 22336 9444
rect 22336 9424 22338 9444
rect 23938 25744 23994 25800
rect 24674 32408 24730 32464
rect 24490 31456 24546 31512
rect 23294 20304 23350 20360
rect 23662 20304 23718 20360
rect 23294 19624 23350 19680
rect 23202 19508 23258 19544
rect 23202 19488 23204 19508
rect 23204 19488 23256 19508
rect 23256 19488 23258 19508
rect 23202 19352 23258 19408
rect 23110 18128 23166 18184
rect 23018 17312 23074 17368
rect 23294 19252 23296 19272
rect 23296 19252 23348 19272
rect 23348 19252 23350 19272
rect 23294 19216 23350 19252
rect 23294 18808 23350 18864
rect 24950 31592 25006 31648
rect 24858 30540 24860 30560
rect 24860 30540 24912 30560
rect 24912 30540 24914 30560
rect 24858 30504 24914 30540
rect 25594 32272 25650 32328
rect 25318 31592 25374 31648
rect 25226 29416 25282 29472
rect 24950 28500 24952 28520
rect 24952 28500 25004 28520
rect 25004 28500 25006 28520
rect 24490 26832 24546 26888
rect 24398 24792 24454 24848
rect 23018 15952 23074 16008
rect 23202 15444 23204 15464
rect 23204 15444 23256 15464
rect 23256 15444 23258 15464
rect 23202 15408 23258 15444
rect 23202 12416 23258 12472
rect 23938 18400 23994 18456
rect 23938 17992 23994 18048
rect 24398 22344 24454 22400
rect 24950 28464 25006 28500
rect 25134 28464 25190 28520
rect 25410 28192 25466 28248
rect 24858 27648 24914 27704
rect 24122 19372 24178 19408
rect 24122 19352 24124 19372
rect 24124 19352 24176 19372
rect 24176 19352 24178 19372
rect 23478 15988 23480 16008
rect 23480 15988 23532 16008
rect 23532 15988 23534 16008
rect 23478 15952 23534 15988
rect 23570 12588 23572 12608
rect 23572 12588 23624 12608
rect 23624 12588 23626 12608
rect 23570 12552 23626 12588
rect 22926 10684 22928 10704
rect 22928 10684 22980 10704
rect 22980 10684 22982 10704
rect 22926 10648 22982 10684
rect 23110 10240 23166 10296
rect 23478 10104 23534 10160
rect 23386 9288 23442 9344
rect 23570 8472 23626 8528
rect 22006 5364 22062 5400
rect 22006 5344 22008 5364
rect 22008 5344 22060 5364
rect 22060 5344 22062 5364
rect 20442 3168 20498 3224
rect 22190 4020 22192 4040
rect 22192 4020 22244 4040
rect 22244 4020 22246 4040
rect 22190 3984 22246 4020
rect 21914 3168 21970 3224
rect 22834 6840 22890 6896
rect 23846 12144 23902 12200
rect 23938 12008 23994 12064
rect 24030 11872 24086 11928
rect 24030 9424 24086 9480
rect 24674 18264 24730 18320
rect 24582 18128 24638 18184
rect 24214 14900 24216 14920
rect 24216 14900 24268 14920
rect 24268 14900 24270 14920
rect 24214 14864 24270 14900
rect 24214 13932 24270 13968
rect 24214 13912 24216 13932
rect 24216 13912 24268 13932
rect 24268 13912 24270 13932
rect 25410 25336 25466 25392
rect 25410 23432 25466 23488
rect 25410 22616 25466 22672
rect 25318 20984 25374 21040
rect 25134 18808 25190 18864
rect 24858 13912 24914 13968
rect 25686 31456 25742 31512
rect 25594 29280 25650 29336
rect 25778 28736 25834 28792
rect 25870 27940 25926 27976
rect 25870 27920 25872 27940
rect 25872 27920 25924 27940
rect 25924 27920 25926 27940
rect 25870 27512 25926 27568
rect 26422 32680 26478 32736
rect 26698 32408 26754 32464
rect 26422 32000 26478 32056
rect 26698 31728 26754 31784
rect 26238 31592 26294 31648
rect 26238 31048 26294 31104
rect 26606 31048 26662 31104
rect 26238 30368 26294 30424
rect 26238 29552 26294 29608
rect 26054 27376 26110 27432
rect 25594 26460 25596 26480
rect 25596 26460 25648 26480
rect 25648 26460 25650 26480
rect 25594 26424 25650 26460
rect 25778 26444 25834 26480
rect 25778 26424 25780 26444
rect 25780 26424 25832 26444
rect 25832 26424 25834 26444
rect 25870 24812 25926 24848
rect 26606 30776 26662 30832
rect 26606 30368 26662 30424
rect 26606 30252 26662 30288
rect 26606 30232 26608 30252
rect 26608 30232 26660 30252
rect 26660 30232 26662 30252
rect 27250 32816 27306 32872
rect 27066 31764 27068 31784
rect 27068 31764 27120 31784
rect 27120 31764 27122 31784
rect 27066 31728 27122 31764
rect 26974 31592 27030 31648
rect 27250 31456 27306 31512
rect 27894 32952 27950 33008
rect 28906 32952 28962 33008
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 28354 32680 28410 32736
rect 28630 32680 28686 32736
rect 28170 32544 28226 32600
rect 28170 32444 28172 32464
rect 28172 32444 28224 32464
rect 28224 32444 28226 32464
rect 28170 32408 28226 32444
rect 27618 31764 27620 31784
rect 27620 31764 27672 31784
rect 27672 31764 27674 31784
rect 27618 31728 27674 31764
rect 27434 31592 27490 31648
rect 27342 30776 27398 30832
rect 27250 30232 27306 30288
rect 27618 30776 27674 30832
rect 27434 30504 27490 30560
rect 26422 27240 26478 27296
rect 26238 26424 26294 26480
rect 25870 24792 25872 24812
rect 25872 24792 25924 24812
rect 25924 24792 25926 24812
rect 25594 22344 25650 22400
rect 26974 28872 27030 28928
rect 26882 28192 26938 28248
rect 27342 29416 27398 29472
rect 26974 27940 27030 27976
rect 26974 27920 26976 27940
rect 26976 27920 27028 27940
rect 27028 27920 27030 27940
rect 26974 27512 27030 27568
rect 26882 27104 26938 27160
rect 26238 21972 26240 21992
rect 26240 21972 26292 21992
rect 26292 21972 26294 21992
rect 26238 21936 26294 21972
rect 26146 20712 26202 20768
rect 25594 19216 25650 19272
rect 25594 18692 25650 18728
rect 25594 18672 25596 18692
rect 25596 18672 25648 18692
rect 25648 18672 25650 18692
rect 25410 18284 25466 18320
rect 25410 18264 25412 18284
rect 25412 18264 25464 18284
rect 25464 18264 25466 18284
rect 24490 10260 24546 10296
rect 24490 10240 24492 10260
rect 24492 10240 24544 10260
rect 24544 10240 24546 10260
rect 24306 9424 24362 9480
rect 24398 9152 24454 9208
rect 24306 8880 24362 8936
rect 25042 10376 25098 10432
rect 25962 19796 25964 19816
rect 25964 19796 26016 19816
rect 26016 19796 26018 19816
rect 25962 19760 26018 19796
rect 25502 17720 25558 17776
rect 25594 14900 25596 14920
rect 25596 14900 25648 14920
rect 25648 14900 25650 14920
rect 25594 14864 25650 14900
rect 26146 18128 26202 18184
rect 26514 20576 26570 20632
rect 25778 14320 25834 14376
rect 25318 10648 25374 10704
rect 25686 11056 25742 11112
rect 26054 12416 26110 12472
rect 25594 10376 25650 10432
rect 25410 9696 25466 9752
rect 26238 10104 26294 10160
rect 27250 28736 27306 28792
rect 27618 30676 27620 30696
rect 27620 30676 27672 30696
rect 27672 30676 27674 30696
rect 27618 30640 27674 30676
rect 27710 30232 27766 30288
rect 28262 32272 28318 32328
rect 28078 31320 28134 31376
rect 28078 31048 28134 31104
rect 27986 30640 28042 30696
rect 27802 29824 27858 29880
rect 27710 29688 27766 29744
rect 27710 29416 27766 29472
rect 27342 27648 27398 27704
rect 27250 27240 27306 27296
rect 27158 27104 27214 27160
rect 27158 26832 27214 26888
rect 27618 27376 27674 27432
rect 28262 31592 28318 31648
rect 28262 31320 28318 31376
rect 28262 30268 28264 30288
rect 28264 30268 28316 30288
rect 28316 30268 28318 30288
rect 28262 30232 28318 30268
rect 28078 29960 28134 30016
rect 28078 29824 28134 29880
rect 27986 29552 28042 29608
rect 28262 29588 28264 29608
rect 28264 29588 28316 29608
rect 28316 29588 28318 29608
rect 28262 29552 28318 29588
rect 28262 29164 28318 29200
rect 28262 29144 28264 29164
rect 28264 29144 28316 29164
rect 28316 29144 28318 29164
rect 26606 19080 26662 19136
rect 26698 18808 26754 18864
rect 26514 16632 26570 16688
rect 26698 11892 26754 11928
rect 26698 11872 26700 11892
rect 26700 11872 26752 11892
rect 26752 11872 26754 11892
rect 26238 9560 26294 9616
rect 26054 9424 26110 9480
rect 26146 9152 26202 9208
rect 25502 8200 25558 8256
rect 24950 7268 25006 7304
rect 24950 7248 24952 7268
rect 24952 7248 25004 7268
rect 25004 7248 25006 7268
rect 23846 4548 23902 4584
rect 23846 4528 23848 4548
rect 23848 4528 23900 4548
rect 23900 4528 23902 4548
rect 23570 4140 23626 4176
rect 23570 4120 23572 4140
rect 23572 4120 23624 4140
rect 23624 4120 23626 4140
rect 23938 3984 23994 4040
rect 26054 7928 26110 7984
rect 27158 24676 27214 24712
rect 27158 24656 27160 24676
rect 27160 24656 27212 24676
rect 27212 24656 27214 24676
rect 27066 20460 27122 20496
rect 27066 20440 27068 20460
rect 27068 20440 27120 20460
rect 27120 20440 27122 20460
rect 27526 24148 27528 24168
rect 27528 24148 27580 24168
rect 27580 24148 27582 24168
rect 27526 24112 27582 24148
rect 28262 28756 28318 28792
rect 28262 28736 28264 28756
rect 28264 28736 28316 28756
rect 28316 28736 28318 28756
rect 28262 28500 28264 28520
rect 28264 28500 28316 28520
rect 28316 28500 28318 28520
rect 28262 28464 28318 28500
rect 28262 27104 28318 27160
rect 28814 31628 28816 31648
rect 28816 31628 28868 31648
rect 28868 31628 28870 31648
rect 28814 31592 28870 31628
rect 28538 30912 28594 30968
rect 28722 30776 28778 30832
rect 28446 29688 28502 29744
rect 28446 28872 28502 28928
rect 28446 28736 28502 28792
rect 28906 30252 28962 30288
rect 28906 30232 28908 30252
rect 28908 30232 28960 30252
rect 28960 30232 28962 30252
rect 29182 31728 29238 31784
rect 29182 30132 29184 30152
rect 29184 30132 29236 30152
rect 29236 30132 29238 30152
rect 29182 30096 29238 30132
rect 27986 20712 28042 20768
rect 27434 18264 27490 18320
rect 26974 16768 27030 16824
rect 27250 14864 27306 14920
rect 26790 9560 26846 9616
rect 26790 9288 26846 9344
rect 26698 8744 26754 8800
rect 26698 8492 26754 8528
rect 26698 8472 26700 8492
rect 26700 8472 26752 8492
rect 26752 8472 26754 8492
rect 27250 13776 27306 13832
rect 27618 17040 27674 17096
rect 27618 15272 27674 15328
rect 27250 11756 27306 11792
rect 27250 11736 27252 11756
rect 27252 11736 27304 11756
rect 27304 11736 27306 11756
rect 26882 9016 26938 9072
rect 27066 8916 27068 8936
rect 27068 8916 27120 8936
rect 27120 8916 27122 8936
rect 27066 8880 27122 8916
rect 26974 8200 27030 8256
rect 26790 7928 26846 7984
rect 26054 5616 26110 5672
rect 22282 3168 22338 3224
rect 27710 14456 27766 14512
rect 27618 14184 27674 14240
rect 27894 16108 27950 16144
rect 28170 22480 28226 22536
rect 28814 27920 28870 27976
rect 28630 27512 28686 27568
rect 28262 20440 28318 20496
rect 27894 16088 27896 16108
rect 27896 16088 27948 16108
rect 27948 16088 27950 16108
rect 27710 11872 27766 11928
rect 27342 9016 27398 9072
rect 27802 7948 27858 7984
rect 27802 7928 27804 7948
rect 27804 7928 27856 7948
rect 27856 7928 27858 7948
rect 28814 24792 28870 24848
rect 28722 24656 28778 24712
rect 28722 24384 28778 24440
rect 28814 23432 28870 23488
rect 29366 30252 29422 30288
rect 29366 30232 29368 30252
rect 29368 30232 29420 30252
rect 29420 30232 29422 30252
rect 29550 31728 29606 31784
rect 29918 32000 29974 32056
rect 29366 25644 29368 25664
rect 29368 25644 29420 25664
rect 29420 25644 29422 25664
rect 29366 25608 29422 25644
rect 28998 22208 29054 22264
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 31114 32716 31116 32736
rect 31116 32716 31168 32736
rect 31168 32716 31170 32736
rect 30194 32544 30250 32600
rect 31114 32680 31170 32716
rect 30378 32136 30434 32192
rect 30654 32308 30656 32328
rect 30656 32308 30708 32328
rect 30708 32308 30710 32328
rect 30654 32272 30710 32308
rect 30470 32000 30526 32056
rect 30194 31456 30250 31512
rect 30470 31628 30472 31648
rect 30472 31628 30524 31648
rect 30524 31628 30526 31648
rect 30470 31592 30526 31628
rect 30838 32000 30894 32056
rect 31022 32272 31078 32328
rect 30286 31204 30342 31240
rect 30286 31184 30288 31204
rect 30288 31184 30340 31204
rect 30340 31184 30342 31204
rect 30838 30504 30894 30560
rect 30010 29028 30066 29064
rect 30010 29008 30012 29028
rect 30012 29008 30064 29028
rect 30064 29008 30066 29028
rect 30010 28328 30066 28384
rect 29918 28076 29974 28112
rect 29918 28056 29920 28076
rect 29920 28056 29972 28076
rect 29972 28056 29974 28076
rect 30102 27532 30158 27568
rect 30102 27512 30104 27532
rect 30104 27512 30156 27532
rect 30156 27512 30158 27532
rect 30010 24928 30066 24984
rect 30194 25644 30196 25664
rect 30196 25644 30248 25664
rect 30248 25644 30250 25664
rect 30194 25608 30250 25644
rect 30378 29416 30434 29472
rect 30654 29960 30710 30016
rect 30746 29572 30802 29608
rect 30746 29552 30748 29572
rect 30748 29552 30800 29572
rect 30800 29552 30802 29572
rect 30378 27512 30434 27568
rect 31114 30252 31170 30288
rect 31114 30232 31116 30252
rect 31116 30232 31168 30252
rect 31168 30232 31170 30252
rect 31022 29960 31078 30016
rect 31022 27920 31078 27976
rect 31298 32680 31354 32736
rect 31850 32544 31906 32600
rect 31574 32428 31630 32464
rect 31574 32408 31576 32428
rect 31576 32408 31628 32428
rect 31628 32408 31630 32428
rect 32218 32680 32274 32736
rect 32402 32272 32458 32328
rect 31942 32136 31998 32192
rect 32218 32000 32274 32056
rect 31022 27512 31078 27568
rect 30930 24284 30932 24304
rect 30932 24284 30984 24304
rect 30984 24284 30986 24304
rect 30930 24248 30986 24284
rect 30930 23432 30986 23488
rect 30378 19352 30434 19408
rect 29274 12416 29330 12472
rect 28998 11600 29054 11656
rect 28262 9560 28318 9616
rect 28170 7112 28226 7168
rect 27802 6704 27858 6760
rect 27526 6296 27582 6352
rect 29090 10532 29146 10568
rect 29090 10512 29092 10532
rect 29092 10512 29144 10532
rect 29144 10512 29146 10532
rect 30654 17332 30710 17368
rect 30654 17312 30656 17332
rect 30656 17312 30708 17332
rect 30708 17312 30710 17332
rect 28722 8880 28778 8936
rect 28538 7948 28594 7984
rect 28538 7928 28540 7948
rect 28540 7928 28592 7948
rect 28592 7928 28594 7948
rect 28538 7384 28594 7440
rect 29182 9832 29238 9888
rect 28998 9696 29054 9752
rect 29826 9696 29882 9752
rect 29274 8492 29330 8528
rect 29274 8472 29276 8492
rect 29276 8472 29328 8492
rect 29328 8472 29330 8492
rect 30102 11756 30158 11792
rect 30654 13776 30710 13832
rect 30562 12280 30618 12336
rect 30654 12008 30710 12064
rect 30102 11736 30104 11756
rect 30104 11736 30156 11756
rect 30156 11736 30158 11756
rect 30286 11600 30342 11656
rect 30194 10240 30250 10296
rect 31482 29164 31538 29200
rect 31482 29144 31484 29164
rect 31484 29144 31536 29164
rect 31536 29144 31538 29164
rect 31390 27784 31446 27840
rect 31666 29416 31722 29472
rect 31666 26832 31722 26888
rect 31298 24928 31354 24984
rect 32034 25472 32090 25528
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 32586 32272 32642 32328
rect 32586 32020 32642 32056
rect 32586 32000 32588 32020
rect 32588 32000 32640 32020
rect 32640 32000 32642 32020
rect 34426 32408 34482 32464
rect 32310 25880 32366 25936
rect 32218 25336 32274 25392
rect 31482 24248 31538 24304
rect 31298 23704 31354 23760
rect 31298 22072 31354 22128
rect 32218 25064 32274 25120
rect 31298 19352 31354 19408
rect 32770 25472 32826 25528
rect 34058 30368 34114 30424
rect 33414 29008 33470 29064
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 30930 11872 30986 11928
rect 30838 11192 30894 11248
rect 31022 11464 31078 11520
rect 31574 15564 31630 15600
rect 31574 15544 31576 15564
rect 31576 15544 31628 15564
rect 31628 15544 31630 15564
rect 31574 12960 31630 13016
rect 32126 15156 32182 15192
rect 32126 15136 32128 15156
rect 32128 15136 32180 15156
rect 32180 15136 32182 15156
rect 31574 11872 31630 11928
rect 31390 11464 31446 11520
rect 31298 10512 31354 10568
rect 31206 10260 31262 10296
rect 31206 10240 31208 10260
rect 31208 10240 31260 10260
rect 31260 10240 31262 10260
rect 31390 10376 31446 10432
rect 30838 9288 30894 9344
rect 30930 8508 30932 8528
rect 30932 8508 30984 8528
rect 30984 8508 30986 8528
rect 30930 8472 30986 8508
rect 30838 8336 30894 8392
rect 31390 9424 31446 9480
rect 31666 11328 31722 11384
rect 31850 11192 31906 11248
rect 32034 11600 32090 11656
rect 32034 10920 32090 10976
rect 31666 9424 31722 9480
rect 32494 13388 32550 13424
rect 32494 13368 32496 13388
rect 32496 13368 32548 13388
rect 32548 13368 32550 13388
rect 32402 11464 32458 11520
rect 32402 10920 32458 10976
rect 32954 18128 33010 18184
rect 32678 12144 32734 12200
rect 32954 11872 33010 11928
rect 32494 9988 32550 10024
rect 32494 9968 32496 9988
rect 32496 9968 32548 9988
rect 32548 9968 32550 9988
rect 31942 5908 31998 5944
rect 31942 5888 31944 5908
rect 31944 5888 31996 5908
rect 31996 5888 31998 5908
rect 32494 9424 32550 9480
rect 32310 8336 32366 8392
rect 33966 24928 34022 24984
rect 33690 13776 33746 13832
rect 33138 9696 33194 9752
rect 32954 8608 33010 8664
rect 33046 7520 33102 7576
rect 35806 29008 35862 29064
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35990 24520 36046 24576
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34518 20712 34574 20768
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35254 21392 35310 21448
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35254 19216 35310 19272
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 36082 23840 36138 23896
rect 36082 22480 36138 22536
rect 36082 21800 36138 21856
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 35806 21392 35862 21448
rect 36082 21120 36138 21176
rect 35806 20848 35862 20904
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35254 16496 35310 16552
rect 34794 16088 34850 16144
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 33506 9580 33562 9616
rect 33506 9560 33508 9580
rect 33508 9560 33560 9580
rect 33560 9560 33562 9580
rect 34426 10260 34482 10296
rect 34426 10240 34428 10260
rect 34428 10240 34480 10260
rect 34480 10240 34482 10260
rect 34242 9696 34298 9752
rect 34058 9560 34114 9616
rect 30378 5092 30434 5128
rect 30378 5072 30380 5092
rect 30380 5072 30432 5092
rect 30432 5072 30434 5092
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 35530 16088 35586 16144
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 35070 14456 35126 14512
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34794 12280 34850 12336
rect 34978 12164 35034 12200
rect 34978 12144 34980 12164
rect 34980 12144 35032 12164
rect 35032 12144 35034 12164
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 36082 12144 36138 12200
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 35346 9832 35402 9888
rect 35162 9596 35164 9616
rect 35164 9596 35216 9616
rect 35216 9596 35218 9616
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 35162 9560 35218 9596
rect 34978 9424 35034 9480
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35530 9424 35586 9480
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 36450 27920 36506 27976
rect 36082 3476 36084 3496
rect 36084 3476 36136 3496
rect 36136 3476 36138 3496
rect 36082 3440 36138 3476
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 17401 36682 17467 36685
rect 18413 36682 18479 36685
rect 17401 36680 18479 36682
rect 17401 36624 17406 36680
rect 17462 36624 18418 36680
rect 18474 36624 18479 36680
rect 17401 36622 18479 36624
rect 17401 36619 17467 36622
rect 18413 36619 18479 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 22185 36274 22251 36277
rect 23473 36274 23539 36277
rect 22185 36272 23539 36274
rect 22185 36216 22190 36272
rect 22246 36216 23478 36272
rect 23534 36216 23539 36272
rect 22185 36214 23539 36216
rect 22185 36211 22251 36214
rect 23473 36211 23539 36214
rect 15837 36138 15903 36141
rect 19241 36138 19307 36141
rect 15837 36136 19307 36138
rect 15837 36080 15842 36136
rect 15898 36080 19246 36136
rect 19302 36080 19307 36136
rect 15837 36078 19307 36080
rect 15837 36075 15903 36078
rect 19241 36075 19307 36078
rect 19793 36138 19859 36141
rect 25589 36138 25655 36141
rect 19793 36136 25655 36138
rect 19793 36080 19798 36136
rect 19854 36080 25594 36136
rect 25650 36080 25655 36136
rect 19793 36078 25655 36080
rect 19793 36075 19859 36078
rect 25589 36075 25655 36078
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 0 35458 800 35488
rect 3693 35458 3759 35461
rect 0 35456 3759 35458
rect 0 35400 3698 35456
rect 3754 35400 3759 35456
rect 0 35398 3759 35400
rect 0 35368 800 35398
rect 3693 35395 3759 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 15377 35322 15443 35325
rect 21357 35322 21423 35325
rect 15377 35320 21423 35322
rect 15377 35264 15382 35320
rect 15438 35264 21362 35320
rect 21418 35264 21423 35320
rect 15377 35262 21423 35264
rect 15377 35259 15443 35262
rect 21357 35259 21423 35262
rect 20161 34914 20227 34917
rect 20294 34914 20300 34916
rect 20161 34912 20300 34914
rect 20161 34856 20166 34912
rect 20222 34856 20300 34912
rect 20161 34854 20300 34856
rect 20161 34851 20227 34854
rect 20294 34852 20300 34854
rect 20364 34852 20370 34916
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 16205 34642 16271 34645
rect 18045 34642 18111 34645
rect 16205 34640 18111 34642
rect 16205 34584 16210 34640
rect 16266 34584 18050 34640
rect 18106 34584 18111 34640
rect 16205 34582 18111 34584
rect 16205 34579 16271 34582
rect 18045 34579 18111 34582
rect 12525 34506 12591 34509
rect 13813 34506 13879 34509
rect 12525 34504 13879 34506
rect 12525 34448 12530 34504
rect 12586 34448 13818 34504
rect 13874 34448 13879 34504
rect 12525 34446 13879 34448
rect 12525 34443 12591 34446
rect 13813 34443 13879 34446
rect 16481 34370 16547 34373
rect 17033 34370 17099 34373
rect 18781 34370 18847 34373
rect 16481 34368 18847 34370
rect 16481 34312 16486 34368
rect 16542 34312 17038 34368
rect 17094 34312 18786 34368
rect 18842 34312 18847 34368
rect 16481 34310 18847 34312
rect 16481 34307 16547 34310
rect 17033 34307 17099 34310
rect 18781 34307 18847 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 12341 34098 12407 34101
rect 14917 34098 14983 34101
rect 16941 34098 17007 34101
rect 12341 34096 17007 34098
rect 12341 34040 12346 34096
rect 12402 34040 14922 34096
rect 14978 34040 16946 34096
rect 17002 34040 17007 34096
rect 12341 34038 17007 34040
rect 12341 34035 12407 34038
rect 14917 34035 14983 34038
rect 16941 34035 17007 34038
rect 10869 33962 10935 33965
rect 15285 33962 15351 33965
rect 10869 33960 15351 33962
rect 10869 33904 10874 33960
rect 10930 33904 15290 33960
rect 15346 33904 15351 33960
rect 10869 33902 15351 33904
rect 10869 33899 10935 33902
rect 15285 33899 15351 33902
rect 22001 33962 22067 33965
rect 23105 33962 23171 33965
rect 22001 33960 23171 33962
rect 22001 33904 22006 33960
rect 22062 33904 23110 33960
rect 23166 33904 23171 33960
rect 22001 33902 23171 33904
rect 22001 33899 22067 33902
rect 23105 33899 23171 33902
rect 6545 33826 6611 33829
rect 10593 33826 10659 33829
rect 6545 33824 10659 33826
rect 6545 33768 6550 33824
rect 6606 33768 10598 33824
rect 10654 33768 10659 33824
rect 6545 33766 10659 33768
rect 6545 33763 6611 33766
rect 10593 33763 10659 33766
rect 12157 33826 12223 33829
rect 13721 33826 13787 33829
rect 14457 33826 14523 33829
rect 15193 33826 15259 33829
rect 12157 33824 15259 33826
rect 12157 33768 12162 33824
rect 12218 33768 13726 33824
rect 13782 33768 14462 33824
rect 14518 33768 15198 33824
rect 15254 33768 15259 33824
rect 12157 33766 15259 33768
rect 12157 33763 12223 33766
rect 13721 33763 13787 33766
rect 14457 33763 14523 33766
rect 15193 33763 15259 33766
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 12709 33690 12775 33693
rect 14273 33690 14339 33693
rect 12709 33688 14339 33690
rect 12709 33632 12714 33688
rect 12770 33632 14278 33688
rect 14334 33632 14339 33688
rect 12709 33630 14339 33632
rect 12709 33627 12775 33630
rect 14273 33627 14339 33630
rect 12433 33554 12499 33557
rect 14181 33554 14247 33557
rect 12433 33552 14247 33554
rect 12433 33496 12438 33552
rect 12494 33496 14186 33552
rect 14242 33496 14247 33552
rect 12433 33494 14247 33496
rect 12433 33491 12499 33494
rect 14181 33491 14247 33494
rect 15193 33554 15259 33557
rect 18137 33554 18203 33557
rect 15193 33552 18203 33554
rect 15193 33496 15198 33552
rect 15254 33496 18142 33552
rect 18198 33496 18203 33552
rect 15193 33494 18203 33496
rect 15193 33491 15259 33494
rect 18137 33491 18203 33494
rect 8845 33418 8911 33421
rect 9397 33418 9463 33421
rect 8845 33416 9463 33418
rect 8845 33360 8850 33416
rect 8906 33360 9402 33416
rect 9458 33360 9463 33416
rect 8845 33358 9463 33360
rect 8845 33355 8911 33358
rect 9397 33355 9463 33358
rect 13905 33418 13971 33421
rect 15561 33418 15627 33421
rect 13905 33416 15627 33418
rect 13905 33360 13910 33416
rect 13966 33360 15566 33416
rect 15622 33360 15627 33416
rect 13905 33358 15627 33360
rect 13905 33355 13971 33358
rect 15561 33355 15627 33358
rect 13353 33282 13419 33285
rect 14089 33282 14155 33285
rect 13353 33280 14155 33282
rect 13353 33224 13358 33280
rect 13414 33224 14094 33280
rect 14150 33224 14155 33280
rect 13353 33222 14155 33224
rect 13353 33219 13419 33222
rect 14089 33219 14155 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 9622 33084 9628 33148
rect 9692 33146 9698 33148
rect 18045 33146 18111 33149
rect 9692 33144 18111 33146
rect 9692 33088 18050 33144
rect 18106 33088 18111 33144
rect 9692 33086 18111 33088
rect 9692 33084 9698 33086
rect 18045 33083 18111 33086
rect 4654 32948 4660 33012
rect 4724 33010 4730 33012
rect 4797 33010 4863 33013
rect 4724 33008 4863 33010
rect 4724 32952 4802 33008
rect 4858 32952 4863 33008
rect 4724 32950 4863 32952
rect 4724 32948 4730 32950
rect 4797 32947 4863 32950
rect 5165 33010 5231 33013
rect 6453 33010 6519 33013
rect 7373 33010 7439 33013
rect 5165 33008 7439 33010
rect 5165 32952 5170 33008
rect 5226 32952 6458 33008
rect 6514 32952 7378 33008
rect 7434 32952 7439 33008
rect 5165 32950 7439 32952
rect 5165 32947 5231 32950
rect 6453 32947 6519 32950
rect 7373 32947 7439 32950
rect 10910 32948 10916 33012
rect 10980 33010 10986 33012
rect 18597 33010 18663 33013
rect 10980 33008 18663 33010
rect 10980 32952 18602 33008
rect 18658 32952 18663 33008
rect 10980 32950 18663 32952
rect 10980 32948 10986 32950
rect 18597 32947 18663 32950
rect 20069 33010 20135 33013
rect 27889 33010 27955 33013
rect 28901 33010 28967 33013
rect 20069 33008 28967 33010
rect 20069 32952 20074 33008
rect 20130 32952 27894 33008
rect 27950 32952 28906 33008
rect 28962 32952 28967 33008
rect 20069 32950 28967 32952
rect 20069 32947 20135 32950
rect 27889 32947 27955 32950
rect 28901 32947 28967 32950
rect 4337 32874 4403 32877
rect 6269 32874 6335 32877
rect 4337 32872 6335 32874
rect 4337 32816 4342 32872
rect 4398 32816 6274 32872
rect 6330 32816 6335 32872
rect 4337 32814 6335 32816
rect 4337 32811 4403 32814
rect 6269 32811 6335 32814
rect 20253 32874 20319 32877
rect 23841 32874 23907 32877
rect 20253 32872 23907 32874
rect 20253 32816 20258 32872
rect 20314 32816 23846 32872
rect 23902 32816 23907 32872
rect 20253 32814 23907 32816
rect 20253 32811 20319 32814
rect 23841 32811 23907 32814
rect 24025 32874 24091 32877
rect 27245 32874 27311 32877
rect 24025 32872 27311 32874
rect 24025 32816 24030 32872
rect 24086 32816 27250 32872
rect 27306 32816 27311 32872
rect 24025 32814 27311 32816
rect 24025 32811 24091 32814
rect 27245 32811 27311 32814
rect 0 32738 800 32768
rect 1301 32738 1367 32741
rect 0 32736 1367 32738
rect 0 32680 1306 32736
rect 1362 32680 1367 32736
rect 0 32678 1367 32680
rect 0 32648 800 32678
rect 1301 32675 1367 32678
rect 26417 32738 26483 32741
rect 28349 32738 28415 32741
rect 26417 32736 28415 32738
rect 26417 32680 26422 32736
rect 26478 32680 28354 32736
rect 28410 32680 28415 32736
rect 26417 32678 28415 32680
rect 26417 32675 26483 32678
rect 28349 32675 28415 32678
rect 28625 32738 28691 32741
rect 31109 32738 31175 32741
rect 28625 32736 31175 32738
rect 28625 32680 28630 32736
rect 28686 32680 31114 32736
rect 31170 32680 31175 32736
rect 28625 32678 31175 32680
rect 28625 32675 28691 32678
rect 31109 32675 31175 32678
rect 31293 32738 31359 32741
rect 32213 32738 32279 32741
rect 31293 32736 32279 32738
rect 31293 32680 31298 32736
rect 31354 32680 32218 32736
rect 32274 32680 32279 32736
rect 31293 32678 32279 32680
rect 31293 32675 31359 32678
rect 32213 32675 32279 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 9765 32602 9831 32605
rect 21817 32602 21883 32605
rect 22461 32602 22527 32605
rect 9765 32600 9874 32602
rect 9765 32544 9770 32600
rect 9826 32544 9874 32600
rect 9765 32539 9874 32544
rect 21817 32600 22527 32602
rect 21817 32544 21822 32600
rect 21878 32544 22466 32600
rect 22522 32544 22527 32600
rect 21817 32542 22527 32544
rect 21817 32539 21883 32542
rect 22461 32539 22527 32542
rect 23657 32602 23723 32605
rect 28165 32602 28231 32605
rect 23657 32600 28231 32602
rect 23657 32544 23662 32600
rect 23718 32544 28170 32600
rect 28226 32544 28231 32600
rect 23657 32542 28231 32544
rect 23657 32539 23723 32542
rect 28165 32539 28231 32542
rect 30189 32602 30255 32605
rect 31845 32602 31911 32605
rect 30189 32600 31911 32602
rect 30189 32544 30194 32600
rect 30250 32544 31850 32600
rect 31906 32544 31911 32600
rect 30189 32542 31911 32544
rect 30189 32539 30255 32542
rect 31845 32539 31911 32542
rect 4981 32466 5047 32469
rect 6821 32466 6887 32469
rect 4981 32464 6887 32466
rect 4981 32408 4986 32464
rect 5042 32408 6826 32464
rect 6882 32408 6887 32464
rect 4981 32406 6887 32408
rect 4981 32403 5047 32406
rect 6821 32403 6887 32406
rect 9814 32333 9874 32539
rect 19885 32466 19951 32469
rect 22093 32466 22159 32469
rect 19885 32464 22159 32466
rect 19885 32408 19890 32464
rect 19946 32408 22098 32464
rect 22154 32408 22159 32464
rect 19885 32406 22159 32408
rect 19885 32403 19951 32406
rect 22093 32403 22159 32406
rect 22277 32466 22343 32469
rect 24301 32466 24367 32469
rect 22277 32464 24367 32466
rect 22277 32408 22282 32464
rect 22338 32408 24306 32464
rect 24362 32408 24367 32464
rect 22277 32406 24367 32408
rect 22277 32403 22343 32406
rect 24301 32403 24367 32406
rect 24669 32466 24735 32469
rect 26693 32466 26759 32469
rect 28165 32466 28231 32469
rect 31569 32466 31635 32469
rect 34421 32466 34487 32469
rect 24669 32464 34487 32466
rect 24669 32408 24674 32464
rect 24730 32408 26698 32464
rect 26754 32408 28170 32464
rect 28226 32408 31574 32464
rect 31630 32408 34426 32464
rect 34482 32408 34487 32464
rect 24669 32406 34487 32408
rect 24669 32403 24735 32406
rect 26693 32403 26759 32406
rect 28165 32403 28231 32406
rect 31569 32403 31635 32406
rect 34421 32403 34487 32406
rect 4654 32268 4660 32332
rect 4724 32330 4730 32332
rect 5073 32330 5139 32333
rect 4724 32328 5139 32330
rect 4724 32272 5078 32328
rect 5134 32272 5139 32328
rect 4724 32270 5139 32272
rect 4724 32268 4730 32270
rect 5073 32267 5139 32270
rect 5257 32330 5323 32333
rect 6177 32330 6243 32333
rect 5257 32328 6243 32330
rect 5257 32272 5262 32328
rect 5318 32272 6182 32328
rect 6238 32272 6243 32328
rect 5257 32270 6243 32272
rect 5257 32267 5323 32270
rect 6177 32267 6243 32270
rect 9765 32328 9874 32333
rect 9765 32272 9770 32328
rect 9826 32272 9874 32328
rect 9765 32270 9874 32272
rect 21633 32330 21699 32333
rect 22921 32330 22987 32333
rect 25589 32330 25655 32333
rect 21633 32328 25655 32330
rect 21633 32272 21638 32328
rect 21694 32272 22926 32328
rect 22982 32272 25594 32328
rect 25650 32272 25655 32328
rect 21633 32270 25655 32272
rect 9765 32267 9831 32270
rect 21633 32267 21699 32270
rect 22921 32267 22987 32270
rect 25589 32267 25655 32270
rect 28257 32330 28323 32333
rect 30649 32330 30715 32333
rect 28257 32328 30715 32330
rect 28257 32272 28262 32328
rect 28318 32272 30654 32328
rect 30710 32272 30715 32328
rect 28257 32270 30715 32272
rect 28257 32267 28323 32270
rect 30649 32267 30715 32270
rect 31017 32330 31083 32333
rect 32397 32330 32463 32333
rect 32581 32330 32647 32333
rect 31017 32328 32647 32330
rect 31017 32272 31022 32328
rect 31078 32272 32402 32328
rect 32458 32272 32586 32328
rect 32642 32272 32647 32328
rect 31017 32270 32647 32272
rect 31017 32267 31083 32270
rect 32397 32267 32463 32270
rect 32581 32267 32647 32270
rect 30373 32194 30439 32197
rect 31937 32194 32003 32197
rect 30373 32192 32003 32194
rect 30373 32136 30378 32192
rect 30434 32136 31942 32192
rect 31998 32136 32003 32192
rect 30373 32134 32003 32136
rect 30373 32131 30439 32134
rect 31937 32131 32003 32134
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 2405 32058 2471 32061
rect 0 32056 2471 32058
rect 0 32000 2410 32056
rect 2466 32000 2471 32056
rect 0 31998 2471 32000
rect 0 31968 800 31998
rect 2405 31995 2471 31998
rect 8017 32058 8083 32061
rect 8477 32058 8543 32061
rect 9581 32058 9647 32061
rect 8017 32056 9647 32058
rect 8017 32000 8022 32056
rect 8078 32000 8482 32056
rect 8538 32000 9586 32056
rect 9642 32000 9647 32056
rect 8017 31998 9647 32000
rect 8017 31995 8083 31998
rect 8477 31995 8543 31998
rect 9581 31995 9647 31998
rect 13302 31996 13308 32060
rect 13372 32058 13378 32060
rect 13721 32058 13787 32061
rect 26417 32060 26483 32061
rect 26366 32058 26372 32060
rect 13372 32056 26372 32058
rect 26436 32058 26483 32060
rect 29913 32058 29979 32061
rect 30465 32058 30531 32061
rect 26436 32056 26564 32058
rect 13372 32000 13726 32056
rect 13782 32000 26372 32056
rect 26478 32000 26564 32056
rect 13372 31998 26372 32000
rect 13372 31996 13378 31998
rect 13721 31995 13787 31998
rect 26366 31996 26372 31998
rect 26436 31998 26564 32000
rect 29913 32056 30531 32058
rect 29913 32000 29918 32056
rect 29974 32000 30470 32056
rect 30526 32000 30531 32056
rect 29913 31998 30531 32000
rect 26436 31996 26483 31998
rect 26417 31995 26483 31996
rect 29913 31995 29979 31998
rect 30465 31995 30531 31998
rect 30833 32058 30899 32061
rect 32213 32058 32279 32061
rect 32581 32058 32647 32061
rect 30833 32056 32647 32058
rect 30833 32000 30838 32056
rect 30894 32000 32218 32056
rect 32274 32000 32586 32056
rect 32642 32000 32647 32056
rect 30833 31998 32647 32000
rect 30833 31995 30899 31998
rect 32213 31995 32279 31998
rect 32581 31995 32647 31998
rect 9673 31922 9739 31925
rect 10961 31922 11027 31925
rect 9673 31920 11027 31922
rect 9673 31864 9678 31920
rect 9734 31864 10966 31920
rect 11022 31864 11027 31920
rect 9673 31862 11027 31864
rect 9673 31859 9739 31862
rect 10961 31859 11027 31862
rect 15510 31860 15516 31924
rect 15580 31922 15586 31924
rect 15929 31922 15995 31925
rect 15580 31920 15995 31922
rect 15580 31864 15934 31920
rect 15990 31864 15995 31920
rect 15580 31862 15995 31864
rect 15580 31860 15586 31862
rect 15929 31859 15995 31862
rect 25086 31862 27906 31922
rect 5574 31724 5580 31788
rect 5644 31786 5650 31788
rect 5717 31786 5783 31789
rect 5644 31784 5783 31786
rect 5644 31728 5722 31784
rect 5778 31728 5783 31784
rect 5644 31726 5783 31728
rect 5644 31724 5650 31726
rect 5717 31723 5783 31726
rect 14958 31724 14964 31788
rect 15028 31786 15034 31788
rect 15101 31786 15167 31789
rect 15028 31784 15167 31786
rect 15028 31728 15106 31784
rect 15162 31728 15167 31784
rect 15028 31726 15167 31728
rect 15028 31724 15034 31726
rect 15101 31723 15167 31726
rect 23749 31786 23815 31789
rect 25086 31786 25146 31862
rect 26693 31786 26759 31789
rect 23749 31784 25146 31786
rect 23749 31728 23754 31784
rect 23810 31728 25146 31784
rect 23749 31726 25146 31728
rect 25270 31784 26759 31786
rect 25270 31728 26698 31784
rect 26754 31728 26759 31784
rect 25270 31726 26759 31728
rect 23749 31723 23815 31726
rect 25270 31653 25330 31726
rect 26693 31723 26759 31726
rect 27061 31786 27127 31789
rect 27613 31788 27679 31789
rect 27470 31786 27476 31788
rect 27061 31784 27476 31786
rect 27061 31728 27066 31784
rect 27122 31728 27476 31784
rect 27061 31726 27476 31728
rect 27061 31723 27127 31726
rect 27470 31724 27476 31726
rect 27540 31724 27546 31788
rect 27613 31784 27660 31788
rect 27724 31786 27730 31788
rect 27846 31786 27906 31862
rect 29177 31786 29243 31789
rect 29545 31786 29611 31789
rect 27613 31728 27618 31784
rect 27613 31724 27660 31728
rect 27724 31726 27770 31786
rect 27846 31784 29611 31786
rect 27846 31728 29182 31784
rect 29238 31728 29550 31784
rect 29606 31728 29611 31784
rect 27846 31726 29611 31728
rect 27724 31724 27730 31726
rect 27613 31723 27679 31724
rect 29177 31723 29243 31726
rect 29545 31723 29611 31726
rect 5441 31650 5507 31653
rect 5574 31650 5580 31652
rect 5441 31648 5580 31650
rect 5441 31592 5446 31648
rect 5502 31592 5580 31648
rect 5441 31590 5580 31592
rect 5441 31587 5507 31590
rect 5574 31588 5580 31590
rect 5644 31588 5650 31652
rect 6269 31650 6335 31653
rect 6637 31650 6703 31653
rect 6269 31648 6703 31650
rect 6269 31592 6274 31648
rect 6330 31592 6642 31648
rect 6698 31592 6703 31648
rect 6269 31590 6703 31592
rect 6269 31587 6335 31590
rect 6637 31587 6703 31590
rect 22553 31650 22619 31653
rect 24025 31650 24091 31653
rect 24945 31650 25011 31653
rect 22553 31648 24091 31650
rect 22553 31592 22558 31648
rect 22614 31592 24030 31648
rect 24086 31592 24091 31648
rect 22553 31590 24091 31592
rect 22553 31587 22619 31590
rect 24025 31587 24091 31590
rect 24166 31648 25011 31650
rect 24166 31592 24950 31648
rect 25006 31592 25011 31648
rect 24166 31590 25011 31592
rect 25270 31648 25379 31653
rect 25270 31592 25318 31648
rect 25374 31592 25379 31648
rect 25270 31590 25379 31592
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 23013 31514 23079 31517
rect 24166 31514 24226 31590
rect 24945 31587 25011 31590
rect 25313 31587 25379 31590
rect 26233 31650 26299 31653
rect 26969 31650 27035 31653
rect 27429 31650 27495 31653
rect 28257 31652 28323 31653
rect 26233 31648 27495 31650
rect 26233 31592 26238 31648
rect 26294 31592 26974 31648
rect 27030 31592 27434 31648
rect 27490 31592 27495 31648
rect 26233 31590 27495 31592
rect 26233 31587 26299 31590
rect 26969 31587 27035 31590
rect 27429 31587 27495 31590
rect 28206 31588 28212 31652
rect 28276 31650 28323 31652
rect 28809 31650 28875 31653
rect 30465 31650 30531 31653
rect 28276 31648 28368 31650
rect 28318 31592 28368 31648
rect 28276 31590 28368 31592
rect 28809 31648 30531 31650
rect 28809 31592 28814 31648
rect 28870 31592 30470 31648
rect 30526 31592 30531 31648
rect 28809 31590 30531 31592
rect 28276 31588 28323 31590
rect 28257 31587 28323 31588
rect 28809 31587 28875 31590
rect 30465 31587 30531 31590
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 23013 31512 24226 31514
rect 23013 31456 23018 31512
rect 23074 31456 24226 31512
rect 23013 31454 24226 31456
rect 24485 31514 24551 31517
rect 25681 31514 25747 31517
rect 27245 31516 27311 31517
rect 27245 31514 27292 31516
rect 24485 31512 25747 31514
rect 24485 31456 24490 31512
rect 24546 31456 25686 31512
rect 25742 31456 25747 31512
rect 24485 31454 25747 31456
rect 27200 31512 27292 31514
rect 27356 31514 27362 31516
rect 30189 31514 30255 31517
rect 27356 31512 30255 31514
rect 27200 31456 27250 31512
rect 27356 31456 30194 31512
rect 30250 31456 30255 31512
rect 27200 31454 27292 31456
rect 23013 31451 23079 31454
rect 24485 31451 24551 31454
rect 25681 31451 25747 31454
rect 27245 31452 27292 31454
rect 27356 31454 30255 31456
rect 27356 31452 27362 31454
rect 27245 31451 27311 31452
rect 30189 31451 30255 31454
rect 0 31378 800 31408
rect 1301 31378 1367 31381
rect 0 31376 1367 31378
rect 0 31320 1306 31376
rect 1362 31320 1367 31376
rect 0 31318 1367 31320
rect 0 31288 800 31318
rect 1301 31315 1367 31318
rect 28073 31378 28139 31381
rect 28257 31378 28323 31381
rect 28073 31376 28323 31378
rect 28073 31320 28078 31376
rect 28134 31320 28262 31376
rect 28318 31320 28323 31376
rect 28073 31318 28323 31320
rect 28073 31315 28139 31318
rect 28257 31315 28323 31318
rect 5717 31242 5783 31245
rect 8569 31242 8635 31245
rect 5717 31240 8635 31242
rect 5717 31184 5722 31240
rect 5778 31184 8574 31240
rect 8630 31184 8635 31240
rect 5717 31182 8635 31184
rect 5717 31179 5783 31182
rect 8569 31179 8635 31182
rect 12065 31242 12131 31245
rect 15377 31244 15443 31245
rect 15326 31242 15332 31244
rect 12065 31240 15332 31242
rect 15396 31242 15443 31244
rect 15561 31242 15627 31245
rect 30281 31242 30347 31245
rect 15396 31240 15488 31242
rect 12065 31184 12070 31240
rect 12126 31184 15332 31240
rect 15438 31184 15488 31240
rect 12065 31182 15332 31184
rect 12065 31179 12131 31182
rect 15326 31180 15332 31182
rect 15396 31182 15488 31184
rect 15561 31240 30347 31242
rect 15561 31184 15566 31240
rect 15622 31184 30286 31240
rect 30342 31184 30347 31240
rect 15561 31182 30347 31184
rect 15396 31180 15443 31182
rect 15377 31179 15443 31180
rect 15561 31179 15627 31182
rect 30281 31179 30347 31182
rect 13537 31106 13603 31109
rect 26233 31106 26299 31109
rect 13537 31104 26299 31106
rect 13537 31048 13542 31104
rect 13598 31048 26238 31104
rect 26294 31048 26299 31104
rect 13537 31046 26299 31048
rect 13537 31043 13603 31046
rect 26233 31043 26299 31046
rect 26601 31106 26667 31109
rect 28073 31106 28139 31109
rect 26601 31104 28139 31106
rect 26601 31048 26606 31104
rect 26662 31048 28078 31104
rect 28134 31048 28139 31104
rect 26601 31046 28139 31048
rect 26601 31043 26667 31046
rect 28073 31043 28139 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 5717 30970 5783 30973
rect 9121 30970 9187 30973
rect 5717 30968 9187 30970
rect 5717 30912 5722 30968
rect 5778 30912 9126 30968
rect 9182 30912 9187 30968
rect 5717 30910 9187 30912
rect 5717 30907 5783 30910
rect 9121 30907 9187 30910
rect 23473 30970 23539 30973
rect 28533 30970 28599 30973
rect 23473 30968 28599 30970
rect 23473 30912 23478 30968
rect 23534 30912 28538 30968
rect 28594 30912 28599 30968
rect 23473 30910 28599 30912
rect 23473 30907 23539 30910
rect 28533 30907 28599 30910
rect 4429 30834 4495 30837
rect 9489 30834 9555 30837
rect 4429 30832 9555 30834
rect 4429 30776 4434 30832
rect 4490 30776 9494 30832
rect 9550 30776 9555 30832
rect 4429 30774 9555 30776
rect 4429 30771 4495 30774
rect 9489 30771 9555 30774
rect 16205 30834 16271 30837
rect 16481 30834 16547 30837
rect 16205 30832 16547 30834
rect 16205 30776 16210 30832
rect 16266 30776 16486 30832
rect 16542 30776 16547 30832
rect 16205 30774 16547 30776
rect 16205 30771 16271 30774
rect 16481 30771 16547 30774
rect 26601 30834 26667 30837
rect 27337 30834 27403 30837
rect 26601 30832 27403 30834
rect 26601 30776 26606 30832
rect 26662 30776 27342 30832
rect 27398 30776 27403 30832
rect 26601 30774 27403 30776
rect 26601 30771 26667 30774
rect 27337 30771 27403 30774
rect 27613 30834 27679 30837
rect 28717 30834 28783 30837
rect 27613 30832 28783 30834
rect 27613 30776 27618 30832
rect 27674 30776 28722 30832
rect 28778 30776 28783 30832
rect 27613 30774 28783 30776
rect 27613 30771 27679 30774
rect 28717 30771 28783 30774
rect 0 30698 800 30728
rect 3141 30698 3207 30701
rect 0 30696 3207 30698
rect 0 30640 3146 30696
rect 3202 30640 3207 30696
rect 0 30638 3207 30640
rect 0 30608 800 30638
rect 3141 30635 3207 30638
rect 4521 30698 4587 30701
rect 4981 30698 5047 30701
rect 27613 30698 27679 30701
rect 27981 30698 28047 30701
rect 4521 30696 6378 30698
rect 4521 30640 4526 30696
rect 4582 30640 4986 30696
rect 5042 30640 6378 30696
rect 4521 30638 6378 30640
rect 4521 30635 4587 30638
rect 4981 30635 5047 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 6318 30428 6378 30638
rect 27613 30696 28047 30698
rect 27613 30640 27618 30696
rect 27674 30640 27986 30696
rect 28042 30640 28047 30696
rect 27613 30638 28047 30640
rect 27613 30635 27679 30638
rect 27981 30635 28047 30638
rect 16205 30562 16271 30565
rect 16389 30562 16455 30565
rect 17861 30562 17927 30565
rect 19609 30562 19675 30565
rect 16205 30560 19675 30562
rect 16205 30504 16210 30560
rect 16266 30504 16394 30560
rect 16450 30504 17866 30560
rect 17922 30504 19614 30560
rect 19670 30504 19675 30560
rect 16205 30502 19675 30504
rect 16205 30499 16271 30502
rect 16389 30499 16455 30502
rect 17861 30499 17927 30502
rect 19609 30499 19675 30502
rect 21357 30562 21423 30565
rect 24853 30562 24919 30565
rect 21357 30560 24919 30562
rect 21357 30504 21362 30560
rect 21418 30504 24858 30560
rect 24914 30504 24919 30560
rect 21357 30502 24919 30504
rect 21357 30499 21423 30502
rect 24853 30499 24919 30502
rect 27429 30562 27495 30565
rect 30833 30562 30899 30565
rect 27429 30560 30899 30562
rect 27429 30504 27434 30560
rect 27490 30504 30838 30560
rect 30894 30504 30899 30560
rect 27429 30502 30899 30504
rect 27429 30499 27495 30502
rect 30833 30499 30899 30502
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 6310 30364 6316 30428
rect 6380 30426 6386 30428
rect 6453 30426 6519 30429
rect 15561 30426 15627 30429
rect 6380 30424 6519 30426
rect 6380 30368 6458 30424
rect 6514 30368 6519 30424
rect 6380 30366 6519 30368
rect 6380 30364 6386 30366
rect 6453 30363 6519 30366
rect 15150 30424 15627 30426
rect 15150 30368 15566 30424
rect 15622 30368 15627 30424
rect 15150 30366 15627 30368
rect 9121 30290 9187 30293
rect 13077 30292 13143 30293
rect 9622 30290 9628 30292
rect 9121 30288 9628 30290
rect 9121 30232 9126 30288
rect 9182 30232 9628 30288
rect 9121 30230 9628 30232
rect 9121 30227 9187 30230
rect 9622 30228 9628 30230
rect 9692 30228 9698 30292
rect 13077 30290 13124 30292
rect 13036 30288 13124 30290
rect 13188 30290 13194 30292
rect 15150 30290 15210 30366
rect 15561 30363 15627 30366
rect 26233 30426 26299 30429
rect 26601 30426 26667 30429
rect 34053 30426 34119 30429
rect 26233 30424 34119 30426
rect 26233 30368 26238 30424
rect 26294 30368 26606 30424
rect 26662 30368 34058 30424
rect 34114 30368 34119 30424
rect 26233 30366 34119 30368
rect 26233 30363 26299 30366
rect 26601 30363 26667 30366
rect 34053 30363 34119 30366
rect 13036 30232 13082 30288
rect 13036 30230 13124 30232
rect 13077 30228 13124 30230
rect 13188 30230 15210 30290
rect 22001 30290 22067 30293
rect 23565 30290 23631 30293
rect 22001 30288 23631 30290
rect 22001 30232 22006 30288
rect 22062 30232 23570 30288
rect 23626 30232 23631 30288
rect 22001 30230 23631 30232
rect 13188 30228 13194 30230
rect 13077 30227 13143 30228
rect 22001 30227 22067 30230
rect 23565 30227 23631 30230
rect 26601 30290 26667 30293
rect 27245 30290 27311 30293
rect 27705 30290 27771 30293
rect 26601 30288 27771 30290
rect 26601 30232 26606 30288
rect 26662 30232 27250 30288
rect 27306 30232 27710 30288
rect 27766 30232 27771 30288
rect 26601 30230 27771 30232
rect 26601 30227 26667 30230
rect 27245 30227 27311 30230
rect 27705 30227 27771 30230
rect 28257 30290 28323 30293
rect 28901 30290 28967 30293
rect 28257 30288 28967 30290
rect 28257 30232 28262 30288
rect 28318 30232 28906 30288
rect 28962 30232 28967 30288
rect 28257 30230 28967 30232
rect 28257 30227 28323 30230
rect 28901 30227 28967 30230
rect 29361 30290 29427 30293
rect 31109 30290 31175 30293
rect 29361 30288 31175 30290
rect 29361 30232 29366 30288
rect 29422 30232 31114 30288
rect 31170 30232 31175 30288
rect 29361 30230 31175 30232
rect 29361 30227 29427 30230
rect 31109 30227 31175 30230
rect 9070 30092 9076 30156
rect 9140 30154 9146 30156
rect 9581 30154 9647 30157
rect 9140 30152 9647 30154
rect 9140 30096 9586 30152
rect 9642 30096 9647 30152
rect 9140 30094 9647 30096
rect 9140 30092 9146 30094
rect 9581 30091 9647 30094
rect 11053 30154 11119 30157
rect 11789 30154 11855 30157
rect 12198 30154 12204 30156
rect 11053 30152 12204 30154
rect 11053 30096 11058 30152
rect 11114 30096 11794 30152
rect 11850 30096 12204 30152
rect 11053 30094 12204 30096
rect 11053 30091 11119 30094
rect 11789 30091 11855 30094
rect 12198 30092 12204 30094
rect 12268 30092 12274 30156
rect 14089 30154 14155 30157
rect 23749 30156 23815 30157
rect 23749 30154 23796 30156
rect 14089 30152 19350 30154
rect 14089 30096 14094 30152
rect 14150 30096 19350 30152
rect 14089 30094 19350 30096
rect 23704 30152 23796 30154
rect 23704 30096 23754 30152
rect 23704 30094 23796 30096
rect 14089 30091 14155 30094
rect 0 30018 800 30048
rect 1301 30018 1367 30021
rect 0 30016 1367 30018
rect 0 29960 1306 30016
rect 1362 29960 1367 30016
rect 0 29958 1367 29960
rect 19290 30018 19350 30094
rect 23749 30092 23796 30094
rect 23860 30092 23866 30156
rect 27470 30092 27476 30156
rect 27540 30154 27546 30156
rect 29177 30154 29243 30157
rect 27540 30152 29243 30154
rect 27540 30096 29182 30152
rect 29238 30096 29243 30152
rect 27540 30094 29243 30096
rect 27540 30092 27546 30094
rect 23749 30091 23815 30092
rect 29177 30091 29243 30094
rect 28073 30018 28139 30021
rect 30649 30018 30715 30021
rect 31017 30018 31083 30021
rect 19290 30016 31083 30018
rect 19290 29960 28078 30016
rect 28134 29960 30654 30016
rect 30710 29960 31022 30016
rect 31078 29960 31083 30016
rect 19290 29958 31083 29960
rect 0 29928 800 29958
rect 1301 29955 1367 29958
rect 28073 29955 28139 29958
rect 30649 29955 30715 29958
rect 31017 29955 31083 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 5349 29882 5415 29885
rect 9305 29882 9371 29885
rect 5349 29880 9371 29882
rect 5349 29824 5354 29880
rect 5410 29824 9310 29880
rect 9366 29824 9371 29880
rect 5349 29822 9371 29824
rect 5349 29819 5415 29822
rect 9305 29819 9371 29822
rect 16665 29882 16731 29885
rect 16941 29882 17007 29885
rect 22737 29882 22803 29885
rect 16665 29880 22803 29882
rect 16665 29824 16670 29880
rect 16726 29824 16946 29880
rect 17002 29824 22742 29880
rect 22798 29824 22803 29880
rect 16665 29822 22803 29824
rect 16665 29819 16731 29822
rect 16941 29819 17007 29822
rect 22737 29819 22803 29822
rect 27797 29882 27863 29885
rect 28073 29882 28139 29885
rect 27797 29880 28139 29882
rect 27797 29824 27802 29880
rect 27858 29824 28078 29880
rect 28134 29824 28139 29880
rect 27797 29822 28139 29824
rect 27797 29819 27863 29822
rect 28073 29819 28139 29822
rect 7281 29746 7347 29749
rect 9121 29746 9187 29749
rect 26182 29746 26188 29748
rect 7281 29744 9187 29746
rect 7281 29688 7286 29744
rect 7342 29688 9126 29744
rect 9182 29688 9187 29744
rect 7281 29686 9187 29688
rect 7281 29683 7347 29686
rect 9121 29683 9187 29686
rect 19290 29686 26188 29746
rect 13353 29610 13419 29613
rect 13721 29610 13787 29613
rect 19290 29610 19350 29686
rect 26182 29684 26188 29686
rect 26252 29746 26258 29748
rect 27705 29746 27771 29749
rect 28206 29746 28212 29748
rect 26252 29744 28212 29746
rect 26252 29688 27710 29744
rect 27766 29688 28212 29744
rect 26252 29686 28212 29688
rect 26252 29684 26258 29686
rect 27705 29683 27771 29686
rect 28206 29684 28212 29686
rect 28276 29746 28282 29748
rect 28441 29746 28507 29749
rect 28276 29744 28507 29746
rect 28276 29688 28446 29744
rect 28502 29688 28507 29744
rect 28276 29686 28507 29688
rect 28276 29684 28282 29686
rect 28441 29683 28507 29686
rect 13353 29608 19350 29610
rect 13353 29552 13358 29608
rect 13414 29552 13726 29608
rect 13782 29552 19350 29608
rect 13353 29550 19350 29552
rect 20989 29610 21055 29613
rect 24158 29610 24164 29612
rect 20989 29608 24164 29610
rect 20989 29552 20994 29608
rect 21050 29552 24164 29608
rect 20989 29550 24164 29552
rect 13353 29547 13419 29550
rect 13721 29547 13787 29550
rect 20989 29547 21055 29550
rect 24158 29548 24164 29550
rect 24228 29548 24234 29612
rect 26233 29610 26299 29613
rect 27981 29610 28047 29613
rect 28257 29610 28323 29613
rect 26233 29608 28323 29610
rect 26233 29552 26238 29608
rect 26294 29552 27986 29608
rect 28042 29552 28262 29608
rect 28318 29552 28323 29608
rect 26233 29550 28323 29552
rect 26233 29547 26299 29550
rect 27981 29547 28047 29550
rect 28257 29547 28323 29550
rect 30741 29610 30807 29613
rect 30966 29610 30972 29612
rect 30741 29608 30972 29610
rect 30741 29552 30746 29608
rect 30802 29552 30972 29608
rect 30741 29550 30972 29552
rect 30741 29547 30807 29550
rect 30966 29548 30972 29550
rect 31036 29548 31042 29612
rect 9990 29412 9996 29476
rect 10060 29474 10066 29476
rect 10225 29474 10291 29477
rect 10060 29472 10291 29474
rect 10060 29416 10230 29472
rect 10286 29416 10291 29472
rect 10060 29414 10291 29416
rect 10060 29412 10066 29414
rect 10225 29411 10291 29414
rect 19609 29474 19675 29477
rect 21725 29474 21791 29477
rect 25221 29476 25287 29477
rect 27337 29476 27403 29477
rect 25221 29474 25268 29476
rect 19609 29472 21791 29474
rect 19609 29416 19614 29472
rect 19670 29416 21730 29472
rect 21786 29416 21791 29472
rect 19609 29414 21791 29416
rect 25176 29472 25268 29474
rect 25176 29416 25226 29472
rect 25176 29414 25268 29416
rect 19609 29411 19675 29414
rect 21725 29411 21791 29414
rect 25221 29412 25268 29414
rect 25332 29412 25338 29476
rect 27286 29474 27292 29476
rect 27246 29414 27292 29474
rect 27356 29472 27403 29476
rect 27398 29416 27403 29472
rect 27286 29412 27292 29414
rect 27356 29412 27403 29416
rect 25221 29411 25287 29412
rect 27337 29411 27403 29412
rect 27705 29474 27771 29477
rect 30373 29474 30439 29477
rect 31661 29474 31727 29477
rect 27705 29472 31727 29474
rect 27705 29416 27710 29472
rect 27766 29416 30378 29472
rect 30434 29416 31666 29472
rect 31722 29416 31727 29472
rect 27705 29414 31727 29416
rect 27705 29411 27771 29414
rect 30373 29411 30439 29414
rect 31661 29411 31727 29414
rect 4870 29408 5186 29409
rect 0 29338 800 29368
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 1301 29338 1367 29341
rect 0 29336 1367 29338
rect 0 29280 1306 29336
rect 1362 29280 1367 29336
rect 0 29278 1367 29280
rect 0 29248 800 29278
rect 1301 29275 1367 29278
rect 12709 29338 12775 29341
rect 13077 29338 13143 29341
rect 13629 29338 13695 29341
rect 12709 29336 13695 29338
rect 12709 29280 12714 29336
rect 12770 29280 13082 29336
rect 13138 29280 13634 29336
rect 13690 29280 13695 29336
rect 12709 29278 13695 29280
rect 12709 29275 12775 29278
rect 13077 29275 13143 29278
rect 13629 29275 13695 29278
rect 21265 29338 21331 29341
rect 25589 29338 25655 29341
rect 21265 29336 25655 29338
rect 21265 29280 21270 29336
rect 21326 29280 25594 29336
rect 25650 29280 25655 29336
rect 21265 29278 25655 29280
rect 21265 29275 21331 29278
rect 25589 29275 25655 29278
rect 1945 29202 2011 29205
rect 5717 29202 5783 29205
rect 1945 29200 5783 29202
rect 1945 29144 1950 29200
rect 2006 29144 5722 29200
rect 5778 29144 5783 29200
rect 1945 29142 5783 29144
rect 1945 29139 2011 29142
rect 5717 29139 5783 29142
rect 11094 29140 11100 29204
rect 11164 29202 11170 29204
rect 13445 29202 13511 29205
rect 11164 29200 13511 29202
rect 11164 29144 13450 29200
rect 13506 29144 13511 29200
rect 11164 29142 13511 29144
rect 11164 29140 11170 29142
rect 13445 29139 13511 29142
rect 13997 29204 14063 29205
rect 13997 29200 14044 29204
rect 14108 29202 14114 29204
rect 17217 29202 17283 29205
rect 18229 29202 18295 29205
rect 13997 29144 14002 29200
rect 13997 29140 14044 29144
rect 14108 29142 14154 29202
rect 17217 29200 18295 29202
rect 17217 29144 17222 29200
rect 17278 29144 18234 29200
rect 18290 29144 18295 29200
rect 17217 29142 18295 29144
rect 14108 29140 14114 29142
rect 13997 29139 14063 29140
rect 17217 29139 17283 29142
rect 18229 29139 18295 29142
rect 21541 29202 21607 29205
rect 23289 29202 23355 29205
rect 21541 29200 23355 29202
rect 21541 29144 21546 29200
rect 21602 29144 23294 29200
rect 23350 29144 23355 29200
rect 21541 29142 23355 29144
rect 21541 29139 21607 29142
rect 23289 29139 23355 29142
rect 28257 29202 28323 29205
rect 31477 29202 31543 29205
rect 28257 29200 31543 29202
rect 28257 29144 28262 29200
rect 28318 29144 31482 29200
rect 31538 29144 31543 29200
rect 28257 29142 31543 29144
rect 28257 29139 28323 29142
rect 31477 29139 31543 29142
rect 13854 29004 13860 29068
rect 13924 29066 13930 29068
rect 14917 29066 14983 29069
rect 13924 29064 14983 29066
rect 13924 29008 14922 29064
rect 14978 29008 14983 29064
rect 13924 29006 14983 29008
rect 13924 29004 13930 29006
rect 14917 29003 14983 29006
rect 15142 29004 15148 29068
rect 15212 29066 15218 29068
rect 15377 29066 15443 29069
rect 15212 29064 15443 29066
rect 15212 29008 15382 29064
rect 15438 29008 15443 29064
rect 15212 29006 15443 29008
rect 15212 29004 15218 29006
rect 15377 29003 15443 29006
rect 18965 29066 19031 29069
rect 30005 29068 30071 29069
rect 19190 29066 19196 29068
rect 18965 29064 19196 29066
rect 18965 29008 18970 29064
rect 19026 29008 19196 29064
rect 18965 29006 19196 29008
rect 18965 29003 19031 29006
rect 19190 29004 19196 29006
rect 19260 29004 19266 29068
rect 30005 29066 30052 29068
rect 29960 29064 30052 29066
rect 29960 29008 30010 29064
rect 29960 29006 30052 29008
rect 30005 29004 30052 29006
rect 30116 29004 30122 29068
rect 33409 29066 33475 29069
rect 33542 29066 33548 29068
rect 33409 29064 33548 29066
rect 33409 29008 33414 29064
rect 33470 29008 33548 29064
rect 33409 29006 33548 29008
rect 30005 29003 30071 29004
rect 33409 29003 33475 29006
rect 33542 29004 33548 29006
rect 33612 29004 33618 29068
rect 34278 29004 34284 29068
rect 34348 29066 34354 29068
rect 35801 29066 35867 29069
rect 34348 29064 35867 29066
rect 34348 29008 35806 29064
rect 35862 29008 35867 29064
rect 34348 29006 35867 29008
rect 34348 29004 34354 29006
rect 35801 29003 35867 29006
rect 21081 28930 21147 28933
rect 21909 28930 21975 28933
rect 21081 28928 21975 28930
rect 21081 28872 21086 28928
rect 21142 28872 21914 28928
rect 21970 28872 21975 28928
rect 21081 28870 21975 28872
rect 21081 28867 21147 28870
rect 21909 28867 21975 28870
rect 26969 28930 27035 28933
rect 27654 28930 27660 28932
rect 26969 28928 27660 28930
rect 26969 28872 26974 28928
rect 27030 28872 27660 28928
rect 26969 28870 27660 28872
rect 26969 28867 27035 28870
rect 27654 28868 27660 28870
rect 27724 28930 27730 28932
rect 28441 28930 28507 28933
rect 27724 28928 28507 28930
rect 27724 28872 28446 28928
rect 28502 28872 28507 28928
rect 27724 28870 28507 28872
rect 27724 28868 27730 28870
rect 28441 28867 28507 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 6269 28794 6335 28797
rect 10910 28794 10916 28796
rect 6269 28792 10916 28794
rect 6269 28736 6274 28792
rect 6330 28736 10916 28792
rect 6269 28734 10916 28736
rect 6269 28731 6335 28734
rect 10910 28732 10916 28734
rect 10980 28732 10986 28796
rect 19425 28794 19491 28797
rect 25773 28794 25839 28797
rect 19425 28792 25839 28794
rect 19425 28736 19430 28792
rect 19486 28736 25778 28792
rect 25834 28736 25839 28792
rect 19425 28734 25839 28736
rect 19425 28731 19491 28734
rect 25773 28731 25839 28734
rect 27245 28794 27311 28797
rect 27654 28794 27660 28796
rect 27245 28792 27660 28794
rect 27245 28736 27250 28792
rect 27306 28736 27660 28792
rect 27245 28734 27660 28736
rect 27245 28731 27311 28734
rect 27654 28732 27660 28734
rect 27724 28732 27730 28796
rect 28257 28794 28323 28797
rect 28441 28794 28507 28797
rect 28257 28792 28507 28794
rect 28257 28736 28262 28792
rect 28318 28736 28446 28792
rect 28502 28736 28507 28792
rect 28257 28734 28507 28736
rect 28257 28731 28323 28734
rect 28441 28731 28507 28734
rect 0 28658 800 28688
rect 1301 28658 1367 28661
rect 0 28656 1367 28658
rect 0 28600 1306 28656
rect 1362 28600 1367 28656
rect 0 28598 1367 28600
rect 0 28568 800 28598
rect 1301 28595 1367 28598
rect 21357 28658 21423 28661
rect 29126 28658 29132 28660
rect 21357 28656 29132 28658
rect 21357 28600 21362 28656
rect 21418 28600 29132 28656
rect 21357 28598 29132 28600
rect 21357 28595 21423 28598
rect 29126 28596 29132 28598
rect 29196 28596 29202 28660
rect 5257 28522 5323 28525
rect 12433 28522 12499 28525
rect 5257 28520 12499 28522
rect 5257 28464 5262 28520
rect 5318 28464 12438 28520
rect 12494 28464 12499 28520
rect 5257 28462 12499 28464
rect 5257 28459 5323 28462
rect 12433 28459 12499 28462
rect 15561 28522 15627 28525
rect 15694 28522 15700 28524
rect 15561 28520 15700 28522
rect 15561 28464 15566 28520
rect 15622 28464 15700 28520
rect 15561 28462 15700 28464
rect 15561 28459 15627 28462
rect 15694 28460 15700 28462
rect 15764 28522 15770 28524
rect 16665 28522 16731 28525
rect 15764 28520 16731 28522
rect 15764 28464 16670 28520
rect 16726 28464 16731 28520
rect 15764 28462 16731 28464
rect 15764 28460 15770 28462
rect 16665 28459 16731 28462
rect 18229 28522 18295 28525
rect 24945 28522 25011 28525
rect 18229 28520 25011 28522
rect 18229 28464 18234 28520
rect 18290 28464 24950 28520
rect 25006 28464 25011 28520
rect 18229 28462 25011 28464
rect 18229 28459 18295 28462
rect 18830 28389 18890 28462
rect 24945 28459 25011 28462
rect 25129 28522 25195 28525
rect 28257 28522 28323 28525
rect 25129 28520 28323 28522
rect 25129 28464 25134 28520
rect 25190 28464 28262 28520
rect 28318 28464 28323 28520
rect 25129 28462 28323 28464
rect 25129 28459 25195 28462
rect 28257 28459 28323 28462
rect 18781 28384 18890 28389
rect 18781 28328 18786 28384
rect 18842 28328 18890 28384
rect 18781 28326 18890 28328
rect 21725 28386 21791 28389
rect 30005 28386 30071 28389
rect 21725 28384 30071 28386
rect 21725 28328 21730 28384
rect 21786 28328 30010 28384
rect 30066 28328 30071 28384
rect 21725 28326 30071 28328
rect 18781 28323 18847 28326
rect 21725 28323 21791 28326
rect 30005 28323 30071 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 15469 28250 15535 28253
rect 19241 28250 19307 28253
rect 15469 28248 19307 28250
rect 15469 28192 15474 28248
rect 15530 28192 19246 28248
rect 19302 28192 19307 28248
rect 15469 28190 19307 28192
rect 15469 28187 15535 28190
rect 19241 28187 19307 28190
rect 25405 28250 25471 28253
rect 26366 28250 26372 28252
rect 25405 28248 26372 28250
rect 25405 28192 25410 28248
rect 25466 28192 26372 28248
rect 25405 28190 26372 28192
rect 25405 28187 25471 28190
rect 26366 28188 26372 28190
rect 26436 28250 26442 28252
rect 26877 28250 26943 28253
rect 26436 28248 26943 28250
rect 26436 28192 26882 28248
rect 26938 28192 26943 28248
rect 26436 28190 26943 28192
rect 26436 28188 26442 28190
rect 26877 28187 26943 28190
rect 9765 28114 9831 28117
rect 10777 28114 10843 28117
rect 9765 28112 10843 28114
rect 9765 28056 9770 28112
rect 9826 28056 10782 28112
rect 10838 28056 10843 28112
rect 9765 28054 10843 28056
rect 9765 28051 9831 28054
rect 10777 28051 10843 28054
rect 22921 28114 22987 28117
rect 25998 28114 26004 28116
rect 22921 28112 26004 28114
rect 22921 28056 22926 28112
rect 22982 28056 26004 28112
rect 22921 28054 26004 28056
rect 22921 28051 22987 28054
rect 25998 28052 26004 28054
rect 26068 28114 26074 28116
rect 29913 28114 29979 28117
rect 26068 28112 29979 28114
rect 26068 28056 29918 28112
rect 29974 28056 29979 28112
rect 26068 28054 29979 28056
rect 26068 28052 26074 28054
rect 29913 28051 29979 28054
rect 0 27978 800 28008
rect 1393 27978 1459 27981
rect 0 27976 1459 27978
rect 0 27920 1398 27976
rect 1454 27920 1459 27976
rect 0 27918 1459 27920
rect 0 27888 800 27918
rect 1393 27915 1459 27918
rect 9673 27978 9739 27981
rect 16389 27978 16455 27981
rect 25865 27978 25931 27981
rect 26969 27978 27035 27981
rect 9673 27976 16455 27978
rect 9673 27920 9678 27976
rect 9734 27920 16394 27976
rect 16450 27920 16455 27976
rect 9673 27918 16455 27920
rect 9673 27915 9739 27918
rect 16389 27915 16455 27918
rect 19290 27976 27035 27978
rect 19290 27920 25870 27976
rect 25926 27920 26974 27976
rect 27030 27920 27035 27976
rect 19290 27918 27035 27920
rect 12801 27844 12867 27845
rect 12750 27842 12756 27844
rect 12674 27782 12756 27842
rect 12820 27842 12867 27844
rect 19290 27842 19350 27918
rect 25865 27915 25931 27918
rect 26969 27915 27035 27918
rect 27654 27916 27660 27980
rect 27724 27978 27730 27980
rect 28809 27978 28875 27981
rect 27724 27976 28875 27978
rect 27724 27920 28814 27976
rect 28870 27920 28875 27976
rect 27724 27918 28875 27920
rect 27724 27916 27730 27918
rect 28809 27915 28875 27918
rect 31017 27978 31083 27981
rect 36445 27978 36511 27981
rect 31017 27976 36511 27978
rect 31017 27920 31022 27976
rect 31078 27920 36450 27976
rect 36506 27920 36511 27976
rect 31017 27918 36511 27920
rect 31017 27915 31083 27918
rect 36445 27915 36511 27918
rect 22829 27844 22895 27845
rect 22829 27842 22876 27844
rect 12820 27840 19350 27842
rect 12862 27784 19350 27840
rect 12750 27780 12756 27782
rect 12820 27782 19350 27784
rect 22784 27840 22876 27842
rect 22784 27784 22834 27840
rect 22784 27782 22876 27784
rect 12820 27780 12867 27782
rect 12801 27779 12867 27780
rect 22829 27780 22876 27782
rect 22940 27780 22946 27844
rect 23105 27842 23171 27845
rect 30414 27842 30420 27844
rect 23105 27840 30420 27842
rect 23105 27784 23110 27840
rect 23166 27784 30420 27840
rect 23105 27782 30420 27784
rect 22829 27779 22895 27780
rect 23105 27779 23171 27782
rect 30414 27780 30420 27782
rect 30484 27842 30490 27844
rect 31385 27842 31451 27845
rect 30484 27840 31451 27842
rect 30484 27784 31390 27840
rect 31446 27784 31451 27840
rect 30484 27782 31451 27784
rect 30484 27780 30490 27782
rect 31385 27779 31451 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 7189 27706 7255 27709
rect 7741 27706 7807 27709
rect 7189 27704 7807 27706
rect 7189 27648 7194 27704
rect 7250 27648 7746 27704
rect 7802 27648 7807 27704
rect 7189 27646 7807 27648
rect 7189 27643 7255 27646
rect 7741 27643 7807 27646
rect 18454 27644 18460 27708
rect 18524 27706 18530 27708
rect 18965 27706 19031 27709
rect 18524 27704 19031 27706
rect 18524 27648 18970 27704
rect 19026 27648 19031 27704
rect 18524 27646 19031 27648
rect 18524 27644 18530 27646
rect 18965 27643 19031 27646
rect 19977 27706 20043 27709
rect 24853 27706 24919 27709
rect 27337 27708 27403 27709
rect 19977 27704 27170 27706
rect 19977 27648 19982 27704
rect 20038 27648 24858 27704
rect 24914 27648 27170 27704
rect 19977 27646 27170 27648
rect 19977 27643 20043 27646
rect 24853 27643 24919 27646
rect 9397 27570 9463 27573
rect 9806 27570 9812 27572
rect 9397 27568 9812 27570
rect 9397 27512 9402 27568
rect 9458 27512 9812 27568
rect 9397 27510 9812 27512
rect 9397 27507 9463 27510
rect 9806 27508 9812 27510
rect 9876 27508 9882 27572
rect 25865 27570 25931 27573
rect 26182 27570 26188 27572
rect 25865 27568 26188 27570
rect 25865 27512 25870 27568
rect 25926 27512 26188 27568
rect 25865 27510 26188 27512
rect 25865 27507 25931 27510
rect 26182 27508 26188 27510
rect 26252 27570 26258 27572
rect 26969 27570 27035 27573
rect 26252 27568 27035 27570
rect 26252 27512 26974 27568
rect 27030 27512 27035 27568
rect 26252 27510 27035 27512
rect 27110 27570 27170 27646
rect 27286 27644 27292 27708
rect 27356 27706 27403 27708
rect 27356 27704 27448 27706
rect 27398 27648 27448 27704
rect 27356 27646 27448 27648
rect 27356 27644 27403 27646
rect 27337 27643 27403 27644
rect 28625 27570 28691 27573
rect 27110 27568 28691 27570
rect 27110 27512 28630 27568
rect 28686 27512 28691 27568
rect 27110 27510 28691 27512
rect 26252 27508 26258 27510
rect 26969 27507 27035 27510
rect 28625 27507 28691 27510
rect 30097 27570 30163 27573
rect 30373 27570 30439 27573
rect 31017 27572 31083 27573
rect 30097 27568 30439 27570
rect 30097 27512 30102 27568
rect 30158 27512 30378 27568
rect 30434 27512 30439 27568
rect 30097 27510 30439 27512
rect 30097 27507 30163 27510
rect 30373 27507 30439 27510
rect 30966 27508 30972 27572
rect 31036 27570 31083 27572
rect 31036 27568 31128 27570
rect 31078 27512 31128 27568
rect 31036 27510 31128 27512
rect 31036 27508 31083 27510
rect 31017 27507 31083 27508
rect 26049 27434 26115 27437
rect 27613 27434 27679 27437
rect 26049 27432 27679 27434
rect 26049 27376 26054 27432
rect 26110 27376 27618 27432
rect 27674 27376 27679 27432
rect 26049 27374 27679 27376
rect 26049 27371 26115 27374
rect 27613 27371 27679 27374
rect 5758 27236 5764 27300
rect 5828 27298 5834 27300
rect 5901 27298 5967 27301
rect 5828 27296 5967 27298
rect 5828 27240 5906 27296
rect 5962 27240 5967 27296
rect 5828 27238 5967 27240
rect 5828 27236 5834 27238
rect 5901 27235 5967 27238
rect 7598 27236 7604 27300
rect 7668 27298 7674 27300
rect 8017 27298 8083 27301
rect 7668 27296 8083 27298
rect 7668 27240 8022 27296
rect 8078 27240 8083 27296
rect 7668 27238 8083 27240
rect 7668 27236 7674 27238
rect 8017 27235 8083 27238
rect 12433 27298 12499 27301
rect 26417 27298 26483 27301
rect 27245 27298 27311 27301
rect 12433 27296 27311 27298
rect 12433 27240 12438 27296
rect 12494 27240 26422 27296
rect 26478 27240 27250 27296
rect 27306 27240 27311 27296
rect 12433 27238 27311 27240
rect 12433 27235 12499 27238
rect 26417 27235 26483 27238
rect 27245 27235 27311 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 26877 27162 26943 27165
rect 27153 27162 27219 27165
rect 28257 27162 28323 27165
rect 26877 27160 28323 27162
rect 26877 27104 26882 27160
rect 26938 27104 27158 27160
rect 27214 27104 28262 27160
rect 28318 27104 28323 27160
rect 26877 27102 28323 27104
rect 26877 27099 26943 27102
rect 27153 27099 27219 27102
rect 28257 27099 28323 27102
rect 16389 27026 16455 27029
rect 18597 27026 18663 27029
rect 16389 27024 18663 27026
rect 16389 26968 16394 27024
rect 16450 26968 18602 27024
rect 18658 26968 18663 27024
rect 16389 26966 18663 26968
rect 16389 26963 16455 26966
rect 18597 26963 18663 26966
rect 24485 26890 24551 26893
rect 27153 26890 27219 26893
rect 24485 26888 27219 26890
rect 24485 26832 24490 26888
rect 24546 26832 27158 26888
rect 27214 26832 27219 26888
rect 24485 26830 27219 26832
rect 24485 26827 24551 26830
rect 27153 26827 27219 26830
rect 31518 26828 31524 26892
rect 31588 26890 31594 26892
rect 31661 26890 31727 26893
rect 31588 26888 31727 26890
rect 31588 26832 31666 26888
rect 31722 26832 31727 26888
rect 31588 26830 31727 26832
rect 31588 26828 31594 26830
rect 31661 26827 31727 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 20713 26618 20779 26621
rect 21398 26618 21404 26620
rect 20713 26616 21404 26618
rect 20713 26560 20718 26616
rect 20774 26560 21404 26616
rect 20713 26558 21404 26560
rect 20713 26555 20779 26558
rect 21398 26556 21404 26558
rect 21468 26556 21474 26620
rect 18229 26482 18295 26485
rect 18505 26482 18571 26485
rect 16944 26480 18571 26482
rect 16944 26424 18234 26480
rect 18290 26424 18510 26480
rect 18566 26424 18571 26480
rect 16944 26422 18571 26424
rect 16944 26349 17004 26422
rect 18229 26419 18295 26422
rect 18505 26419 18571 26422
rect 20253 26482 20319 26485
rect 22134 26482 22140 26484
rect 20253 26480 22140 26482
rect 20253 26424 20258 26480
rect 20314 26424 22140 26480
rect 20253 26422 22140 26424
rect 20253 26419 20319 26422
rect 22134 26420 22140 26422
rect 22204 26420 22210 26484
rect 23289 26482 23355 26485
rect 25589 26482 25655 26485
rect 23289 26480 25655 26482
rect 23289 26424 23294 26480
rect 23350 26424 25594 26480
rect 25650 26424 25655 26480
rect 23289 26422 25655 26424
rect 23289 26419 23355 26422
rect 25589 26419 25655 26422
rect 25773 26482 25839 26485
rect 26233 26482 26299 26485
rect 25773 26480 26299 26482
rect 25773 26424 25778 26480
rect 25834 26424 26238 26480
rect 26294 26424 26299 26480
rect 25773 26422 26299 26424
rect 25773 26419 25839 26422
rect 26233 26419 26299 26422
rect 8385 26348 8451 26349
rect 8334 26346 8340 26348
rect 8294 26286 8340 26346
rect 8404 26344 8451 26348
rect 8446 26288 8451 26344
rect 8334 26284 8340 26286
rect 8404 26284 8451 26288
rect 8385 26283 8451 26284
rect 10593 26346 10659 26349
rect 12709 26346 12775 26349
rect 10593 26344 12775 26346
rect 10593 26288 10598 26344
rect 10654 26288 12714 26344
rect 12770 26288 12775 26344
rect 10593 26286 12775 26288
rect 10593 26283 10659 26286
rect 12709 26283 12775 26286
rect 14273 26346 14339 26349
rect 14825 26346 14891 26349
rect 16614 26346 16620 26348
rect 14273 26344 16620 26346
rect 14273 26288 14278 26344
rect 14334 26288 14830 26344
rect 14886 26288 16620 26344
rect 14273 26286 16620 26288
rect 14273 26283 14339 26286
rect 14825 26283 14891 26286
rect 16614 26284 16620 26286
rect 16684 26346 16690 26348
rect 16941 26346 17007 26349
rect 16684 26344 17007 26346
rect 16684 26288 16946 26344
rect 17002 26288 17007 26344
rect 16684 26286 17007 26288
rect 16684 26284 16690 26286
rect 16941 26283 17007 26286
rect 17166 26284 17172 26348
rect 17236 26346 17242 26348
rect 17309 26346 17375 26349
rect 17236 26344 17375 26346
rect 17236 26288 17314 26344
rect 17370 26288 17375 26344
rect 17236 26286 17375 26288
rect 17236 26284 17242 26286
rect 17309 26283 17375 26286
rect 17493 26346 17559 26349
rect 17902 26346 17908 26348
rect 17493 26344 17908 26346
rect 17493 26288 17498 26344
rect 17554 26288 17908 26344
rect 17493 26286 17908 26288
rect 17493 26283 17559 26286
rect 17902 26284 17908 26286
rect 17972 26284 17978 26348
rect 21030 26284 21036 26348
rect 21100 26346 21106 26348
rect 21909 26346 21975 26349
rect 21100 26344 21975 26346
rect 21100 26288 21914 26344
rect 21970 26288 21975 26344
rect 21100 26286 21975 26288
rect 21100 26284 21106 26286
rect 21909 26283 21975 26286
rect 22185 26346 22251 26349
rect 22686 26346 22692 26348
rect 22185 26344 22692 26346
rect 22185 26288 22190 26344
rect 22246 26288 22692 26344
rect 22185 26286 22692 26288
rect 22185 26283 22251 26286
rect 22686 26284 22692 26286
rect 22756 26284 22762 26348
rect 14733 26210 14799 26213
rect 21173 26210 21239 26213
rect 14733 26208 21239 26210
rect 14733 26152 14738 26208
rect 14794 26152 21178 26208
rect 21234 26152 21239 26208
rect 14733 26150 21239 26152
rect 14733 26147 14799 26150
rect 21173 26147 21239 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 16665 26074 16731 26077
rect 17309 26074 17375 26077
rect 16665 26072 17375 26074
rect 16665 26016 16670 26072
rect 16726 26016 17314 26072
rect 17370 26016 17375 26072
rect 16665 26014 17375 26016
rect 16665 26011 16731 26014
rect 17309 26011 17375 26014
rect 11053 25938 11119 25941
rect 12065 25938 12131 25941
rect 12801 25938 12867 25941
rect 32305 25940 32371 25941
rect 11053 25936 12867 25938
rect 11053 25880 11058 25936
rect 11114 25880 12070 25936
rect 12126 25880 12806 25936
rect 12862 25880 12867 25936
rect 11053 25878 12867 25880
rect 11053 25875 11119 25878
rect 12065 25875 12131 25878
rect 12801 25875 12867 25878
rect 32254 25876 32260 25940
rect 32324 25938 32371 25940
rect 32324 25936 32416 25938
rect 32366 25880 32416 25936
rect 32324 25878 32416 25880
rect 32324 25876 32371 25878
rect 32305 25875 32371 25876
rect 23933 25802 23999 25805
rect 24158 25802 24164 25804
rect 23933 25800 24164 25802
rect 23933 25744 23938 25800
rect 23994 25744 24164 25800
rect 23933 25742 24164 25744
rect 23933 25739 23999 25742
rect 24158 25740 24164 25742
rect 24228 25740 24234 25804
rect 7833 25668 7899 25669
rect 29361 25668 29427 25669
rect 7782 25604 7788 25668
rect 7852 25666 7899 25668
rect 7852 25664 7944 25666
rect 7894 25608 7944 25664
rect 7852 25606 7944 25608
rect 7852 25604 7899 25606
rect 29310 25604 29316 25668
rect 29380 25666 29427 25668
rect 30189 25666 30255 25669
rect 29380 25664 30255 25666
rect 29422 25608 30194 25664
rect 30250 25608 30255 25664
rect 29380 25606 30255 25608
rect 29380 25604 29427 25606
rect 7833 25603 7899 25604
rect 29361 25603 29427 25604
rect 30189 25603 30255 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 10225 25530 10291 25533
rect 11145 25530 11211 25533
rect 10225 25528 11211 25530
rect 10225 25472 10230 25528
rect 10286 25472 11150 25528
rect 11206 25472 11211 25528
rect 10225 25470 11211 25472
rect 10225 25467 10291 25470
rect 11145 25467 11211 25470
rect 32029 25530 32095 25533
rect 32765 25530 32831 25533
rect 32029 25528 32831 25530
rect 32029 25472 32034 25528
rect 32090 25472 32770 25528
rect 32826 25472 32831 25528
rect 32029 25470 32831 25472
rect 32029 25467 32095 25470
rect 32765 25467 32831 25470
rect 22001 25394 22067 25397
rect 25405 25394 25471 25397
rect 22001 25392 25471 25394
rect 22001 25336 22006 25392
rect 22062 25336 25410 25392
rect 25466 25336 25471 25392
rect 22001 25334 25471 25336
rect 22001 25331 22067 25334
rect 25405 25331 25471 25334
rect 32213 25394 32279 25397
rect 32213 25392 32322 25394
rect 32213 25336 32218 25392
rect 32274 25336 32322 25392
rect 32213 25331 32322 25336
rect 5717 25256 5783 25261
rect 5717 25200 5722 25256
rect 5778 25200 5783 25256
rect 5717 25195 5783 25200
rect 20529 25258 20595 25261
rect 21357 25258 21423 25261
rect 20529 25256 21423 25258
rect 20529 25200 20534 25256
rect 20590 25200 21362 25256
rect 21418 25200 21423 25256
rect 20529 25198 21423 25200
rect 20529 25195 20595 25198
rect 21357 25195 21423 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 5720 24986 5780 25195
rect 32262 25125 32322 25331
rect 5942 25060 5948 25124
rect 6012 25122 6018 25124
rect 6085 25122 6151 25125
rect 6012 25120 6151 25122
rect 6012 25064 6090 25120
rect 6146 25064 6151 25120
rect 6012 25062 6151 25064
rect 6012 25060 6018 25062
rect 6085 25059 6151 25062
rect 11053 25122 11119 25125
rect 12157 25122 12223 25125
rect 11053 25120 12223 25122
rect 11053 25064 11058 25120
rect 11114 25064 12162 25120
rect 12218 25064 12223 25120
rect 11053 25062 12223 25064
rect 11053 25059 11119 25062
rect 12157 25059 12223 25062
rect 32213 25120 32322 25125
rect 32213 25064 32218 25120
rect 32274 25064 32322 25120
rect 32213 25062 32322 25064
rect 32213 25059 32279 25062
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 6085 24986 6151 24989
rect 5720 24984 6151 24986
rect 5720 24928 6090 24984
rect 6146 24928 6151 24984
rect 5720 24926 6151 24928
rect 6085 24923 6151 24926
rect 10869 24986 10935 24989
rect 12341 24986 12407 24989
rect 10869 24984 12407 24986
rect 10869 24928 10874 24984
rect 10930 24928 12346 24984
rect 12402 24928 12407 24984
rect 10869 24926 12407 24928
rect 10869 24923 10935 24926
rect 12341 24923 12407 24926
rect 18270 24924 18276 24988
rect 18340 24986 18346 24988
rect 20529 24986 20595 24989
rect 18340 24984 20595 24986
rect 18340 24928 20534 24984
rect 20590 24928 20595 24984
rect 18340 24926 20595 24928
rect 18340 24924 18346 24926
rect 20529 24923 20595 24926
rect 30005 24986 30071 24989
rect 31293 24986 31359 24989
rect 33961 24986 34027 24989
rect 30005 24984 34027 24986
rect 30005 24928 30010 24984
rect 30066 24928 31298 24984
rect 31354 24928 33966 24984
rect 34022 24928 34027 24984
rect 30005 24926 34027 24928
rect 30005 24923 30071 24926
rect 31293 24923 31359 24926
rect 33961 24923 34027 24926
rect 3141 24850 3207 24853
rect 8845 24850 8911 24853
rect 3141 24848 8911 24850
rect 3141 24792 3146 24848
rect 3202 24792 8850 24848
rect 8906 24792 8911 24848
rect 3141 24790 8911 24792
rect 3141 24787 3207 24790
rect 8845 24787 8911 24790
rect 12249 24850 12315 24853
rect 14038 24850 14044 24852
rect 12249 24848 14044 24850
rect 12249 24792 12254 24848
rect 12310 24792 14044 24848
rect 12249 24790 14044 24792
rect 12249 24787 12315 24790
rect 14038 24788 14044 24790
rect 14108 24788 14114 24852
rect 15101 24850 15167 24853
rect 16573 24850 16639 24853
rect 15101 24848 16639 24850
rect 15101 24792 15106 24848
rect 15162 24792 16578 24848
rect 16634 24792 16639 24848
rect 15101 24790 16639 24792
rect 15101 24787 15167 24790
rect 16573 24787 16639 24790
rect 24393 24850 24459 24853
rect 25865 24850 25931 24853
rect 24393 24848 25931 24850
rect 24393 24792 24398 24848
rect 24454 24792 25870 24848
rect 25926 24792 25931 24848
rect 24393 24790 25931 24792
rect 24393 24787 24459 24790
rect 25865 24787 25931 24790
rect 28809 24850 28875 24853
rect 28809 24848 29010 24850
rect 28809 24792 28814 24848
rect 28870 24792 29010 24848
rect 28809 24790 29010 24792
rect 28809 24787 28875 24790
rect 8753 24714 8819 24717
rect 12709 24714 12775 24717
rect 12893 24714 12959 24717
rect 8753 24712 12959 24714
rect 8753 24656 8758 24712
rect 8814 24656 12714 24712
rect 12770 24656 12898 24712
rect 12954 24656 12959 24712
rect 8753 24654 12959 24656
rect 8753 24651 8819 24654
rect 12709 24651 12775 24654
rect 12893 24651 12959 24654
rect 16665 24714 16731 24717
rect 16941 24714 17007 24717
rect 16665 24712 17007 24714
rect 16665 24656 16670 24712
rect 16726 24656 16946 24712
rect 17002 24656 17007 24712
rect 16665 24654 17007 24656
rect 16665 24651 16731 24654
rect 16941 24651 17007 24654
rect 27153 24714 27219 24717
rect 28717 24714 28783 24717
rect 27153 24712 28783 24714
rect 27153 24656 27158 24712
rect 27214 24656 28722 24712
rect 28778 24656 28783 24712
rect 27153 24654 28783 24656
rect 27153 24651 27219 24654
rect 28717 24651 28783 24654
rect 10501 24578 10567 24581
rect 12750 24578 12756 24580
rect 10501 24576 12756 24578
rect 10501 24520 10506 24576
rect 10562 24520 12756 24576
rect 10501 24518 12756 24520
rect 10501 24515 10567 24518
rect 12750 24516 12756 24518
rect 12820 24516 12826 24580
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 12525 24442 12591 24445
rect 12934 24442 12940 24444
rect 12525 24440 12940 24442
rect 12525 24384 12530 24440
rect 12586 24384 12940 24440
rect 12525 24382 12940 24384
rect 12525 24379 12591 24382
rect 12934 24380 12940 24382
rect 13004 24380 13010 24444
rect 16798 24380 16804 24444
rect 16868 24442 16874 24444
rect 16941 24442 17007 24445
rect 16868 24440 17007 24442
rect 16868 24384 16946 24440
rect 17002 24384 17007 24440
rect 16868 24382 17007 24384
rect 16868 24380 16874 24382
rect 16941 24379 17007 24382
rect 28717 24442 28783 24445
rect 28950 24442 29010 24790
rect 35985 24578 36051 24581
rect 36782 24578 37582 24608
rect 35985 24576 37582 24578
rect 35985 24520 35990 24576
rect 36046 24520 37582 24576
rect 35985 24518 37582 24520
rect 35985 24515 36051 24518
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 36782 24488 37582 24518
rect 34930 24447 35246 24448
rect 28717 24440 29010 24442
rect 28717 24384 28722 24440
rect 28778 24384 29010 24440
rect 28717 24382 29010 24384
rect 28717 24379 28783 24382
rect 5441 24306 5507 24309
rect 9765 24306 9831 24309
rect 13077 24308 13143 24309
rect 11094 24306 11100 24308
rect 5441 24304 9690 24306
rect 5441 24248 5446 24304
rect 5502 24248 9690 24304
rect 5441 24246 9690 24248
rect 5441 24243 5507 24246
rect 4061 24170 4127 24173
rect 7373 24170 7439 24173
rect 4061 24168 7439 24170
rect 4061 24112 4066 24168
rect 4122 24112 7378 24168
rect 7434 24112 7439 24168
rect 4061 24110 7439 24112
rect 9630 24170 9690 24246
rect 9765 24304 11100 24306
rect 9765 24248 9770 24304
rect 9826 24248 11100 24304
rect 9765 24246 11100 24248
rect 9765 24243 9831 24246
rect 11094 24244 11100 24246
rect 11164 24244 11170 24308
rect 13077 24306 13124 24308
rect 13032 24304 13124 24306
rect 13032 24248 13082 24304
rect 13032 24246 13124 24248
rect 13077 24244 13124 24246
rect 13188 24244 13194 24308
rect 30925 24306 30991 24309
rect 31477 24306 31543 24309
rect 30925 24304 31543 24306
rect 30925 24248 30930 24304
rect 30986 24248 31482 24304
rect 31538 24248 31543 24304
rect 30925 24246 31543 24248
rect 13077 24243 13143 24244
rect 30925 24243 30991 24246
rect 31477 24243 31543 24246
rect 10409 24170 10475 24173
rect 9630 24168 10475 24170
rect 9630 24112 10414 24168
rect 10470 24112 10475 24168
rect 9630 24110 10475 24112
rect 4061 24107 4127 24110
rect 7373 24107 7439 24110
rect 10409 24107 10475 24110
rect 16297 24170 16363 24173
rect 19241 24170 19307 24173
rect 20805 24172 20871 24173
rect 27521 24172 27587 24173
rect 20805 24170 20852 24172
rect 16297 24168 19307 24170
rect 16297 24112 16302 24168
rect 16358 24112 19246 24168
rect 19302 24112 19307 24168
rect 16297 24110 19307 24112
rect 20760 24168 20852 24170
rect 20760 24112 20810 24168
rect 20760 24110 20852 24112
rect 16297 24107 16363 24110
rect 19241 24107 19307 24110
rect 20805 24108 20852 24110
rect 20916 24108 20922 24172
rect 27470 24170 27476 24172
rect 27430 24110 27476 24170
rect 27540 24168 27587 24172
rect 27582 24112 27587 24168
rect 27470 24108 27476 24110
rect 27540 24108 27587 24112
rect 20805 24107 20871 24108
rect 27521 24107 27587 24108
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 19609 23898 19675 23901
rect 23606 23898 23612 23900
rect 19609 23896 23612 23898
rect 19609 23840 19614 23896
rect 19670 23840 23612 23896
rect 19609 23838 23612 23840
rect 19609 23835 19675 23838
rect 23606 23836 23612 23838
rect 23676 23836 23682 23900
rect 36077 23898 36143 23901
rect 36782 23898 37582 23928
rect 36077 23896 37582 23898
rect 36077 23840 36082 23896
rect 36138 23840 37582 23896
rect 36077 23838 37582 23840
rect 36077 23835 36143 23838
rect 36782 23808 37582 23838
rect 5349 23762 5415 23765
rect 6545 23762 6611 23765
rect 7373 23762 7439 23765
rect 5349 23760 7439 23762
rect 5349 23704 5354 23760
rect 5410 23704 6550 23760
rect 6606 23704 7378 23760
rect 7434 23704 7439 23760
rect 5349 23702 7439 23704
rect 5349 23699 5415 23702
rect 6545 23699 6611 23702
rect 7373 23699 7439 23702
rect 14590 23700 14596 23764
rect 14660 23762 14666 23764
rect 15653 23762 15719 23765
rect 14660 23760 15719 23762
rect 14660 23704 15658 23760
rect 15714 23704 15719 23760
rect 14660 23702 15719 23704
rect 14660 23700 14666 23702
rect 15653 23699 15719 23702
rect 21214 23700 21220 23764
rect 21284 23762 21290 23764
rect 22645 23762 22711 23765
rect 21284 23760 22711 23762
rect 21284 23704 22650 23760
rect 22706 23704 22711 23760
rect 21284 23702 22711 23704
rect 21284 23700 21290 23702
rect 22645 23699 22711 23702
rect 30782 23700 30788 23764
rect 30852 23762 30858 23764
rect 31293 23762 31359 23765
rect 30852 23760 31359 23762
rect 30852 23704 31298 23760
rect 31354 23704 31359 23760
rect 30852 23702 31359 23704
rect 30852 23700 30858 23702
rect 31293 23699 31359 23702
rect 2865 23626 2931 23629
rect 5901 23626 5967 23629
rect 2865 23624 5967 23626
rect 2865 23568 2870 23624
rect 2926 23568 5906 23624
rect 5962 23568 5967 23624
rect 2865 23566 5967 23568
rect 2865 23563 2931 23566
rect 5901 23563 5967 23566
rect 6085 23626 6151 23629
rect 9765 23626 9831 23629
rect 6085 23624 9831 23626
rect 6085 23568 6090 23624
rect 6146 23568 9770 23624
rect 9826 23568 9831 23624
rect 6085 23566 9831 23568
rect 6085 23563 6151 23566
rect 9765 23563 9831 23566
rect 11329 23626 11395 23629
rect 11462 23626 11468 23628
rect 11329 23624 11468 23626
rect 11329 23568 11334 23624
rect 11390 23568 11468 23624
rect 11329 23566 11468 23568
rect 11329 23563 11395 23566
rect 11462 23564 11468 23566
rect 11532 23564 11538 23628
rect 13721 23626 13787 23629
rect 14222 23626 14228 23628
rect 13721 23624 14228 23626
rect 13721 23568 13726 23624
rect 13782 23568 14228 23624
rect 13721 23566 14228 23568
rect 13721 23563 13787 23566
rect 14222 23564 14228 23566
rect 14292 23626 14298 23628
rect 15469 23626 15535 23629
rect 14292 23624 15535 23626
rect 14292 23568 15474 23624
rect 15530 23568 15535 23624
rect 14292 23566 15535 23568
rect 14292 23564 14298 23566
rect 15469 23563 15535 23566
rect 5073 23490 5139 23493
rect 7373 23490 7439 23493
rect 5073 23488 7439 23490
rect 5073 23432 5078 23488
rect 5134 23432 7378 23488
rect 7434 23432 7439 23488
rect 5073 23430 7439 23432
rect 5073 23427 5139 23430
rect 7373 23427 7439 23430
rect 9581 23492 9647 23493
rect 9581 23488 9628 23492
rect 9692 23490 9698 23492
rect 13261 23490 13327 23493
rect 13486 23490 13492 23492
rect 9581 23432 9586 23488
rect 9581 23428 9628 23432
rect 9692 23430 9738 23490
rect 13261 23488 13492 23490
rect 13261 23432 13266 23488
rect 13322 23432 13492 23488
rect 13261 23430 13492 23432
rect 9692 23428 9698 23430
rect 9581 23427 9647 23428
rect 13261 23427 13327 23430
rect 13486 23428 13492 23430
rect 13556 23428 13562 23492
rect 13997 23490 14063 23493
rect 17401 23490 17467 23493
rect 13997 23488 17467 23490
rect 13997 23432 14002 23488
rect 14058 23432 17406 23488
rect 17462 23432 17467 23488
rect 13997 23430 17467 23432
rect 13997 23427 14063 23430
rect 17401 23427 17467 23430
rect 17769 23490 17835 23493
rect 19885 23490 19951 23493
rect 17769 23488 19951 23490
rect 17769 23432 17774 23488
rect 17830 23432 19890 23488
rect 19946 23432 19951 23488
rect 17769 23430 19951 23432
rect 17769 23427 17835 23430
rect 19885 23427 19951 23430
rect 25405 23490 25471 23493
rect 28809 23490 28875 23493
rect 25405 23488 28875 23490
rect 25405 23432 25410 23488
rect 25466 23432 28814 23488
rect 28870 23432 28875 23488
rect 25405 23430 28875 23432
rect 25405 23427 25471 23430
rect 28809 23427 28875 23430
rect 30925 23490 30991 23493
rect 31150 23490 31156 23492
rect 30925 23488 31156 23490
rect 30925 23432 30930 23488
rect 30986 23432 31156 23488
rect 30925 23430 31156 23432
rect 30925 23427 30991 23430
rect 31150 23428 31156 23430
rect 31220 23428 31226 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 5165 23354 5231 23357
rect 6637 23354 6703 23357
rect 8109 23354 8175 23357
rect 9397 23354 9463 23357
rect 5165 23352 9463 23354
rect 5165 23296 5170 23352
rect 5226 23296 6642 23352
rect 6698 23296 8114 23352
rect 8170 23296 9402 23352
rect 9458 23296 9463 23352
rect 5165 23294 9463 23296
rect 5165 23291 5231 23294
rect 6637 23291 6703 23294
rect 8109 23291 8175 23294
rect 9397 23291 9463 23294
rect 11973 23354 12039 23357
rect 15285 23354 15351 23357
rect 17033 23356 17099 23357
rect 11973 23352 15351 23354
rect 11973 23296 11978 23352
rect 12034 23296 15290 23352
rect 15346 23296 15351 23352
rect 11973 23294 15351 23296
rect 11973 23291 12039 23294
rect 15285 23291 15351 23294
rect 16982 23292 16988 23356
rect 17052 23354 17099 23356
rect 17861 23354 17927 23357
rect 19333 23354 19399 23357
rect 17052 23352 17144 23354
rect 17094 23296 17144 23352
rect 17052 23294 17144 23296
rect 17861 23352 19399 23354
rect 17861 23296 17866 23352
rect 17922 23296 19338 23352
rect 19394 23296 19399 23352
rect 17861 23294 19399 23296
rect 17052 23292 17099 23294
rect 17033 23291 17099 23292
rect 17861 23291 17927 23294
rect 19333 23291 19399 23294
rect 5257 23218 5323 23221
rect 8385 23218 8451 23221
rect 9581 23218 9647 23221
rect 5257 23216 9647 23218
rect 5257 23160 5262 23216
rect 5318 23160 8390 23216
rect 8446 23160 9586 23216
rect 9642 23160 9647 23216
rect 5257 23158 9647 23160
rect 5257 23155 5323 23158
rect 8385 23155 8451 23158
rect 9581 23155 9647 23158
rect 12617 23218 12683 23221
rect 13629 23218 13695 23221
rect 12617 23216 13695 23218
rect 12617 23160 12622 23216
rect 12678 23160 13634 23216
rect 13690 23160 13695 23216
rect 12617 23158 13695 23160
rect 12617 23155 12683 23158
rect 13629 23155 13695 23158
rect 14733 23218 14799 23221
rect 18137 23218 18203 23221
rect 14733 23216 18203 23218
rect 14733 23160 14738 23216
rect 14794 23160 18142 23216
rect 18198 23160 18203 23216
rect 14733 23158 18203 23160
rect 14733 23155 14799 23158
rect 18137 23155 18203 23158
rect 19057 23218 19123 23221
rect 19977 23218 20043 23221
rect 19057 23216 20043 23218
rect 19057 23160 19062 23216
rect 19118 23160 19982 23216
rect 20038 23160 20043 23216
rect 19057 23158 20043 23160
rect 19057 23155 19123 23158
rect 19977 23155 20043 23158
rect 2630 23020 2636 23084
rect 2700 23082 2706 23084
rect 7189 23082 7255 23085
rect 2700 23080 7255 23082
rect 2700 23024 7194 23080
rect 7250 23024 7255 23080
rect 2700 23022 7255 23024
rect 2700 23020 2706 23022
rect 7189 23019 7255 23022
rect 11053 23082 11119 23085
rect 11605 23082 11671 23085
rect 11881 23082 11947 23085
rect 11053 23080 11947 23082
rect 11053 23024 11058 23080
rect 11114 23024 11610 23080
rect 11666 23024 11886 23080
rect 11942 23024 11947 23080
rect 11053 23022 11947 23024
rect 11053 23019 11119 23022
rect 11605 23019 11671 23022
rect 11881 23019 11947 23022
rect 12341 23082 12407 23085
rect 16297 23082 16363 23085
rect 12341 23080 16363 23082
rect 12341 23024 12346 23080
rect 12402 23024 16302 23080
rect 16358 23024 16363 23080
rect 12341 23022 16363 23024
rect 12341 23019 12407 23022
rect 16297 23019 16363 23022
rect 16798 23020 16804 23084
rect 16868 23082 16874 23084
rect 16941 23082 17007 23085
rect 18781 23082 18847 23085
rect 18965 23082 19031 23085
rect 16868 23080 19031 23082
rect 16868 23024 16946 23080
rect 17002 23024 18786 23080
rect 18842 23024 18970 23080
rect 19026 23024 19031 23080
rect 16868 23022 19031 23024
rect 16868 23020 16874 23022
rect 16941 23019 17007 23022
rect 18781 23019 18847 23022
rect 18965 23019 19031 23022
rect 3918 22884 3924 22948
rect 3988 22946 3994 22948
rect 4245 22946 4311 22949
rect 6361 22948 6427 22949
rect 6310 22946 6316 22948
rect 3988 22944 4311 22946
rect 3988 22888 4250 22944
rect 4306 22888 4311 22944
rect 3988 22886 4311 22888
rect 6270 22886 6316 22946
rect 6380 22944 6427 22948
rect 6422 22888 6427 22944
rect 3988 22884 3994 22886
rect 4245 22883 4311 22886
rect 6310 22884 6316 22886
rect 6380 22884 6427 22888
rect 6361 22883 6427 22884
rect 14365 22946 14431 22949
rect 14825 22946 14891 22949
rect 14365 22944 14891 22946
rect 14365 22888 14370 22944
rect 14426 22888 14830 22944
rect 14886 22888 14891 22944
rect 14365 22886 14891 22888
rect 14365 22883 14431 22886
rect 14825 22883 14891 22886
rect 17033 22946 17099 22949
rect 19149 22946 19215 22949
rect 17033 22944 19215 22946
rect 17033 22888 17038 22944
rect 17094 22888 19154 22944
rect 19210 22888 19215 22944
rect 17033 22886 19215 22888
rect 17033 22883 17099 22886
rect 19149 22883 19215 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 4429 22810 4495 22813
rect 5809 22810 5875 22813
rect 6085 22810 6151 22813
rect 7649 22810 7715 22813
rect 4429 22808 4722 22810
rect 4429 22752 4434 22808
rect 4490 22752 4722 22808
rect 4429 22750 4722 22752
rect 4429 22747 4495 22750
rect 4662 22674 4722 22750
rect 5809 22808 6010 22810
rect 5809 22752 5814 22808
rect 5870 22752 6010 22808
rect 5809 22750 6010 22752
rect 5809 22747 5875 22750
rect 5950 22677 6010 22750
rect 6085 22808 7715 22810
rect 6085 22752 6090 22808
rect 6146 22752 7654 22808
rect 7710 22752 7715 22808
rect 6085 22750 7715 22752
rect 6085 22747 6151 22750
rect 7649 22747 7715 22750
rect 19190 22748 19196 22812
rect 19260 22810 19266 22812
rect 29494 22810 29500 22812
rect 19260 22750 29500 22810
rect 19260 22748 19266 22750
rect 29494 22748 29500 22750
rect 29564 22748 29570 22812
rect 4889 22674 4955 22677
rect 4662 22672 4955 22674
rect 4662 22616 4894 22672
rect 4950 22616 4955 22672
rect 4662 22614 4955 22616
rect 4889 22611 4955 22614
rect 5625 22674 5691 22677
rect 5809 22674 5875 22677
rect 5625 22672 5875 22674
rect 5625 22616 5630 22672
rect 5686 22616 5814 22672
rect 5870 22616 5875 22672
rect 5625 22614 5875 22616
rect 5950 22674 6059 22677
rect 6637 22674 6703 22677
rect 9029 22674 9095 22677
rect 5950 22672 9095 22674
rect 5950 22616 5998 22672
rect 6054 22616 6642 22672
rect 6698 22616 9034 22672
rect 9090 22616 9095 22672
rect 5950 22614 9095 22616
rect 5625 22611 5691 22614
rect 5809 22611 5875 22614
rect 5993 22611 6059 22614
rect 6637 22611 6703 22614
rect 9029 22611 9095 22614
rect 10501 22674 10567 22677
rect 12157 22674 12223 22677
rect 10501 22672 12223 22674
rect 10501 22616 10506 22672
rect 10562 22616 12162 22672
rect 12218 22616 12223 22672
rect 10501 22614 12223 22616
rect 10501 22611 10567 22614
rect 12157 22611 12223 22614
rect 13445 22674 13511 22677
rect 18229 22674 18295 22677
rect 13445 22672 18295 22674
rect 13445 22616 13450 22672
rect 13506 22616 18234 22672
rect 18290 22616 18295 22672
rect 13445 22614 18295 22616
rect 13445 22611 13511 22614
rect 18229 22611 18295 22614
rect 25405 22676 25471 22677
rect 25405 22672 25452 22676
rect 25516 22674 25522 22676
rect 25405 22616 25410 22672
rect 25405 22612 25452 22616
rect 25516 22614 25562 22674
rect 25516 22612 25522 22614
rect 25405 22611 25471 22612
rect 5165 22538 5231 22541
rect 5533 22538 5599 22541
rect 9121 22540 9187 22541
rect 5165 22536 5599 22538
rect 5165 22480 5170 22536
rect 5226 22480 5538 22536
rect 5594 22480 5599 22536
rect 5165 22478 5599 22480
rect 5165 22475 5231 22478
rect 5533 22475 5599 22478
rect 9070 22476 9076 22540
rect 9140 22538 9187 22540
rect 10593 22538 10659 22541
rect 11605 22538 11671 22541
rect 9140 22536 9232 22538
rect 9182 22480 9232 22536
rect 9140 22478 9232 22480
rect 10593 22536 11671 22538
rect 10593 22480 10598 22536
rect 10654 22480 11610 22536
rect 11666 22480 11671 22536
rect 10593 22478 11671 22480
rect 9140 22476 9187 22478
rect 9121 22475 9187 22476
rect 10593 22475 10659 22478
rect 11605 22475 11671 22478
rect 14641 22538 14707 22541
rect 15837 22538 15903 22541
rect 14641 22536 15903 22538
rect 14641 22480 14646 22536
rect 14702 22480 15842 22536
rect 15898 22480 15903 22536
rect 14641 22478 15903 22480
rect 14641 22475 14707 22478
rect 15837 22475 15903 22478
rect 21582 22476 21588 22540
rect 21652 22538 21658 22540
rect 22001 22538 22067 22541
rect 21652 22536 22067 22538
rect 21652 22480 22006 22536
rect 22062 22480 22067 22536
rect 21652 22478 22067 22480
rect 21652 22476 21658 22478
rect 22001 22475 22067 22478
rect 28165 22540 28231 22541
rect 28165 22536 28212 22540
rect 28276 22538 28282 22540
rect 36077 22538 36143 22541
rect 36782 22538 37582 22568
rect 28165 22480 28170 22536
rect 28165 22476 28212 22480
rect 28276 22478 28322 22538
rect 36077 22536 37582 22538
rect 36077 22480 36082 22536
rect 36138 22480 37582 22536
rect 36077 22478 37582 22480
rect 28276 22476 28282 22478
rect 28165 22475 28231 22476
rect 36077 22475 36143 22478
rect 36782 22448 37582 22478
rect 8109 22404 8175 22405
rect 8109 22400 8156 22404
rect 8220 22402 8226 22404
rect 11789 22402 11855 22405
rect 15377 22402 15443 22405
rect 15653 22402 15719 22405
rect 24393 22404 24459 22405
rect 24342 22402 24348 22404
rect 8109 22344 8114 22400
rect 8109 22340 8156 22344
rect 8220 22342 8266 22402
rect 11789 22400 11898 22402
rect 11789 22344 11794 22400
rect 11850 22344 11898 22400
rect 8220 22340 8226 22342
rect 8109 22339 8175 22340
rect 11789 22339 11898 22344
rect 15377 22400 15719 22402
rect 15377 22344 15382 22400
rect 15438 22344 15658 22400
rect 15714 22344 15719 22400
rect 15377 22342 15719 22344
rect 24302 22342 24348 22402
rect 24412 22400 24459 22404
rect 24454 22344 24459 22400
rect 15377 22339 15443 22342
rect 15653 22339 15719 22342
rect 24342 22340 24348 22342
rect 24412 22340 24459 22344
rect 24894 22340 24900 22404
rect 24964 22402 24970 22404
rect 25589 22402 25655 22405
rect 24964 22400 25655 22402
rect 24964 22344 25594 22400
rect 25650 22344 25655 22400
rect 24964 22342 25655 22344
rect 24964 22340 24970 22342
rect 24393 22339 24459 22340
rect 25589 22339 25655 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 9673 22266 9739 22269
rect 10041 22266 10107 22269
rect 9673 22264 10107 22266
rect 9673 22208 9678 22264
rect 9734 22208 10046 22264
rect 10102 22208 10107 22264
rect 9673 22206 10107 22208
rect 11838 22266 11898 22339
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 12065 22266 12131 22269
rect 11838 22264 12131 22266
rect 11838 22208 12070 22264
rect 12126 22208 12131 22264
rect 11838 22206 12131 22208
rect 9673 22203 9739 22206
rect 10041 22203 10107 22206
rect 12065 22203 12131 22206
rect 28993 22266 29059 22269
rect 32806 22266 32812 22268
rect 28993 22264 32812 22266
rect 28993 22208 28998 22264
rect 29054 22208 32812 22264
rect 28993 22206 32812 22208
rect 28993 22203 29059 22206
rect 32806 22204 32812 22206
rect 32876 22204 32882 22268
rect 8661 22130 8727 22133
rect 8526 22128 8727 22130
rect 8526 22072 8666 22128
rect 8722 22072 8727 22128
rect 8526 22070 8727 22072
rect 8526 21997 8586 22070
rect 8661 22067 8727 22070
rect 11278 22068 11284 22132
rect 11348 22130 11354 22132
rect 13854 22130 13860 22132
rect 11348 22070 13860 22130
rect 11348 22068 11354 22070
rect 13854 22068 13860 22070
rect 13924 22068 13930 22132
rect 15377 22130 15443 22133
rect 16573 22130 16639 22133
rect 17677 22130 17743 22133
rect 15377 22128 17743 22130
rect 15377 22072 15382 22128
rect 15438 22072 16578 22128
rect 16634 22072 17682 22128
rect 17738 22072 17743 22128
rect 15377 22070 17743 22072
rect 15377 22067 15443 22070
rect 16573 22067 16639 22070
rect 17677 22067 17743 22070
rect 18505 22130 18571 22133
rect 19609 22130 19675 22133
rect 23013 22132 23079 22133
rect 23013 22130 23060 22132
rect 18505 22128 19675 22130
rect 18505 22072 18510 22128
rect 18566 22072 19614 22128
rect 19670 22072 19675 22128
rect 18505 22070 19675 22072
rect 22968 22128 23060 22130
rect 22968 22072 23018 22128
rect 22968 22070 23060 22072
rect 18505 22067 18571 22070
rect 19609 22067 19675 22070
rect 23013 22068 23060 22070
rect 23124 22068 23130 22132
rect 31293 22130 31359 22133
rect 32438 22130 32444 22132
rect 31293 22128 32444 22130
rect 31293 22072 31298 22128
rect 31354 22072 32444 22128
rect 31293 22070 32444 22072
rect 23013 22067 23079 22068
rect 31293 22067 31359 22070
rect 32438 22068 32444 22070
rect 32508 22068 32514 22132
rect 6678 21932 6684 21996
rect 6748 21994 6754 21996
rect 7465 21994 7531 21997
rect 6748 21992 7531 21994
rect 6748 21936 7470 21992
rect 7526 21936 7531 21992
rect 6748 21934 7531 21936
rect 6748 21932 6754 21934
rect 7465 21931 7531 21934
rect 8477 21992 8586 21997
rect 8477 21936 8482 21992
rect 8538 21936 8586 21992
rect 8477 21934 8586 21936
rect 8477 21931 8543 21934
rect 10910 21932 10916 21996
rect 10980 21994 10986 21996
rect 12198 21994 12204 21996
rect 10980 21934 12204 21994
rect 10980 21932 10986 21934
rect 12198 21932 12204 21934
rect 12268 21994 12274 21996
rect 12341 21994 12407 21997
rect 12268 21992 12407 21994
rect 12268 21936 12346 21992
rect 12402 21936 12407 21992
rect 12268 21934 12407 21936
rect 12268 21932 12274 21934
rect 12341 21931 12407 21934
rect 15745 21994 15811 21997
rect 16757 21994 16823 21997
rect 17769 21994 17835 21997
rect 15745 21992 17835 21994
rect 15745 21936 15750 21992
rect 15806 21936 16762 21992
rect 16818 21936 17774 21992
rect 17830 21936 17835 21992
rect 15745 21934 17835 21936
rect 15745 21931 15811 21934
rect 16757 21931 16823 21934
rect 17769 21931 17835 21934
rect 19333 21994 19399 21997
rect 20294 21994 20300 21996
rect 19333 21992 20300 21994
rect 19333 21936 19338 21992
rect 19394 21936 20300 21992
rect 19333 21934 20300 21936
rect 19333 21931 19399 21934
rect 20294 21932 20300 21934
rect 20364 21932 20370 21996
rect 26233 21994 26299 21997
rect 26366 21994 26372 21996
rect 26233 21992 26372 21994
rect 26233 21936 26238 21992
rect 26294 21936 26372 21992
rect 26233 21934 26372 21936
rect 20302 21861 20362 21932
rect 26233 21931 26299 21934
rect 26366 21932 26372 21934
rect 26436 21932 26442 21996
rect 10593 21858 10659 21861
rect 16389 21858 16455 21861
rect 10593 21856 16455 21858
rect 10593 21800 10598 21856
rect 10654 21800 16394 21856
rect 16450 21800 16455 21856
rect 10593 21798 16455 21800
rect 10593 21795 10659 21798
rect 16389 21795 16455 21798
rect 20253 21856 20362 21861
rect 20253 21800 20258 21856
rect 20314 21800 20362 21856
rect 20253 21798 20362 21800
rect 36077 21858 36143 21861
rect 36782 21858 37582 21888
rect 36077 21856 37582 21858
rect 36077 21800 36082 21856
rect 36138 21800 37582 21856
rect 36077 21798 37582 21800
rect 20253 21795 20319 21798
rect 36077 21795 36143 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 36782 21768 37582 21798
rect 35590 21727 35906 21728
rect 15377 21586 15443 21589
rect 15510 21586 15516 21588
rect 15377 21584 15516 21586
rect 15377 21528 15382 21584
rect 15438 21528 15516 21584
rect 15377 21526 15516 21528
rect 15377 21523 15443 21526
rect 15510 21524 15516 21526
rect 15580 21524 15586 21588
rect 15009 21450 15075 21453
rect 19241 21450 19307 21453
rect 15009 21448 19307 21450
rect 15009 21392 15014 21448
rect 15070 21392 19246 21448
rect 19302 21392 19307 21448
rect 15009 21390 19307 21392
rect 15009 21387 15075 21390
rect 19241 21387 19307 21390
rect 35249 21450 35315 21453
rect 35801 21450 35867 21453
rect 35249 21448 35867 21450
rect 35249 21392 35254 21448
rect 35310 21392 35806 21448
rect 35862 21392 35867 21448
rect 35249 21390 35867 21392
rect 35249 21387 35315 21390
rect 35801 21387 35867 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 12249 21178 12315 21181
rect 12985 21178 13051 21181
rect 13302 21178 13308 21180
rect 12249 21176 13308 21178
rect 12249 21120 12254 21176
rect 12310 21120 12990 21176
rect 13046 21120 13308 21176
rect 12249 21118 13308 21120
rect 12249 21115 12315 21118
rect 12985 21115 13051 21118
rect 13302 21116 13308 21118
rect 13372 21116 13378 21180
rect 36077 21178 36143 21181
rect 36782 21178 37582 21208
rect 36077 21176 37582 21178
rect 36077 21120 36082 21176
rect 36138 21120 37582 21176
rect 36077 21118 37582 21120
rect 36077 21115 36143 21118
rect 36782 21088 37582 21118
rect 21357 21042 21423 21045
rect 25313 21042 25379 21045
rect 21357 21040 25379 21042
rect 21357 20984 21362 21040
rect 21418 20984 25318 21040
rect 25374 20984 25379 21040
rect 21357 20982 25379 20984
rect 21357 20979 21423 20982
rect 25313 20979 25379 20982
rect 4613 20906 4679 20909
rect 5390 20906 5396 20908
rect 4613 20904 5396 20906
rect 4613 20848 4618 20904
rect 4674 20848 5396 20904
rect 4613 20846 5396 20848
rect 4613 20843 4679 20846
rect 5390 20844 5396 20846
rect 5460 20844 5466 20908
rect 5625 20906 5691 20909
rect 7833 20906 7899 20909
rect 5625 20904 7899 20906
rect 5625 20848 5630 20904
rect 5686 20848 7838 20904
rect 7894 20848 7899 20904
rect 5625 20846 7899 20848
rect 5625 20843 5691 20846
rect 7833 20843 7899 20846
rect 15326 20844 15332 20908
rect 15396 20906 15402 20908
rect 17033 20906 17099 20909
rect 35801 20906 35867 20909
rect 15396 20904 35867 20906
rect 15396 20848 17038 20904
rect 17094 20848 35806 20904
rect 35862 20848 35867 20904
rect 15396 20846 35867 20848
rect 15396 20844 15402 20846
rect 17033 20843 17099 20846
rect 35801 20843 35867 20846
rect 20478 20708 20484 20772
rect 20548 20770 20554 20772
rect 26141 20770 26207 20773
rect 20548 20768 26207 20770
rect 20548 20712 26146 20768
rect 26202 20712 26207 20768
rect 20548 20710 26207 20712
rect 20548 20708 20554 20710
rect 26141 20707 26207 20710
rect 27654 20708 27660 20772
rect 27724 20770 27730 20772
rect 27981 20770 28047 20773
rect 27724 20768 28047 20770
rect 27724 20712 27986 20768
rect 28042 20712 28047 20768
rect 27724 20710 28047 20712
rect 27724 20708 27730 20710
rect 27981 20707 28047 20710
rect 34094 20708 34100 20772
rect 34164 20770 34170 20772
rect 34513 20770 34579 20773
rect 34164 20768 34579 20770
rect 34164 20712 34518 20768
rect 34574 20712 34579 20768
rect 34164 20710 34579 20712
rect 34164 20708 34170 20710
rect 34513 20707 34579 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 8293 20636 8359 20637
rect 16205 20636 16271 20637
rect 8293 20632 8340 20636
rect 8404 20634 8410 20636
rect 8293 20576 8298 20632
rect 8293 20572 8340 20576
rect 8404 20574 8450 20634
rect 16205 20632 16252 20636
rect 16316 20634 16322 20636
rect 26509 20634 26575 20637
rect 16205 20576 16210 20632
rect 8404 20572 8410 20574
rect 16205 20572 16252 20576
rect 16316 20574 16362 20634
rect 26509 20632 27124 20634
rect 26509 20576 26514 20632
rect 26570 20576 27124 20632
rect 26509 20574 27124 20576
rect 16316 20572 16322 20574
rect 8293 20571 8359 20572
rect 16205 20571 16271 20572
rect 26509 20571 26575 20574
rect 27064 20501 27124 20574
rect 5073 20498 5139 20501
rect 5942 20498 5948 20500
rect 5073 20496 5948 20498
rect 5073 20440 5078 20496
rect 5134 20440 5948 20496
rect 5073 20438 5948 20440
rect 5073 20435 5139 20438
rect 5942 20436 5948 20438
rect 6012 20436 6018 20500
rect 8109 20498 8175 20501
rect 9121 20498 9187 20501
rect 8109 20496 9187 20498
rect 8109 20440 8114 20496
rect 8170 20440 9126 20496
rect 9182 20440 9187 20496
rect 8109 20438 9187 20440
rect 8109 20435 8175 20438
rect 9121 20435 9187 20438
rect 17585 20498 17651 20501
rect 21081 20498 21147 20501
rect 17585 20496 21147 20498
rect 17585 20440 17590 20496
rect 17646 20440 21086 20496
rect 21142 20440 21147 20496
rect 17585 20438 21147 20440
rect 17585 20435 17651 20438
rect 21081 20435 21147 20438
rect 27061 20498 27127 20501
rect 28257 20498 28323 20501
rect 27061 20496 28323 20498
rect 27061 20440 27066 20496
rect 27122 20440 28262 20496
rect 28318 20440 28323 20496
rect 27061 20438 28323 20440
rect 27061 20435 27127 20438
rect 28257 20435 28323 20438
rect 7005 20362 7071 20365
rect 9397 20362 9463 20365
rect 7005 20360 9463 20362
rect 7005 20304 7010 20360
rect 7066 20304 9402 20360
rect 9458 20304 9463 20360
rect 7005 20302 9463 20304
rect 7005 20299 7071 20302
rect 9397 20299 9463 20302
rect 16665 20362 16731 20365
rect 18321 20362 18387 20365
rect 19241 20362 19307 20365
rect 16665 20360 19307 20362
rect 16665 20304 16670 20360
rect 16726 20304 18326 20360
rect 18382 20304 19246 20360
rect 19302 20304 19307 20360
rect 16665 20302 19307 20304
rect 16665 20299 16731 20302
rect 18321 20299 18387 20302
rect 19241 20299 19307 20302
rect 20805 20362 20871 20365
rect 23289 20362 23355 20365
rect 23657 20362 23723 20365
rect 20805 20360 23723 20362
rect 20805 20304 20810 20360
rect 20866 20304 23294 20360
rect 23350 20304 23662 20360
rect 23718 20304 23723 20360
rect 20805 20302 23723 20304
rect 20805 20299 20871 20302
rect 23289 20299 23355 20302
rect 23657 20299 23723 20302
rect 10869 20226 10935 20229
rect 11646 20226 11652 20228
rect 10869 20224 11652 20226
rect 10869 20168 10874 20224
rect 10930 20168 11652 20224
rect 10869 20166 11652 20168
rect 10869 20163 10935 20166
rect 11646 20164 11652 20166
rect 11716 20164 11722 20228
rect 14641 20226 14707 20229
rect 17217 20226 17283 20229
rect 14641 20224 17283 20226
rect 14641 20168 14646 20224
rect 14702 20168 17222 20224
rect 17278 20168 17283 20224
rect 14641 20166 17283 20168
rect 14641 20163 14707 20166
rect 17217 20163 17283 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 16757 20090 16823 20093
rect 17953 20090 18019 20093
rect 16757 20088 18019 20090
rect 16757 20032 16762 20088
rect 16818 20032 17958 20088
rect 18014 20032 18019 20088
rect 16757 20030 18019 20032
rect 16757 20027 16823 20030
rect 17953 20027 18019 20030
rect 5533 19954 5599 19957
rect 5758 19954 5764 19956
rect 5533 19952 5764 19954
rect 5533 19896 5538 19952
rect 5594 19896 5764 19952
rect 5533 19894 5764 19896
rect 5533 19891 5599 19894
rect 5758 19892 5764 19894
rect 5828 19892 5834 19956
rect 8937 19954 9003 19957
rect 9581 19954 9647 19957
rect 8937 19952 9647 19954
rect 8937 19896 8942 19952
rect 8998 19896 9586 19952
rect 9642 19896 9647 19952
rect 8937 19894 9647 19896
rect 8937 19891 9003 19894
rect 9581 19891 9647 19894
rect 3785 19818 3851 19821
rect 19241 19818 19307 19821
rect 25957 19820 26023 19821
rect 25957 19818 26004 19820
rect 3785 19816 19307 19818
rect 3785 19760 3790 19816
rect 3846 19760 19246 19816
rect 19302 19760 19307 19816
rect 3785 19758 19307 19760
rect 25912 19816 26004 19818
rect 25912 19760 25962 19816
rect 25912 19758 26004 19760
rect 3785 19755 3851 19758
rect 19241 19755 19307 19758
rect 25957 19756 26004 19758
rect 26068 19756 26074 19820
rect 25957 19755 26023 19756
rect 14549 19682 14615 19685
rect 14774 19682 14780 19684
rect 14549 19680 14780 19682
rect 14549 19624 14554 19680
rect 14610 19624 14780 19680
rect 14549 19622 14780 19624
rect 14549 19619 14615 19622
rect 14774 19620 14780 19622
rect 14844 19682 14850 19684
rect 20846 19682 20852 19684
rect 14844 19622 20852 19682
rect 14844 19620 14850 19622
rect 20846 19620 20852 19622
rect 20916 19620 20922 19684
rect 22553 19682 22619 19685
rect 23289 19682 23355 19685
rect 22553 19680 23355 19682
rect 22553 19624 22558 19680
rect 22614 19624 23294 19680
rect 23350 19624 23355 19680
rect 22553 19622 23355 19624
rect 22553 19619 22619 19622
rect 23289 19619 23355 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 8661 19546 8727 19549
rect 9121 19546 9187 19549
rect 9397 19546 9463 19549
rect 8661 19544 9463 19546
rect 8661 19488 8666 19544
rect 8722 19488 9126 19544
rect 9182 19488 9402 19544
rect 9458 19488 9463 19544
rect 8661 19486 9463 19488
rect 8661 19483 8727 19486
rect 9121 19483 9187 19486
rect 9397 19483 9463 19486
rect 16798 19484 16804 19548
rect 16868 19546 16874 19548
rect 17033 19546 17099 19549
rect 22645 19546 22711 19549
rect 16868 19544 22711 19546
rect 16868 19488 17038 19544
rect 17094 19488 22650 19544
rect 22706 19488 22711 19544
rect 16868 19486 22711 19488
rect 16868 19484 16874 19486
rect 17033 19483 17099 19486
rect 22645 19483 22711 19486
rect 23197 19546 23263 19549
rect 31150 19546 31156 19548
rect 23197 19544 31156 19546
rect 23197 19488 23202 19544
rect 23258 19488 31156 19544
rect 23197 19486 31156 19488
rect 23197 19483 23263 19486
rect 31150 19484 31156 19486
rect 31220 19484 31226 19548
rect 7833 19412 7899 19413
rect 7782 19348 7788 19412
rect 7852 19410 7899 19412
rect 7852 19408 7944 19410
rect 7894 19352 7944 19408
rect 7852 19350 7944 19352
rect 7852 19348 7899 19350
rect 8702 19348 8708 19412
rect 8772 19410 8778 19412
rect 8937 19410 9003 19413
rect 8772 19408 9003 19410
rect 8772 19352 8942 19408
rect 8998 19352 9003 19408
rect 8772 19350 9003 19352
rect 8772 19348 8778 19350
rect 7833 19347 7899 19348
rect 8937 19347 9003 19350
rect 9305 19410 9371 19413
rect 10593 19410 10659 19413
rect 9305 19408 10659 19410
rect 9305 19352 9310 19408
rect 9366 19352 10598 19408
rect 10654 19352 10659 19408
rect 9305 19350 10659 19352
rect 9305 19347 9371 19350
rect 10593 19347 10659 19350
rect 16614 19348 16620 19412
rect 16684 19410 16690 19412
rect 16757 19410 16823 19413
rect 16684 19408 16823 19410
rect 16684 19352 16762 19408
rect 16818 19352 16823 19408
rect 16684 19350 16823 19352
rect 16684 19348 16690 19350
rect 16757 19347 16823 19350
rect 19977 19410 20043 19413
rect 19977 19408 20730 19410
rect 19977 19352 19982 19408
rect 20038 19352 20730 19408
rect 19977 19350 20730 19352
rect 19977 19347 20043 19350
rect 15745 19276 15811 19277
rect 15694 19274 15700 19276
rect 15654 19214 15700 19274
rect 15764 19272 15811 19276
rect 15806 19216 15811 19272
rect 15694 19212 15700 19214
rect 15764 19212 15811 19216
rect 20670 19274 20730 19350
rect 22134 19348 22140 19412
rect 22204 19410 22210 19412
rect 22553 19410 22619 19413
rect 22829 19412 22895 19413
rect 22829 19410 22876 19412
rect 22204 19408 22619 19410
rect 22204 19352 22558 19408
rect 22614 19352 22619 19408
rect 22204 19350 22619 19352
rect 22784 19408 22876 19410
rect 22784 19352 22834 19408
rect 22784 19350 22876 19352
rect 22204 19348 22210 19350
rect 22553 19347 22619 19350
rect 22829 19348 22876 19350
rect 22940 19348 22946 19412
rect 23197 19410 23263 19413
rect 24117 19410 24183 19413
rect 30373 19412 30439 19413
rect 25262 19410 25268 19412
rect 23197 19408 25268 19410
rect 23197 19352 23202 19408
rect 23258 19352 24122 19408
rect 24178 19352 25268 19408
rect 23197 19350 25268 19352
rect 22829 19347 22895 19348
rect 23197 19347 23263 19350
rect 24117 19347 24183 19350
rect 25262 19348 25268 19350
rect 25332 19348 25338 19412
rect 30373 19410 30420 19412
rect 30292 19408 30420 19410
rect 30484 19410 30490 19412
rect 31293 19410 31359 19413
rect 30484 19408 31359 19410
rect 30292 19352 30378 19408
rect 30484 19352 31298 19408
rect 31354 19352 31359 19408
rect 30292 19350 30420 19352
rect 30373 19348 30420 19350
rect 30484 19350 31359 19352
rect 30484 19348 30490 19350
rect 30373 19347 30439 19348
rect 31293 19347 31359 19350
rect 23289 19274 23355 19277
rect 25589 19274 25655 19277
rect 20670 19214 22110 19274
rect 15745 19211 15811 19212
rect 8753 19138 8819 19141
rect 10041 19138 10107 19141
rect 12065 19138 12131 19141
rect 8753 19136 12131 19138
rect 8753 19080 8758 19136
rect 8814 19080 10046 19136
rect 10102 19080 12070 19136
rect 12126 19080 12131 19136
rect 8753 19078 12131 19080
rect 8753 19075 8819 19078
rect 10041 19075 10107 19078
rect 12065 19075 12131 19078
rect 18229 19138 18295 19141
rect 21214 19138 21220 19140
rect 18229 19136 21220 19138
rect 18229 19080 18234 19136
rect 18290 19080 21220 19136
rect 18229 19078 21220 19080
rect 18229 19075 18295 19078
rect 21214 19076 21220 19078
rect 21284 19076 21290 19140
rect 22050 19138 22110 19214
rect 23289 19272 25655 19274
rect 23289 19216 23294 19272
rect 23350 19216 25594 19272
rect 25650 19216 25655 19272
rect 23289 19214 25655 19216
rect 23289 19211 23355 19214
rect 25589 19211 25655 19214
rect 35249 19274 35315 19277
rect 35382 19274 35388 19276
rect 35249 19272 35388 19274
rect 35249 19216 35254 19272
rect 35310 19216 35388 19272
rect 35249 19214 35388 19216
rect 35249 19211 35315 19214
rect 35382 19212 35388 19214
rect 35452 19212 35458 19276
rect 26601 19138 26667 19141
rect 22050 19136 26667 19138
rect 22050 19080 26606 19136
rect 26662 19080 26667 19136
rect 22050 19078 26667 19080
rect 26601 19075 26667 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 16757 19002 16823 19005
rect 16982 19002 16988 19004
rect 16757 19000 16988 19002
rect 16757 18944 16762 19000
rect 16818 18944 16988 19000
rect 16757 18942 16988 18944
rect 16757 18939 16823 18942
rect 16982 18940 16988 18942
rect 17052 18940 17058 19004
rect 18638 18940 18644 19004
rect 18708 19002 18714 19004
rect 21030 19002 21036 19004
rect 18708 18942 21036 19002
rect 18708 18940 18714 18942
rect 21030 18940 21036 18942
rect 21100 18940 21106 19004
rect 3877 18868 3943 18869
rect 3877 18864 3924 18868
rect 3988 18866 3994 18868
rect 3877 18808 3882 18864
rect 3877 18804 3924 18808
rect 3988 18806 4034 18866
rect 3988 18804 3994 18806
rect 12750 18804 12756 18868
rect 12820 18866 12826 18868
rect 18137 18866 18203 18869
rect 12820 18864 18203 18866
rect 12820 18808 18142 18864
rect 18198 18808 18203 18864
rect 12820 18806 18203 18808
rect 12820 18804 12826 18806
rect 3877 18803 3943 18804
rect 18137 18803 18203 18806
rect 23289 18866 23355 18869
rect 24894 18866 24900 18868
rect 23289 18864 24900 18866
rect 23289 18808 23294 18864
rect 23350 18808 24900 18864
rect 23289 18806 24900 18808
rect 23289 18803 23355 18806
rect 24894 18804 24900 18806
rect 24964 18866 24970 18868
rect 25129 18866 25195 18869
rect 24964 18864 25195 18866
rect 24964 18808 25134 18864
rect 25190 18808 25195 18864
rect 24964 18806 25195 18808
rect 24964 18804 24970 18806
rect 25129 18803 25195 18806
rect 26693 18868 26759 18869
rect 26693 18864 26740 18868
rect 26804 18866 26810 18868
rect 26693 18808 26698 18864
rect 26693 18804 26740 18808
rect 26804 18806 26850 18866
rect 26804 18804 26810 18806
rect 26693 18803 26759 18804
rect 11789 18730 11855 18733
rect 12985 18730 13051 18733
rect 11789 18728 13051 18730
rect 11789 18672 11794 18728
rect 11850 18672 12990 18728
rect 13046 18672 13051 18728
rect 11789 18670 13051 18672
rect 11789 18667 11855 18670
rect 12985 18667 13051 18670
rect 25589 18730 25655 18733
rect 27654 18730 27660 18732
rect 25589 18728 27660 18730
rect 25589 18672 25594 18728
rect 25650 18672 27660 18728
rect 25589 18670 27660 18672
rect 25589 18667 25655 18670
rect 27654 18668 27660 18670
rect 27724 18668 27730 18732
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 7598 18396 7604 18460
rect 7668 18458 7674 18460
rect 7741 18458 7807 18461
rect 7668 18456 7807 18458
rect 7668 18400 7746 18456
rect 7802 18400 7807 18456
rect 7668 18398 7807 18400
rect 7668 18396 7674 18398
rect 7741 18395 7807 18398
rect 23933 18458 23999 18461
rect 23933 18456 24042 18458
rect 23933 18400 23938 18456
rect 23994 18400 24042 18456
rect 23933 18395 24042 18400
rect 18597 18322 18663 18325
rect 19701 18322 19767 18325
rect 23982 18322 24042 18395
rect 24669 18322 24735 18325
rect 18597 18320 24735 18322
rect 18597 18264 18602 18320
rect 18658 18264 19706 18320
rect 19762 18264 24674 18320
rect 24730 18264 24735 18320
rect 18597 18262 24735 18264
rect 18597 18259 18663 18262
rect 19701 18259 19767 18262
rect 24669 18259 24735 18262
rect 25405 18322 25471 18325
rect 25630 18322 25636 18324
rect 25405 18320 25636 18322
rect 25405 18264 25410 18320
rect 25466 18264 25636 18320
rect 25405 18262 25636 18264
rect 25405 18259 25471 18262
rect 25630 18260 25636 18262
rect 25700 18260 25706 18324
rect 27429 18322 27495 18325
rect 28022 18322 28028 18324
rect 25822 18320 28028 18322
rect 25822 18264 27434 18320
rect 27490 18264 28028 18320
rect 25822 18262 28028 18264
rect 4429 18186 4495 18189
rect 8477 18186 8543 18189
rect 10409 18186 10475 18189
rect 14917 18186 14983 18189
rect 4429 18184 4676 18186
rect 4429 18128 4434 18184
rect 4490 18128 4676 18184
rect 4429 18126 4676 18128
rect 4429 18123 4495 18126
rect 4616 18053 4676 18126
rect 8477 18184 14983 18186
rect 8477 18128 8482 18184
rect 8538 18128 10414 18184
rect 10470 18128 14922 18184
rect 14978 18128 14983 18184
rect 8477 18126 14983 18128
rect 8477 18123 8543 18126
rect 10409 18123 10475 18126
rect 14917 18123 14983 18126
rect 15326 18124 15332 18188
rect 15396 18186 15402 18188
rect 18270 18186 18276 18188
rect 15396 18126 18276 18186
rect 15396 18124 15402 18126
rect 18270 18124 18276 18126
rect 18340 18124 18346 18188
rect 21541 18186 21607 18189
rect 23105 18186 23171 18189
rect 21541 18184 23171 18186
rect 21541 18128 21546 18184
rect 21602 18128 23110 18184
rect 23166 18128 23171 18184
rect 21541 18126 23171 18128
rect 21541 18123 21607 18126
rect 23105 18123 23171 18126
rect 23606 18124 23612 18188
rect 23676 18186 23682 18188
rect 24577 18186 24643 18189
rect 25822 18186 25882 18262
rect 27429 18259 27495 18262
rect 28022 18260 28028 18262
rect 28092 18260 28098 18324
rect 26141 18188 26207 18189
rect 26141 18186 26188 18188
rect 23676 18184 25882 18186
rect 23676 18128 24582 18184
rect 24638 18128 25882 18184
rect 23676 18126 25882 18128
rect 26096 18184 26188 18186
rect 26096 18128 26146 18184
rect 26096 18126 26188 18128
rect 23676 18124 23682 18126
rect 24577 18123 24643 18126
rect 26141 18124 26188 18126
rect 26252 18124 26258 18188
rect 32070 18124 32076 18188
rect 32140 18186 32146 18188
rect 32806 18186 32812 18188
rect 32140 18126 32812 18186
rect 32140 18124 32146 18126
rect 32806 18124 32812 18126
rect 32876 18186 32882 18188
rect 32949 18186 33015 18189
rect 32876 18184 33015 18186
rect 32876 18128 32954 18184
rect 33010 18128 33015 18184
rect 32876 18126 33015 18128
rect 32876 18124 32882 18126
rect 26141 18123 26207 18124
rect 32949 18123 33015 18126
rect 4613 18048 4679 18053
rect 4613 17992 4618 18048
rect 4674 17992 4679 18048
rect 4613 17987 4679 17992
rect 16113 18050 16179 18053
rect 21909 18052 21975 18053
rect 23933 18052 23999 18053
rect 19374 18050 19380 18052
rect 16113 18048 19380 18050
rect 16113 17992 16118 18048
rect 16174 17992 19380 18048
rect 16113 17990 19380 17992
rect 16113 17987 16179 17990
rect 19374 17988 19380 17990
rect 19444 17988 19450 18052
rect 21909 18048 21956 18052
rect 22020 18050 22026 18052
rect 21909 17992 21914 18048
rect 21909 17988 21956 17992
rect 22020 17990 22066 18050
rect 23933 18048 23980 18052
rect 24044 18050 24050 18052
rect 23933 17992 23938 18048
rect 22020 17988 22026 17990
rect 23933 17988 23980 17992
rect 24044 17990 24090 18050
rect 24044 17988 24050 17990
rect 24158 17988 24164 18052
rect 24228 18050 24234 18052
rect 24894 18050 24900 18052
rect 24228 17990 24900 18050
rect 24228 17988 24234 17990
rect 24894 17988 24900 17990
rect 24964 17988 24970 18052
rect 21909 17987 21975 17988
rect 23933 17987 23999 17988
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 34930 17984 35246 17985
rect 4210 17919 4526 17920
rect 10593 17968 10659 17973
rect 4705 17916 4771 17917
rect 4654 17852 4660 17916
rect 4724 17914 4771 17916
rect 9857 17914 9923 17917
rect 10358 17914 10364 17916
rect 4724 17912 4816 17914
rect 4766 17856 4816 17912
rect 4724 17854 4816 17856
rect 9857 17912 10364 17914
rect 9857 17856 9862 17912
rect 9918 17856 10364 17912
rect 9857 17854 10364 17856
rect 4724 17852 4771 17854
rect 4705 17851 4771 17852
rect 9857 17851 9923 17854
rect 10358 17852 10364 17854
rect 10428 17852 10434 17916
rect 10593 17912 10598 17968
rect 10654 17914 10659 17968
rect 10869 17970 10935 17973
rect 10869 17968 10978 17970
rect 10726 17914 10732 17916
rect 10654 17912 10732 17914
rect 10593 17907 10732 17912
rect 10596 17854 10732 17907
rect 10726 17852 10732 17854
rect 10796 17852 10802 17916
rect 10869 17912 10874 17968
rect 10930 17914 10978 17968
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 10930 17912 12082 17914
rect 10869 17907 12082 17912
rect 10918 17854 12082 17907
rect 4337 17778 4403 17781
rect 5441 17778 5507 17781
rect 4337 17776 5507 17778
rect 4337 17720 4342 17776
rect 4398 17720 5446 17776
rect 5502 17720 5507 17776
rect 4337 17718 5507 17720
rect 4337 17715 4403 17718
rect 5441 17715 5507 17718
rect 10542 17716 10548 17780
rect 10612 17778 10618 17780
rect 10777 17778 10843 17781
rect 10612 17776 10843 17778
rect 10612 17720 10782 17776
rect 10838 17720 10843 17776
rect 10612 17718 10843 17720
rect 10612 17716 10618 17718
rect 10777 17715 10843 17718
rect 11053 17778 11119 17781
rect 11329 17778 11395 17781
rect 11053 17776 11395 17778
rect 11053 17720 11058 17776
rect 11114 17720 11334 17776
rect 11390 17720 11395 17776
rect 11053 17718 11395 17720
rect 12022 17778 12082 17854
rect 12249 17778 12315 17781
rect 12022 17776 12315 17778
rect 12022 17720 12254 17776
rect 12310 17720 12315 17776
rect 12022 17718 12315 17720
rect 11053 17715 11119 17718
rect 11329 17715 11395 17718
rect 12249 17715 12315 17718
rect 21173 17778 21239 17781
rect 25497 17778 25563 17781
rect 21173 17776 25563 17778
rect 21173 17720 21178 17776
rect 21234 17720 25502 17776
rect 25558 17720 25563 17776
rect 21173 17718 25563 17720
rect 21173 17715 21239 17718
rect 25497 17715 25563 17718
rect 3693 17642 3759 17645
rect 4889 17642 4955 17645
rect 3693 17640 4955 17642
rect 3693 17584 3698 17640
rect 3754 17584 4894 17640
rect 4950 17584 4955 17640
rect 3693 17582 4955 17584
rect 3693 17579 3759 17582
rect 4889 17579 4955 17582
rect 10041 17642 10107 17645
rect 10174 17642 10180 17644
rect 10041 17640 10180 17642
rect 10041 17584 10046 17640
rect 10102 17584 10180 17640
rect 10041 17582 10180 17584
rect 10041 17579 10107 17582
rect 10174 17580 10180 17582
rect 10244 17580 10250 17644
rect 21633 17642 21699 17645
rect 22829 17642 22895 17645
rect 28206 17642 28212 17644
rect 21633 17640 28212 17642
rect 21633 17584 21638 17640
rect 21694 17584 22834 17640
rect 22890 17584 28212 17640
rect 21633 17582 28212 17584
rect 21633 17579 21699 17582
rect 22829 17579 22895 17582
rect 28206 17580 28212 17582
rect 28276 17580 28282 17644
rect 9213 17506 9279 17509
rect 11421 17506 11487 17509
rect 9213 17504 11487 17506
rect 9213 17448 9218 17504
rect 9274 17448 11426 17504
rect 11482 17448 11487 17504
rect 9213 17446 11487 17448
rect 9213 17443 9279 17446
rect 11421 17443 11487 17446
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 4245 17370 4311 17373
rect 4705 17370 4771 17373
rect 4245 17368 4771 17370
rect 4245 17312 4250 17368
rect 4306 17312 4710 17368
rect 4766 17312 4771 17368
rect 4245 17310 4771 17312
rect 4245 17307 4311 17310
rect 4705 17307 4771 17310
rect 9806 17308 9812 17372
rect 9876 17370 9882 17372
rect 9949 17370 10015 17373
rect 9876 17368 10015 17370
rect 9876 17312 9954 17368
rect 10010 17312 10015 17368
rect 9876 17310 10015 17312
rect 9876 17308 9882 17310
rect 9949 17307 10015 17310
rect 10133 17370 10199 17373
rect 10409 17370 10475 17373
rect 10133 17368 10475 17370
rect 10133 17312 10138 17368
rect 10194 17312 10414 17368
rect 10470 17312 10475 17368
rect 10133 17310 10475 17312
rect 10133 17307 10199 17310
rect 10409 17307 10475 17310
rect 10777 17370 10843 17373
rect 11605 17370 11671 17373
rect 10777 17368 11671 17370
rect 10777 17312 10782 17368
rect 10838 17312 11610 17368
rect 11666 17312 11671 17368
rect 10777 17310 11671 17312
rect 10777 17307 10843 17310
rect 11605 17307 11671 17310
rect 12934 17308 12940 17372
rect 13004 17370 13010 17372
rect 13077 17370 13143 17373
rect 13537 17370 13603 17373
rect 13004 17368 13603 17370
rect 13004 17312 13082 17368
rect 13138 17312 13542 17368
rect 13598 17312 13603 17368
rect 13004 17310 13603 17312
rect 13004 17308 13010 17310
rect 13077 17307 13143 17310
rect 13537 17307 13603 17310
rect 15142 17308 15148 17372
rect 15212 17370 15218 17372
rect 15285 17370 15351 17373
rect 15212 17368 15351 17370
rect 15212 17312 15290 17368
rect 15346 17312 15351 17368
rect 15212 17310 15351 17312
rect 15212 17308 15218 17310
rect 15285 17307 15351 17310
rect 22461 17370 22527 17373
rect 23013 17370 23079 17373
rect 22461 17368 23079 17370
rect 22461 17312 22466 17368
rect 22522 17312 23018 17368
rect 23074 17312 23079 17368
rect 22461 17310 23079 17312
rect 22461 17307 22527 17310
rect 23013 17307 23079 17310
rect 30649 17370 30715 17373
rect 35382 17370 35388 17372
rect 30649 17368 35388 17370
rect 30649 17312 30654 17368
rect 30710 17312 35388 17368
rect 30649 17310 35388 17312
rect 30649 17307 30715 17310
rect 35382 17308 35388 17310
rect 35452 17308 35458 17372
rect 9581 17234 9647 17237
rect 9949 17234 10015 17237
rect 9581 17232 10015 17234
rect 9581 17176 9586 17232
rect 9642 17176 9954 17232
rect 10010 17176 10015 17232
rect 9581 17174 10015 17176
rect 9581 17171 9647 17174
rect 9949 17171 10015 17174
rect 10358 17172 10364 17236
rect 10428 17234 10434 17236
rect 10961 17234 11027 17237
rect 10428 17232 11027 17234
rect 10428 17176 10966 17232
rect 11022 17176 11027 17232
rect 10428 17174 11027 17176
rect 10428 17172 10434 17174
rect 10961 17171 11027 17174
rect 22553 17234 22619 17237
rect 25630 17234 25636 17236
rect 22553 17232 25636 17234
rect 22553 17176 22558 17232
rect 22614 17176 25636 17232
rect 22553 17174 25636 17176
rect 22553 17171 22619 17174
rect 25630 17172 25636 17174
rect 25700 17172 25706 17236
rect 10726 17036 10732 17100
rect 10796 17098 10802 17100
rect 13721 17098 13787 17101
rect 10796 17096 13787 17098
rect 10796 17040 13726 17096
rect 13782 17040 13787 17096
rect 10796 17038 13787 17040
rect 10796 17036 10802 17038
rect 13721 17035 13787 17038
rect 18045 17098 18111 17101
rect 20478 17098 20484 17100
rect 18045 17096 20484 17098
rect 18045 17040 18050 17096
rect 18106 17040 20484 17096
rect 18045 17038 20484 17040
rect 18045 17035 18111 17038
rect 20478 17036 20484 17038
rect 20548 17036 20554 17100
rect 27613 17098 27679 17101
rect 28574 17098 28580 17100
rect 27613 17096 28580 17098
rect 27613 17040 27618 17096
rect 27674 17040 28580 17096
rect 27613 17038 28580 17040
rect 27613 17035 27679 17038
rect 28574 17036 28580 17038
rect 28644 17036 28650 17100
rect 10542 16900 10548 16964
rect 10612 16962 10618 16964
rect 10777 16962 10843 16965
rect 10612 16960 10843 16962
rect 10612 16904 10782 16960
rect 10838 16904 10843 16960
rect 10612 16902 10843 16904
rect 10612 16900 10618 16902
rect 10777 16899 10843 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 21909 16826 21975 16829
rect 25446 16826 25452 16828
rect 21909 16824 25452 16826
rect 21909 16768 21914 16824
rect 21970 16768 25452 16824
rect 21909 16766 25452 16768
rect 21909 16763 21975 16766
rect 25446 16764 25452 16766
rect 25516 16826 25522 16828
rect 26969 16826 27035 16829
rect 25516 16824 27035 16826
rect 25516 16768 26974 16824
rect 27030 16768 27035 16824
rect 25516 16766 27035 16768
rect 25516 16764 25522 16766
rect 26969 16763 27035 16766
rect 4521 16690 4587 16693
rect 4654 16690 4660 16692
rect 4521 16688 4660 16690
rect 4521 16632 4526 16688
rect 4582 16632 4660 16688
rect 4521 16630 4660 16632
rect 4521 16627 4587 16630
rect 4654 16628 4660 16630
rect 4724 16628 4730 16692
rect 12617 16690 12683 16693
rect 14958 16690 14964 16692
rect 12617 16688 14964 16690
rect 12617 16632 12622 16688
rect 12678 16632 14964 16688
rect 12617 16630 14964 16632
rect 12617 16627 12683 16630
rect 14958 16628 14964 16630
rect 15028 16628 15034 16692
rect 26366 16628 26372 16692
rect 26436 16690 26442 16692
rect 26509 16690 26575 16693
rect 26436 16688 26575 16690
rect 26436 16632 26514 16688
rect 26570 16632 26575 16688
rect 26436 16630 26575 16632
rect 26436 16628 26442 16630
rect 26509 16627 26575 16630
rect 3325 16554 3391 16557
rect 4429 16554 4495 16557
rect 3325 16552 4495 16554
rect 3325 16496 3330 16552
rect 3386 16496 4434 16552
rect 4490 16496 4495 16552
rect 3325 16494 4495 16496
rect 3325 16491 3391 16494
rect 4429 16491 4495 16494
rect 35249 16554 35315 16557
rect 35249 16552 36140 16554
rect 35249 16496 35254 16552
rect 35310 16496 36140 16552
rect 35249 16494 36140 16496
rect 35249 16491 35315 16494
rect 22645 16420 22711 16421
rect 22645 16418 22692 16420
rect 22600 16416 22692 16418
rect 22600 16360 22650 16416
rect 22600 16358 22692 16360
rect 22645 16356 22692 16358
rect 22756 16356 22762 16420
rect 36080 16418 36140 16494
rect 36782 16418 37582 16448
rect 36080 16358 37582 16418
rect 22645 16355 22711 16356
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 36782 16328 37582 16358
rect 35590 16287 35906 16288
rect 17125 16284 17191 16285
rect 17125 16282 17172 16284
rect 17080 16280 17172 16282
rect 17080 16224 17130 16280
rect 17080 16222 17172 16224
rect 17125 16220 17172 16222
rect 17236 16220 17242 16284
rect 17125 16219 17191 16220
rect 2589 16146 2655 16149
rect 3877 16146 3943 16149
rect 7005 16146 7071 16149
rect 2589 16144 7071 16146
rect 2589 16088 2594 16144
rect 2650 16088 3882 16144
rect 3938 16088 7010 16144
rect 7066 16088 7071 16144
rect 2589 16086 7071 16088
rect 2589 16083 2655 16086
rect 3877 16083 3943 16086
rect 7005 16083 7071 16086
rect 12801 16146 12867 16149
rect 15745 16146 15811 16149
rect 12801 16144 15811 16146
rect 12801 16088 12806 16144
rect 12862 16088 15750 16144
rect 15806 16088 15811 16144
rect 12801 16086 15811 16088
rect 12801 16083 12867 16086
rect 15745 16083 15811 16086
rect 21633 16146 21699 16149
rect 27889 16146 27955 16149
rect 21633 16144 27955 16146
rect 21633 16088 21638 16144
rect 21694 16088 27894 16144
rect 27950 16088 27955 16144
rect 21633 16086 27955 16088
rect 21633 16083 21699 16086
rect 27889 16083 27955 16086
rect 34789 16146 34855 16149
rect 35525 16146 35591 16149
rect 34789 16144 35591 16146
rect 34789 16088 34794 16144
rect 34850 16088 35530 16144
rect 35586 16088 35591 16144
rect 34789 16086 35591 16088
rect 34789 16083 34855 16086
rect 35525 16083 35591 16086
rect 15193 16010 15259 16013
rect 16614 16010 16620 16012
rect 15193 16008 16620 16010
rect 15193 15952 15198 16008
rect 15254 15952 16620 16008
rect 15193 15950 16620 15952
rect 15193 15947 15259 15950
rect 16614 15948 16620 15950
rect 16684 15948 16690 16012
rect 22185 16010 22251 16013
rect 23013 16010 23079 16013
rect 22185 16008 23079 16010
rect 22185 15952 22190 16008
rect 22246 15952 23018 16008
rect 23074 15952 23079 16008
rect 22185 15950 23079 15952
rect 22185 15947 22251 15950
rect 23013 15947 23079 15950
rect 23473 16010 23539 16013
rect 23790 16010 23796 16012
rect 23473 16008 23796 16010
rect 23473 15952 23478 16008
rect 23534 15952 23796 16008
rect 23473 15950 23796 15952
rect 23473 15947 23539 15950
rect 23790 15948 23796 15950
rect 23860 16010 23866 16012
rect 23860 15950 35450 16010
rect 23860 15948 23866 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 35390 15738 35450 15950
rect 36782 15738 37582 15768
rect 35390 15678 37582 15738
rect 36782 15648 37582 15678
rect 8334 15540 8340 15604
rect 8404 15602 8410 15604
rect 8569 15602 8635 15605
rect 8404 15600 8635 15602
rect 8404 15544 8574 15600
rect 8630 15544 8635 15600
rect 8404 15542 8635 15544
rect 8404 15540 8410 15542
rect 8569 15539 8635 15542
rect 10041 15602 10107 15605
rect 31569 15604 31635 15605
rect 10174 15602 10180 15604
rect 10041 15600 10180 15602
rect 10041 15544 10046 15600
rect 10102 15544 10180 15600
rect 10041 15542 10180 15544
rect 10041 15539 10107 15542
rect 10174 15540 10180 15542
rect 10244 15540 10250 15604
rect 31518 15540 31524 15604
rect 31588 15602 31635 15604
rect 31588 15600 31680 15602
rect 31630 15544 31680 15600
rect 31588 15542 31680 15544
rect 31588 15540 31635 15542
rect 31569 15539 31635 15540
rect 23197 15466 23263 15469
rect 25078 15466 25084 15468
rect 23197 15464 25084 15466
rect 23197 15408 23202 15464
rect 23258 15408 25084 15464
rect 23197 15406 25084 15408
rect 23197 15403 23263 15406
rect 25078 15404 25084 15406
rect 25148 15404 25154 15468
rect 5257 15330 5323 15333
rect 8753 15330 8819 15333
rect 5257 15328 8819 15330
rect 5257 15272 5262 15328
rect 5318 15272 8758 15328
rect 8814 15272 8819 15328
rect 5257 15270 8819 15272
rect 5257 15267 5323 15270
rect 8753 15267 8819 15270
rect 21582 15268 21588 15332
rect 21652 15330 21658 15332
rect 22093 15330 22159 15333
rect 21652 15328 22159 15330
rect 21652 15272 22098 15328
rect 22154 15272 22159 15328
rect 21652 15270 22159 15272
rect 21652 15268 21658 15270
rect 22093 15267 22159 15270
rect 27613 15330 27679 15333
rect 29310 15330 29316 15332
rect 27613 15328 29316 15330
rect 27613 15272 27618 15328
rect 27674 15272 29316 15328
rect 27613 15270 29316 15272
rect 27613 15267 27679 15270
rect 29310 15268 29316 15270
rect 29380 15268 29386 15332
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 2630 15132 2636 15196
rect 2700 15194 2706 15196
rect 4613 15194 4679 15197
rect 2700 15192 4679 15194
rect 2700 15136 4618 15192
rect 4674 15136 4679 15192
rect 2700 15134 4679 15136
rect 2700 15132 2706 15134
rect 4613 15131 4679 15134
rect 10685 15194 10751 15197
rect 10910 15194 10916 15196
rect 10685 15192 10916 15194
rect 10685 15136 10690 15192
rect 10746 15136 10916 15192
rect 10685 15134 10916 15136
rect 10685 15131 10751 15134
rect 10910 15132 10916 15134
rect 10980 15132 10986 15196
rect 19241 15194 19307 15197
rect 19558 15194 19564 15196
rect 19241 15192 19564 15194
rect 19241 15136 19246 15192
rect 19302 15136 19564 15192
rect 19241 15134 19564 15136
rect 19241 15131 19307 15134
rect 19558 15132 19564 15134
rect 19628 15132 19634 15196
rect 32121 15194 32187 15197
rect 32254 15194 32260 15196
rect 32121 15192 32260 15194
rect 32121 15136 32126 15192
rect 32182 15136 32260 15192
rect 32121 15134 32260 15136
rect 32121 15131 32187 15134
rect 32254 15132 32260 15134
rect 32324 15132 32330 15196
rect 20805 15058 20871 15061
rect 21214 15058 21220 15060
rect 20805 15056 21220 15058
rect 20805 15000 20810 15056
rect 20866 15000 21220 15056
rect 20805 14998 21220 15000
rect 20805 14995 20871 14998
rect 21214 14996 21220 14998
rect 21284 15058 21290 15060
rect 21357 15058 21423 15061
rect 21284 15056 21423 15058
rect 21284 15000 21362 15056
rect 21418 15000 21423 15056
rect 21284 14998 21423 15000
rect 21284 14996 21290 14998
rect 21357 14995 21423 14998
rect 19333 14922 19399 14925
rect 19742 14922 19748 14924
rect 19333 14920 19748 14922
rect 19333 14864 19338 14920
rect 19394 14864 19748 14920
rect 19333 14862 19748 14864
rect 19333 14859 19399 14862
rect 19742 14860 19748 14862
rect 19812 14860 19818 14924
rect 20529 14922 20595 14925
rect 21030 14922 21036 14924
rect 20529 14920 21036 14922
rect 20529 14864 20534 14920
rect 20590 14864 21036 14920
rect 20529 14862 21036 14864
rect 20529 14859 20595 14862
rect 21030 14860 21036 14862
rect 21100 14922 21106 14924
rect 21265 14922 21331 14925
rect 21100 14920 21331 14922
rect 21100 14864 21270 14920
rect 21326 14864 21331 14920
rect 21100 14862 21331 14864
rect 21100 14860 21106 14862
rect 21265 14859 21331 14862
rect 22001 14922 22067 14925
rect 24209 14922 24275 14925
rect 25589 14922 25655 14925
rect 22001 14920 25655 14922
rect 22001 14864 22006 14920
rect 22062 14864 24214 14920
rect 24270 14864 25594 14920
rect 25650 14864 25655 14920
rect 22001 14862 25655 14864
rect 22001 14859 22067 14862
rect 24209 14859 24275 14862
rect 25589 14859 25655 14862
rect 26182 14860 26188 14924
rect 26252 14922 26258 14924
rect 27245 14922 27311 14925
rect 26252 14920 27311 14922
rect 26252 14864 27250 14920
rect 27306 14864 27311 14920
rect 26252 14862 27311 14864
rect 26252 14860 26258 14862
rect 27245 14859 27311 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 8661 14516 8727 14517
rect 9949 14516 10015 14517
rect 11237 14516 11303 14517
rect 8661 14514 8708 14516
rect 8616 14512 8708 14514
rect 8772 14514 8778 14516
rect 9254 14514 9260 14516
rect 8616 14456 8666 14512
rect 8616 14454 8708 14456
rect 8661 14452 8708 14454
rect 8772 14454 9260 14514
rect 8772 14452 8778 14454
rect 9254 14452 9260 14454
rect 9324 14452 9330 14516
rect 9949 14514 9996 14516
rect 9904 14512 9996 14514
rect 9904 14456 9954 14512
rect 9904 14454 9996 14456
rect 9949 14452 9996 14454
rect 10060 14452 10066 14516
rect 11237 14514 11284 14516
rect 11192 14512 11284 14514
rect 11192 14456 11242 14512
rect 11192 14454 11284 14456
rect 11237 14452 11284 14454
rect 11348 14452 11354 14516
rect 27286 14452 27292 14516
rect 27356 14514 27362 14516
rect 27705 14514 27771 14517
rect 27356 14512 27771 14514
rect 27356 14456 27710 14512
rect 27766 14456 27771 14512
rect 27356 14454 27771 14456
rect 27356 14452 27362 14454
rect 8661 14451 8727 14452
rect 9949 14451 10015 14452
rect 11237 14451 11303 14452
rect 27705 14451 27771 14454
rect 35065 14514 35131 14517
rect 35382 14514 35388 14516
rect 35065 14512 35388 14514
rect 35065 14456 35070 14512
rect 35126 14456 35388 14512
rect 35065 14454 35388 14456
rect 35065 14451 35131 14454
rect 35382 14452 35388 14454
rect 35452 14452 35458 14516
rect 20713 14378 20779 14381
rect 25773 14378 25839 14381
rect 20713 14376 25839 14378
rect 20713 14320 20718 14376
rect 20774 14320 25778 14376
rect 25834 14320 25839 14376
rect 20713 14318 25839 14320
rect 20713 14315 20779 14318
rect 25773 14315 25839 14318
rect 27613 14242 27679 14245
rect 28206 14242 28212 14244
rect 27613 14240 28212 14242
rect 27613 14184 27618 14240
rect 27674 14184 28212 14240
rect 27613 14182 28212 14184
rect 27613 14179 27679 14182
rect 28206 14180 28212 14182
rect 28276 14180 28282 14244
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 14774 13908 14780 13972
rect 14844 13970 14850 13972
rect 15009 13970 15075 13973
rect 14844 13968 15075 13970
rect 14844 13912 15014 13968
rect 15070 13912 15075 13968
rect 14844 13910 15075 13912
rect 14844 13908 14850 13910
rect 15009 13907 15075 13910
rect 19701 13970 19767 13973
rect 24209 13970 24275 13973
rect 24853 13970 24919 13973
rect 19701 13968 24919 13970
rect 19701 13912 19706 13968
rect 19762 13912 24214 13968
rect 24270 13912 24858 13968
rect 24914 13912 24919 13968
rect 19701 13910 24919 13912
rect 19701 13907 19767 13910
rect 24209 13907 24275 13910
rect 24853 13907 24919 13910
rect 4613 13836 4679 13837
rect 4613 13832 4660 13836
rect 4724 13834 4730 13836
rect 4613 13776 4618 13832
rect 4613 13772 4660 13776
rect 4724 13774 4770 13834
rect 27245 13832 27311 13837
rect 27245 13776 27250 13832
rect 27306 13776 27311 13832
rect 4724 13772 4730 13774
rect 4613 13771 4679 13772
rect 27245 13771 27311 13776
rect 30649 13834 30715 13837
rect 33685 13834 33751 13837
rect 30649 13832 33751 13834
rect 30649 13776 30654 13832
rect 30710 13776 33690 13832
rect 33746 13776 33751 13832
rect 30649 13774 33751 13776
rect 30649 13771 30715 13774
rect 33685 13771 33751 13774
rect 8293 13698 8359 13701
rect 9070 13698 9076 13700
rect 8293 13696 9076 13698
rect 8293 13640 8298 13696
rect 8354 13640 9076 13696
rect 8293 13638 9076 13640
rect 8293 13635 8359 13638
rect 9070 13636 9076 13638
rect 9140 13636 9146 13700
rect 27248 13698 27308 13771
rect 30598 13698 30604 13700
rect 27248 13638 30604 13698
rect 30598 13636 30604 13638
rect 30668 13636 30674 13700
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 15009 13562 15075 13565
rect 21541 13562 21607 13565
rect 15009 13560 21607 13562
rect 15009 13504 15014 13560
rect 15070 13504 21546 13560
rect 21602 13504 21607 13560
rect 15009 13502 21607 13504
rect 15009 13499 15075 13502
rect 21541 13499 21607 13502
rect 9397 13426 9463 13429
rect 10225 13426 10291 13429
rect 9397 13424 10291 13426
rect 9397 13368 9402 13424
rect 9458 13368 10230 13424
rect 10286 13368 10291 13424
rect 9397 13366 10291 13368
rect 9397 13363 9463 13366
rect 10225 13363 10291 13366
rect 19333 13426 19399 13429
rect 20161 13426 20227 13429
rect 19333 13424 20227 13426
rect 19333 13368 19338 13424
rect 19394 13368 20166 13424
rect 20222 13368 20227 13424
rect 19333 13366 20227 13368
rect 19333 13363 19399 13366
rect 20161 13363 20227 13366
rect 30046 13364 30052 13428
rect 30116 13426 30122 13428
rect 32489 13426 32555 13429
rect 30116 13424 32555 13426
rect 30116 13368 32494 13424
rect 32550 13368 32555 13424
rect 30116 13366 32555 13368
rect 30116 13364 30122 13366
rect 32489 13363 32555 13366
rect 5441 13290 5507 13293
rect 5574 13290 5580 13292
rect 5441 13288 5580 13290
rect 5441 13232 5446 13288
rect 5502 13232 5580 13288
rect 5441 13230 5580 13232
rect 5441 13227 5507 13230
rect 5574 13228 5580 13230
rect 5644 13228 5650 13292
rect 18873 13290 18939 13293
rect 19333 13290 19399 13293
rect 19885 13290 19951 13293
rect 18873 13288 19074 13290
rect 18873 13232 18878 13288
rect 18934 13232 19074 13288
rect 18873 13230 19074 13232
rect 18873 13227 18939 13230
rect 19014 13154 19074 13230
rect 19333 13288 19951 13290
rect 19333 13232 19338 13288
rect 19394 13232 19890 13288
rect 19946 13232 19951 13288
rect 19333 13230 19951 13232
rect 19333 13227 19399 13230
rect 19885 13227 19951 13230
rect 19149 13154 19215 13157
rect 19014 13152 19215 13154
rect 19014 13096 19154 13152
rect 19210 13096 19215 13152
rect 19014 13094 19215 13096
rect 19149 13091 19215 13094
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 19333 13020 19399 13021
rect 19333 13018 19380 13020
rect 19288 13016 19380 13018
rect 19288 12960 19338 13016
rect 19288 12958 19380 12960
rect 19333 12956 19380 12958
rect 19444 12956 19450 13020
rect 25998 12956 26004 13020
rect 26068 13018 26074 13020
rect 31569 13018 31635 13021
rect 26068 13016 31635 13018
rect 26068 12960 31574 13016
rect 31630 12960 31635 13016
rect 26068 12958 31635 12960
rect 26068 12956 26074 12958
rect 19333 12955 19399 12956
rect 31569 12955 31635 12958
rect 2037 12882 2103 12885
rect 3918 12882 3924 12884
rect 2037 12880 3924 12882
rect 2037 12824 2042 12880
rect 2098 12824 3924 12880
rect 2037 12822 3924 12824
rect 2037 12819 2103 12822
rect 3918 12820 3924 12822
rect 3988 12882 3994 12884
rect 4061 12882 4127 12885
rect 3988 12880 4127 12882
rect 3988 12824 4066 12880
rect 4122 12824 4127 12880
rect 3988 12822 4127 12824
rect 3988 12820 3994 12822
rect 4061 12819 4127 12822
rect 8477 12882 8543 12885
rect 10869 12882 10935 12885
rect 17585 12884 17651 12885
rect 17534 12882 17540 12884
rect 8477 12880 10935 12882
rect 8477 12824 8482 12880
rect 8538 12824 10874 12880
rect 10930 12824 10935 12880
rect 8477 12822 10935 12824
rect 17494 12822 17540 12882
rect 17604 12880 17651 12884
rect 17646 12824 17651 12880
rect 8477 12819 8543 12822
rect 10869 12819 10935 12822
rect 17534 12820 17540 12822
rect 17604 12820 17651 12824
rect 17585 12819 17651 12820
rect 3877 12746 3943 12749
rect 5533 12746 5599 12749
rect 6177 12746 6243 12749
rect 3877 12744 5599 12746
rect 3877 12688 3882 12744
rect 3938 12688 5538 12744
rect 5594 12688 5599 12744
rect 3877 12686 5599 12688
rect 3877 12683 3943 12686
rect 5533 12683 5599 12686
rect 6134 12744 6243 12746
rect 6134 12688 6182 12744
rect 6238 12688 6243 12744
rect 6134 12683 6243 12688
rect 7189 12748 7255 12749
rect 7189 12744 7236 12748
rect 7300 12746 7306 12748
rect 7189 12688 7194 12744
rect 7189 12684 7236 12688
rect 7300 12686 7346 12746
rect 7300 12684 7306 12686
rect 7189 12683 7255 12684
rect 4889 12610 4955 12613
rect 5165 12610 5231 12613
rect 4889 12608 5231 12610
rect 4889 12552 4894 12608
rect 4950 12552 5170 12608
rect 5226 12552 5231 12608
rect 4889 12550 5231 12552
rect 4889 12547 4955 12550
rect 5165 12547 5231 12550
rect 5809 12610 5875 12613
rect 6134 12610 6194 12683
rect 5809 12608 6194 12610
rect 5809 12552 5814 12608
rect 5870 12552 6194 12608
rect 5809 12550 6194 12552
rect 19333 12610 19399 12613
rect 21173 12610 21239 12613
rect 23565 12610 23631 12613
rect 19333 12608 23631 12610
rect 19333 12552 19338 12608
rect 19394 12552 21178 12608
rect 21234 12552 23570 12608
rect 23626 12552 23631 12608
rect 19333 12550 23631 12552
rect 5809 12547 5875 12550
rect 19333 12547 19399 12550
rect 21173 12547 21239 12550
rect 23565 12547 23631 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 4705 12474 4771 12477
rect 5758 12474 5764 12476
rect 4705 12472 5764 12474
rect 4705 12416 4710 12472
rect 4766 12416 5764 12472
rect 4705 12414 5764 12416
rect 4705 12411 4771 12414
rect 5758 12412 5764 12414
rect 5828 12474 5834 12476
rect 22277 12474 22343 12477
rect 23197 12474 23263 12477
rect 5828 12414 6930 12474
rect 5828 12412 5834 12414
rect 4337 12338 4403 12341
rect 6729 12338 6795 12341
rect 4337 12336 6795 12338
rect 4337 12280 4342 12336
rect 4398 12280 6734 12336
rect 6790 12280 6795 12336
rect 4337 12278 6795 12280
rect 4337 12275 4403 12278
rect 6729 12275 6795 12278
rect 4797 12202 4863 12205
rect 4662 12200 4863 12202
rect 4662 12144 4802 12200
rect 4858 12144 4863 12200
rect 4662 12142 4863 12144
rect 4662 11658 4722 12142
rect 4797 12139 4863 12142
rect 4981 12202 5047 12205
rect 6870 12202 6930 12414
rect 22277 12472 23263 12474
rect 22277 12416 22282 12472
rect 22338 12416 23202 12472
rect 23258 12416 23263 12472
rect 22277 12414 23263 12416
rect 22277 12411 22343 12414
rect 23197 12411 23263 12414
rect 26049 12474 26115 12477
rect 29269 12474 29335 12477
rect 26049 12472 29335 12474
rect 26049 12416 26054 12472
rect 26110 12416 29274 12472
rect 29330 12416 29335 12472
rect 26049 12414 29335 12416
rect 26049 12411 26115 12414
rect 29269 12411 29335 12414
rect 30422 12414 31034 12474
rect 17125 12338 17191 12341
rect 17677 12338 17743 12341
rect 17125 12336 17743 12338
rect 17125 12280 17130 12336
rect 17186 12280 17682 12336
rect 17738 12280 17743 12336
rect 17125 12278 17743 12280
rect 17125 12275 17191 12278
rect 17677 12275 17743 12278
rect 18321 12338 18387 12341
rect 30422 12338 30482 12414
rect 18321 12336 30482 12338
rect 18321 12280 18326 12336
rect 18382 12280 30482 12336
rect 18321 12278 30482 12280
rect 30557 12338 30623 12341
rect 30782 12338 30788 12340
rect 30557 12336 30788 12338
rect 30557 12280 30562 12336
rect 30618 12280 30788 12336
rect 30557 12278 30788 12280
rect 18321 12275 18387 12278
rect 30557 12275 30623 12278
rect 30782 12276 30788 12278
rect 30852 12276 30858 12340
rect 30974 12338 31034 12414
rect 32990 12338 32996 12340
rect 30974 12278 32996 12338
rect 32990 12276 32996 12278
rect 33060 12338 33066 12340
rect 34789 12338 34855 12341
rect 33060 12336 34855 12338
rect 33060 12280 34794 12336
rect 34850 12280 34855 12336
rect 33060 12278 34855 12280
rect 33060 12276 33066 12278
rect 34789 12275 34855 12278
rect 8017 12202 8083 12205
rect 4981 12200 5458 12202
rect 4981 12144 4986 12200
rect 5042 12144 5458 12200
rect 4981 12142 5458 12144
rect 6870 12200 8083 12202
rect 6870 12144 8022 12200
rect 8078 12144 8083 12200
rect 6870 12142 8083 12144
rect 4981 12139 5047 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 5257 11928 5323 11933
rect 5257 11872 5262 11928
rect 5318 11872 5323 11928
rect 5257 11867 5323 11872
rect 4889 11794 4955 11797
rect 5260 11794 5320 11867
rect 4889 11792 5320 11794
rect 4889 11736 4894 11792
rect 4950 11736 5320 11792
rect 4889 11734 5320 11736
rect 4889 11731 4955 11734
rect 5398 11661 5458 12142
rect 8017 12139 8083 12142
rect 16757 12202 16823 12205
rect 18597 12202 18663 12205
rect 21265 12202 21331 12205
rect 23841 12202 23907 12205
rect 16757 12200 18154 12202
rect 16757 12144 16762 12200
rect 16818 12144 18154 12200
rect 16757 12142 18154 12144
rect 16757 12139 16823 12142
rect 6913 12066 6979 12069
rect 7741 12066 7807 12069
rect 6913 12064 7807 12066
rect 6913 12008 6918 12064
rect 6974 12008 7746 12064
rect 7802 12008 7807 12064
rect 6913 12006 7807 12008
rect 6913 12003 6979 12006
rect 7741 12003 7807 12006
rect 8385 11930 8451 11933
rect 16665 11932 16731 11933
rect 8342 11928 8451 11930
rect 8342 11872 8390 11928
rect 8446 11872 8451 11928
rect 8342 11867 8451 11872
rect 16614 11868 16620 11932
rect 16684 11930 16731 11932
rect 18094 11930 18154 12142
rect 18597 12200 23907 12202
rect 18597 12144 18602 12200
rect 18658 12144 21270 12200
rect 21326 12144 23846 12200
rect 23902 12144 23907 12200
rect 18597 12142 23907 12144
rect 18597 12139 18663 12142
rect 21265 12139 21331 12142
rect 23841 12139 23907 12142
rect 32673 12202 32739 12205
rect 34973 12202 35039 12205
rect 36077 12202 36143 12205
rect 32673 12200 36143 12202
rect 32673 12144 32678 12200
rect 32734 12144 34978 12200
rect 35034 12144 36082 12200
rect 36138 12144 36143 12200
rect 32673 12142 36143 12144
rect 32673 12139 32739 12142
rect 34973 12139 35039 12142
rect 36077 12139 36143 12142
rect 23933 12066 23999 12069
rect 30649 12066 30715 12069
rect 23933 12064 30715 12066
rect 23933 12008 23938 12064
rect 23994 12008 30654 12064
rect 30710 12008 30715 12064
rect 23933 12006 30715 12008
rect 23933 12003 23999 12006
rect 30649 12003 30715 12006
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 24025 11930 24091 11933
rect 26693 11932 26759 11933
rect 26693 11930 26740 11932
rect 16684 11928 16776 11930
rect 16726 11872 16776 11928
rect 16684 11870 16776 11872
rect 18094 11928 24091 11930
rect 18094 11872 24030 11928
rect 24086 11872 24091 11928
rect 18094 11870 24091 11872
rect 26648 11928 26740 11930
rect 26648 11872 26698 11928
rect 26648 11870 26740 11872
rect 16684 11868 16731 11870
rect 16665 11867 16731 11868
rect 24025 11867 24091 11870
rect 26693 11868 26740 11870
rect 26804 11868 26810 11932
rect 27705 11930 27771 11933
rect 30925 11930 30991 11933
rect 27705 11928 30991 11930
rect 27705 11872 27710 11928
rect 27766 11872 30930 11928
rect 30986 11872 30991 11928
rect 27705 11870 30991 11872
rect 26693 11867 26759 11868
rect 27705 11867 27771 11870
rect 30925 11867 30991 11870
rect 31569 11930 31635 11933
rect 32949 11930 33015 11933
rect 31569 11928 33015 11930
rect 31569 11872 31574 11928
rect 31630 11872 32954 11928
rect 33010 11872 33015 11928
rect 31569 11870 33015 11872
rect 31569 11867 31635 11870
rect 32949 11867 33015 11870
rect 8342 11661 8402 11867
rect 17493 11794 17559 11797
rect 21449 11794 21515 11797
rect 17493 11792 21515 11794
rect 17493 11736 17498 11792
rect 17554 11736 21454 11792
rect 21510 11736 21515 11792
rect 17493 11734 21515 11736
rect 17493 11731 17559 11734
rect 21449 11731 21515 11734
rect 25078 11732 25084 11796
rect 25148 11794 25154 11796
rect 26182 11794 26188 11796
rect 25148 11734 26188 11794
rect 25148 11732 25154 11734
rect 26182 11732 26188 11734
rect 26252 11794 26258 11796
rect 27245 11794 27311 11797
rect 30097 11796 30163 11797
rect 26252 11792 27311 11794
rect 26252 11736 27250 11792
rect 27306 11736 27311 11792
rect 26252 11734 27311 11736
rect 26252 11732 26258 11734
rect 27245 11731 27311 11734
rect 30046 11732 30052 11796
rect 30116 11794 30163 11796
rect 30116 11792 30208 11794
rect 30158 11736 30208 11792
rect 30116 11734 30208 11736
rect 30116 11732 30163 11734
rect 30097 11731 30163 11732
rect 5165 11658 5231 11661
rect 4662 11656 5231 11658
rect 4662 11600 5170 11656
rect 5226 11600 5231 11656
rect 4662 11598 5231 11600
rect 5398 11656 5507 11661
rect 5398 11600 5446 11656
rect 5502 11600 5507 11656
rect 5398 11598 5507 11600
rect 8342 11656 8451 11661
rect 8342 11600 8390 11656
rect 8446 11600 8451 11656
rect 8342 11598 8451 11600
rect 5165 11595 5231 11598
rect 5441 11595 5507 11598
rect 8385 11595 8451 11598
rect 10593 11658 10659 11661
rect 26366 11658 26372 11660
rect 10593 11656 26372 11658
rect 10593 11600 10598 11656
rect 10654 11600 26372 11656
rect 10593 11598 26372 11600
rect 10593 11595 10659 11598
rect 26366 11596 26372 11598
rect 26436 11596 26442 11660
rect 28993 11658 29059 11661
rect 30281 11658 30347 11661
rect 32029 11658 32095 11661
rect 28993 11656 29194 11658
rect 28993 11600 28998 11656
rect 29054 11600 29194 11656
rect 28993 11598 29194 11600
rect 28993 11595 29059 11598
rect 14549 11522 14615 11525
rect 17585 11522 17651 11525
rect 14549 11520 17651 11522
rect 14549 11464 14554 11520
rect 14610 11464 17590 11520
rect 17646 11464 17651 11520
rect 14549 11462 17651 11464
rect 29134 11522 29194 11598
rect 30281 11656 32095 11658
rect 30281 11600 30286 11656
rect 30342 11600 32034 11656
rect 32090 11600 32095 11656
rect 30281 11598 32095 11600
rect 30281 11595 30347 11598
rect 32029 11595 32095 11598
rect 31017 11522 31083 11525
rect 29134 11520 31083 11522
rect 29134 11464 31022 11520
rect 31078 11464 31083 11520
rect 29134 11462 31083 11464
rect 14549 11459 14615 11462
rect 17585 11459 17651 11462
rect 31017 11459 31083 11462
rect 31385 11522 31451 11525
rect 32397 11522 32463 11525
rect 31385 11520 32463 11522
rect 31385 11464 31390 11520
rect 31446 11464 32402 11520
rect 32458 11464 32463 11520
rect 31385 11462 32463 11464
rect 31385 11459 31451 11462
rect 32397 11459 32463 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 16481 11386 16547 11389
rect 17677 11386 17743 11389
rect 16481 11384 17743 11386
rect 16481 11328 16486 11384
rect 16542 11328 17682 11384
rect 17738 11328 17743 11384
rect 16481 11326 17743 11328
rect 16481 11323 16547 11326
rect 17677 11323 17743 11326
rect 25630 11324 25636 11388
rect 25700 11386 25706 11388
rect 31661 11386 31727 11389
rect 25700 11384 31727 11386
rect 25700 11328 31666 11384
rect 31722 11328 31727 11384
rect 25700 11326 31727 11328
rect 25700 11324 25706 11326
rect 31661 11323 31727 11326
rect 17493 11250 17559 11253
rect 30414 11250 30420 11252
rect 17493 11248 30420 11250
rect 17493 11192 17498 11248
rect 17554 11192 30420 11248
rect 17493 11190 30420 11192
rect 17493 11187 17559 11190
rect 30414 11188 30420 11190
rect 30484 11250 30490 11252
rect 30833 11250 30899 11253
rect 30484 11248 30899 11250
rect 30484 11192 30838 11248
rect 30894 11192 30899 11248
rect 30484 11190 30899 11192
rect 30484 11188 30490 11190
rect 30833 11187 30899 11190
rect 31845 11250 31911 11253
rect 31845 11248 31954 11250
rect 31845 11192 31850 11248
rect 31906 11192 31954 11248
rect 31845 11187 31954 11192
rect 16665 11114 16731 11117
rect 17217 11114 17283 11117
rect 16665 11112 17283 11114
rect 16665 11056 16670 11112
rect 16726 11056 17222 11112
rect 17278 11056 17283 11112
rect 16665 11054 17283 11056
rect 16665 11051 16731 11054
rect 17217 11051 17283 11054
rect 20253 11114 20319 11117
rect 25681 11114 25747 11117
rect 20253 11112 25747 11114
rect 20253 11056 20258 11112
rect 20314 11056 25686 11112
rect 25742 11056 25747 11112
rect 20253 11054 25747 11056
rect 20253 11051 20319 11054
rect 25681 11051 25747 11054
rect 31894 10978 31954 11187
rect 32029 10978 32095 10981
rect 31894 10976 32095 10978
rect 31894 10920 32034 10976
rect 32090 10920 32095 10976
rect 31894 10918 32095 10920
rect 32029 10915 32095 10918
rect 32254 10916 32260 10980
rect 32324 10978 32330 10980
rect 32397 10978 32463 10981
rect 32324 10976 32463 10978
rect 32324 10920 32402 10976
rect 32458 10920 32463 10976
rect 32324 10918 32463 10920
rect 32324 10916 32330 10918
rect 32397 10915 32463 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 3325 10706 3391 10709
rect 5809 10706 5875 10709
rect 3325 10704 5875 10706
rect 3325 10648 3330 10704
rect 3386 10648 5814 10704
rect 5870 10648 5875 10704
rect 3325 10646 5875 10648
rect 3325 10643 3391 10646
rect 5809 10643 5875 10646
rect 14457 10706 14523 10709
rect 17769 10706 17835 10709
rect 14457 10704 17835 10706
rect 14457 10648 14462 10704
rect 14518 10648 17774 10704
rect 17830 10648 17835 10704
rect 14457 10646 17835 10648
rect 14457 10643 14523 10646
rect 17769 10643 17835 10646
rect 17953 10706 18019 10709
rect 20069 10706 20135 10709
rect 20897 10706 20963 10709
rect 17953 10704 20963 10706
rect 17953 10648 17958 10704
rect 18014 10648 20074 10704
rect 20130 10648 20902 10704
rect 20958 10648 20963 10704
rect 17953 10646 20963 10648
rect 17953 10643 18019 10646
rect 20069 10643 20135 10646
rect 20897 10643 20963 10646
rect 21357 10706 21423 10709
rect 22921 10706 22987 10709
rect 23054 10706 23060 10708
rect 21357 10704 23060 10706
rect 21357 10648 21362 10704
rect 21418 10648 22926 10704
rect 22982 10648 23060 10704
rect 21357 10646 23060 10648
rect 21357 10643 21423 10646
rect 22921 10643 22987 10646
rect 23054 10644 23060 10646
rect 23124 10644 23130 10708
rect 25313 10706 25379 10709
rect 25630 10706 25636 10708
rect 25313 10704 25636 10706
rect 25313 10648 25318 10704
rect 25374 10648 25636 10704
rect 25313 10646 25636 10648
rect 25313 10643 25379 10646
rect 25630 10644 25636 10646
rect 25700 10644 25706 10708
rect 18689 10570 18755 10573
rect 21541 10570 21607 10573
rect 18689 10568 21607 10570
rect 18689 10512 18694 10568
rect 18750 10512 21546 10568
rect 21602 10512 21607 10568
rect 18689 10510 21607 10512
rect 18689 10507 18755 10510
rect 21541 10507 21607 10510
rect 29085 10570 29151 10573
rect 31293 10570 31359 10573
rect 29085 10568 31359 10570
rect 29085 10512 29090 10568
rect 29146 10512 31298 10568
rect 31354 10512 31359 10568
rect 29085 10510 31359 10512
rect 29085 10507 29151 10510
rect 31293 10507 31359 10510
rect 19609 10434 19675 10437
rect 25037 10434 25103 10437
rect 25589 10434 25655 10437
rect 19609 10432 25655 10434
rect 19609 10376 19614 10432
rect 19670 10376 25042 10432
rect 25098 10376 25594 10432
rect 25650 10376 25655 10432
rect 19609 10374 25655 10376
rect 19609 10371 19675 10374
rect 25037 10371 25103 10374
rect 25589 10371 25655 10374
rect 30598 10372 30604 10436
rect 30668 10434 30674 10436
rect 31385 10434 31451 10437
rect 30668 10432 31451 10434
rect 30668 10376 31390 10432
rect 31446 10376 31451 10432
rect 30668 10374 31451 10376
rect 30668 10372 30674 10374
rect 31385 10371 31451 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 23105 10298 23171 10301
rect 24342 10298 24348 10300
rect 23105 10296 24348 10298
rect 23105 10240 23110 10296
rect 23166 10240 24348 10296
rect 23105 10238 24348 10240
rect 23105 10235 23171 10238
rect 24342 10236 24348 10238
rect 24412 10298 24418 10300
rect 24485 10298 24551 10301
rect 24412 10296 24551 10298
rect 24412 10240 24490 10296
rect 24546 10240 24551 10296
rect 24412 10238 24551 10240
rect 24412 10236 24418 10238
rect 24485 10235 24551 10238
rect 29494 10236 29500 10300
rect 29564 10298 29570 10300
rect 30189 10298 30255 10301
rect 31201 10300 31267 10301
rect 29564 10296 30255 10298
rect 29564 10240 30194 10296
rect 30250 10240 30255 10296
rect 29564 10238 30255 10240
rect 29564 10236 29570 10238
rect 30189 10235 30255 10238
rect 31150 10236 31156 10300
rect 31220 10298 31267 10300
rect 34278 10298 34284 10300
rect 31220 10296 31312 10298
rect 31262 10240 31312 10296
rect 31220 10238 31312 10240
rect 31710 10238 34284 10298
rect 31220 10236 31267 10238
rect 31201 10235 31267 10236
rect 3918 10100 3924 10164
rect 3988 10162 3994 10164
rect 4705 10162 4771 10165
rect 3988 10160 4771 10162
rect 3988 10104 4710 10160
rect 4766 10104 4771 10160
rect 3988 10102 4771 10104
rect 3988 10100 3994 10102
rect 4705 10099 4771 10102
rect 8293 10162 8359 10165
rect 8937 10162 9003 10165
rect 17401 10162 17467 10165
rect 8293 10160 17467 10162
rect 8293 10104 8298 10160
rect 8354 10104 8942 10160
rect 8998 10104 17406 10160
rect 17462 10104 17467 10160
rect 8293 10102 17467 10104
rect 8293 10099 8359 10102
rect 8937 10099 9003 10102
rect 17401 10099 17467 10102
rect 19885 10162 19951 10165
rect 21633 10162 21699 10165
rect 23473 10162 23539 10165
rect 19885 10160 23539 10162
rect 19885 10104 19890 10160
rect 19946 10104 21638 10160
rect 21694 10104 23478 10160
rect 23534 10104 23539 10160
rect 19885 10102 23539 10104
rect 19885 10099 19951 10102
rect 21633 10099 21699 10102
rect 23473 10099 23539 10102
rect 26233 10162 26299 10165
rect 31710 10162 31770 10238
rect 34278 10236 34284 10238
rect 34348 10298 34354 10300
rect 34421 10298 34487 10301
rect 34348 10296 34487 10298
rect 34348 10240 34426 10296
rect 34482 10240 34487 10296
rect 34348 10238 34487 10240
rect 34348 10236 34354 10238
rect 34421 10235 34487 10238
rect 26233 10160 31770 10162
rect 26233 10104 26238 10160
rect 26294 10104 31770 10160
rect 26233 10102 31770 10104
rect 26233 10099 26299 10102
rect 2221 10026 2287 10029
rect 4245 10026 4311 10029
rect 32489 10028 32555 10029
rect 32438 10026 32444 10028
rect 2221 10024 4311 10026
rect 2221 9968 2226 10024
rect 2282 9968 4250 10024
rect 4306 9968 4311 10024
rect 2221 9966 4311 9968
rect 32398 9966 32444 10026
rect 32508 10024 32555 10028
rect 32550 9968 32555 10024
rect 2221 9963 2287 9966
rect 3880 9893 3940 9966
rect 4245 9963 4311 9966
rect 32438 9964 32444 9966
rect 32508 9964 32555 9968
rect 32489 9963 32555 9964
rect 3877 9888 3943 9893
rect 3877 9832 3882 9888
rect 3938 9832 3943 9888
rect 3877 9827 3943 9832
rect 29177 9890 29243 9893
rect 35341 9890 35407 9893
rect 29177 9888 35407 9890
rect 29177 9832 29182 9888
rect 29238 9832 35346 9888
rect 35402 9832 35407 9888
rect 29177 9830 35407 9832
rect 29177 9827 29243 9830
rect 35341 9827 35407 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 18505 9754 18571 9757
rect 25405 9754 25471 9757
rect 28993 9754 29059 9757
rect 29821 9754 29887 9757
rect 18505 9752 29887 9754
rect 18505 9696 18510 9752
rect 18566 9696 25410 9752
rect 25466 9696 28998 9752
rect 29054 9696 29826 9752
rect 29882 9696 29887 9752
rect 18505 9694 29887 9696
rect 18505 9691 18571 9694
rect 25405 9691 25471 9694
rect 28993 9691 29059 9694
rect 29821 9691 29887 9694
rect 33133 9754 33199 9757
rect 34094 9754 34100 9756
rect 33133 9752 34100 9754
rect 33133 9696 33138 9752
rect 33194 9696 34100 9752
rect 33133 9694 34100 9696
rect 33133 9691 33199 9694
rect 34094 9692 34100 9694
rect 34164 9754 34170 9756
rect 34237 9754 34303 9757
rect 34164 9752 34303 9754
rect 34164 9696 34242 9752
rect 34298 9696 34303 9752
rect 34164 9694 34303 9696
rect 34164 9692 34170 9694
rect 34237 9691 34303 9694
rect 4981 9618 5047 9621
rect 5441 9618 5507 9621
rect 5574 9618 5580 9620
rect 4981 9616 5580 9618
rect 4981 9560 4986 9616
rect 5042 9560 5446 9616
rect 5502 9560 5580 9616
rect 4981 9558 5580 9560
rect 4981 9555 5047 9558
rect 5441 9555 5507 9558
rect 5574 9556 5580 9558
rect 5644 9556 5650 9620
rect 7373 9618 7439 9621
rect 8845 9618 8911 9621
rect 7373 9616 8911 9618
rect 7373 9560 7378 9616
rect 7434 9560 8850 9616
rect 8906 9560 8911 9616
rect 7373 9558 8911 9560
rect 7373 9555 7439 9558
rect 8845 9555 8911 9558
rect 19558 9556 19564 9620
rect 19628 9618 19634 9620
rect 20069 9618 20135 9621
rect 26233 9618 26299 9621
rect 26785 9618 26851 9621
rect 19628 9616 20135 9618
rect 19628 9560 20074 9616
rect 20130 9560 20135 9616
rect 19628 9558 20135 9560
rect 19628 9556 19634 9558
rect 20069 9555 20135 9558
rect 22050 9616 26851 9618
rect 22050 9560 26238 9616
rect 26294 9560 26790 9616
rect 26846 9560 26851 9616
rect 22050 9558 26851 9560
rect 12525 9482 12591 9485
rect 12750 9482 12756 9484
rect 12525 9480 12756 9482
rect 12525 9424 12530 9480
rect 12586 9424 12756 9480
rect 12525 9422 12756 9424
rect 12525 9419 12591 9422
rect 12750 9420 12756 9422
rect 12820 9420 12826 9484
rect 20805 9482 20871 9485
rect 22050 9482 22110 9558
rect 26233 9555 26299 9558
rect 26785 9555 26851 9558
rect 28257 9618 28323 9621
rect 33501 9618 33567 9621
rect 28257 9616 33567 9618
rect 28257 9560 28262 9616
rect 28318 9560 33506 9616
rect 33562 9560 33567 9616
rect 28257 9558 33567 9560
rect 28257 9555 28323 9558
rect 33501 9555 33567 9558
rect 34053 9618 34119 9621
rect 35157 9618 35223 9621
rect 34053 9616 35223 9618
rect 34053 9560 34058 9616
rect 34114 9560 35162 9616
rect 35218 9560 35223 9616
rect 34053 9558 35223 9560
rect 34053 9555 34119 9558
rect 35157 9555 35223 9558
rect 20805 9480 22110 9482
rect 20805 9424 20810 9480
rect 20866 9424 22110 9480
rect 20805 9422 22110 9424
rect 22277 9482 22343 9485
rect 24025 9482 24091 9485
rect 24301 9482 24367 9485
rect 22277 9480 24367 9482
rect 22277 9424 22282 9480
rect 22338 9424 24030 9480
rect 24086 9424 24306 9480
rect 24362 9424 24367 9480
rect 22277 9422 24367 9424
rect 20805 9419 20871 9422
rect 22277 9419 22343 9422
rect 24025 9419 24091 9422
rect 24301 9419 24367 9422
rect 26049 9482 26115 9485
rect 31385 9482 31451 9485
rect 26049 9480 31451 9482
rect 26049 9424 26054 9480
rect 26110 9424 31390 9480
rect 31446 9424 31451 9480
rect 26049 9422 31451 9424
rect 26049 9419 26115 9422
rect 31385 9419 31451 9422
rect 31661 9482 31727 9485
rect 32489 9482 32555 9485
rect 34973 9482 35039 9485
rect 35525 9482 35591 9485
rect 31661 9480 35591 9482
rect 31661 9424 31666 9480
rect 31722 9424 32494 9480
rect 32550 9424 34978 9480
rect 35034 9424 35530 9480
rect 35586 9424 35591 9480
rect 31661 9422 35591 9424
rect 31661 9419 31727 9422
rect 32489 9419 32555 9422
rect 34973 9419 35039 9422
rect 35525 9419 35591 9422
rect 7005 9346 7071 9349
rect 8753 9346 8819 9349
rect 7005 9344 8819 9346
rect 7005 9288 7010 9344
rect 7066 9288 8758 9344
rect 8814 9288 8819 9344
rect 7005 9286 8819 9288
rect 7005 9283 7071 9286
rect 8753 9283 8819 9286
rect 23381 9346 23447 9349
rect 26785 9346 26851 9349
rect 30833 9346 30899 9349
rect 23381 9344 30899 9346
rect 23381 9288 23386 9344
rect 23442 9288 26790 9344
rect 26846 9288 30838 9344
rect 30894 9288 30899 9344
rect 23381 9286 30899 9288
rect 23381 9283 23447 9286
rect 26785 9283 26851 9286
rect 30833 9283 30899 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4889 9210 4955 9213
rect 9029 9210 9095 9213
rect 4889 9208 9095 9210
rect 4889 9152 4894 9208
rect 4950 9152 9034 9208
rect 9090 9152 9095 9208
rect 4889 9150 9095 9152
rect 4889 9147 4955 9150
rect 9029 9147 9095 9150
rect 17585 9210 17651 9213
rect 17902 9210 17908 9212
rect 17585 9208 17908 9210
rect 17585 9152 17590 9208
rect 17646 9152 17908 9208
rect 17585 9150 17908 9152
rect 17585 9147 17651 9150
rect 17902 9148 17908 9150
rect 17972 9148 17978 9212
rect 18965 9210 19031 9213
rect 24393 9210 24459 9213
rect 18965 9208 24459 9210
rect 18965 9152 18970 9208
rect 19026 9152 24398 9208
rect 24454 9152 24459 9208
rect 18965 9150 24459 9152
rect 18965 9147 19031 9150
rect 24393 9147 24459 9150
rect 26141 9212 26207 9213
rect 26141 9208 26188 9212
rect 26252 9210 26258 9212
rect 26141 9152 26146 9208
rect 26141 9148 26188 9152
rect 26252 9150 26298 9210
rect 26252 9148 26258 9150
rect 26141 9147 26207 9148
rect 3693 9074 3759 9077
rect 4889 9074 4955 9077
rect 3693 9072 4955 9074
rect 3693 9016 3698 9072
rect 3754 9016 4894 9072
rect 4950 9016 4955 9072
rect 3693 9014 4955 9016
rect 3693 9011 3759 9014
rect 4889 9011 4955 9014
rect 5625 9074 5691 9077
rect 5758 9074 5764 9076
rect 5625 9072 5764 9074
rect 5625 9016 5630 9072
rect 5686 9016 5764 9072
rect 5625 9014 5764 9016
rect 5625 9011 5691 9014
rect 5758 9012 5764 9014
rect 5828 9012 5834 9076
rect 13813 9074 13879 9077
rect 26877 9074 26943 9077
rect 27337 9074 27403 9077
rect 13813 9072 27403 9074
rect 13813 9016 13818 9072
rect 13874 9016 26882 9072
rect 26938 9016 27342 9072
rect 27398 9016 27403 9072
rect 13813 9014 27403 9016
rect 13813 9011 13879 9014
rect 26877 9011 26943 9014
rect 27337 9011 27403 9014
rect 4705 8940 4771 8941
rect 4654 8876 4660 8940
rect 4724 8938 4771 8940
rect 18229 8938 18295 8941
rect 19241 8938 19307 8941
rect 4724 8936 4816 8938
rect 4766 8880 4816 8936
rect 4724 8878 4816 8880
rect 18229 8936 19307 8938
rect 18229 8880 18234 8936
rect 18290 8880 19246 8936
rect 19302 8880 19307 8936
rect 18229 8878 19307 8880
rect 4724 8876 4771 8878
rect 4705 8875 4771 8876
rect 18229 8875 18295 8878
rect 19241 8875 19307 8878
rect 24301 8938 24367 8941
rect 27061 8938 27127 8941
rect 28717 8938 28783 8941
rect 24301 8936 28783 8938
rect 24301 8880 24306 8936
rect 24362 8880 27066 8936
rect 27122 8880 28722 8936
rect 28778 8880 28783 8936
rect 24301 8878 28783 8880
rect 24301 8875 24367 8878
rect 27061 8875 27127 8878
rect 28717 8875 28783 8878
rect 8201 8802 8267 8805
rect 26693 8802 26759 8805
rect 8201 8800 26759 8802
rect 8201 8744 8206 8800
rect 8262 8744 26698 8800
rect 26754 8744 26759 8800
rect 8201 8742 26759 8744
rect 8201 8739 8267 8742
rect 26693 8739 26759 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 6678 8604 6684 8668
rect 6748 8666 6754 8668
rect 7741 8666 7807 8669
rect 32949 8668 33015 8669
rect 32949 8666 32996 8668
rect 6748 8664 7807 8666
rect 6748 8608 7746 8664
rect 7802 8608 7807 8664
rect 6748 8606 7807 8608
rect 32904 8664 32996 8666
rect 32904 8608 32954 8664
rect 32904 8606 32996 8608
rect 6748 8604 6754 8606
rect 7741 8603 7807 8606
rect 32949 8604 32996 8606
rect 33060 8604 33066 8668
rect 32949 8603 33015 8604
rect 4889 8530 4955 8533
rect 9673 8532 9739 8533
rect 5390 8530 5396 8532
rect 4889 8528 5396 8530
rect 4889 8472 4894 8528
rect 4950 8472 5396 8528
rect 4889 8470 5396 8472
rect 4889 8467 4955 8470
rect 5390 8468 5396 8470
rect 5460 8468 5466 8532
rect 9622 8468 9628 8532
rect 9692 8530 9739 8532
rect 20253 8530 20319 8533
rect 21357 8530 21423 8533
rect 9692 8528 9784 8530
rect 9734 8472 9784 8528
rect 9692 8470 9784 8472
rect 20253 8528 21423 8530
rect 20253 8472 20258 8528
rect 20314 8472 21362 8528
rect 21418 8472 21423 8528
rect 20253 8470 21423 8472
rect 9692 8468 9739 8470
rect 9673 8467 9739 8468
rect 20253 8467 20319 8470
rect 21357 8467 21423 8470
rect 23565 8530 23631 8533
rect 26693 8530 26759 8533
rect 23565 8528 26759 8530
rect 23565 8472 23570 8528
rect 23626 8472 26698 8528
rect 26754 8472 26759 8528
rect 23565 8470 26759 8472
rect 23565 8467 23631 8470
rect 26693 8467 26759 8470
rect 29269 8530 29335 8533
rect 30925 8530 30991 8533
rect 29269 8528 30991 8530
rect 29269 8472 29274 8528
rect 29330 8472 30930 8528
rect 30986 8472 30991 8528
rect 29269 8470 30991 8472
rect 29269 8467 29335 8470
rect 30925 8467 30991 8470
rect 4429 8394 4495 8397
rect 11053 8396 11119 8397
rect 11053 8394 11100 8396
rect 4429 8392 11100 8394
rect 4429 8336 4434 8392
rect 4490 8336 11058 8392
rect 4429 8334 11100 8336
rect 4429 8331 4495 8334
rect 11053 8332 11100 8334
rect 11164 8332 11170 8396
rect 16389 8394 16455 8397
rect 19057 8394 19123 8397
rect 16389 8392 19123 8394
rect 16389 8336 16394 8392
rect 16450 8336 19062 8392
rect 19118 8336 19123 8392
rect 16389 8334 19123 8336
rect 11053 8331 11119 8332
rect 16389 8331 16455 8334
rect 19057 8331 19123 8334
rect 30833 8394 30899 8397
rect 32305 8394 32371 8397
rect 30833 8392 32371 8394
rect 30833 8336 30838 8392
rect 30894 8336 32310 8392
rect 32366 8336 32371 8392
rect 30833 8334 32371 8336
rect 30833 8331 30899 8334
rect 32305 8331 32371 8334
rect 25497 8258 25563 8261
rect 26366 8258 26372 8260
rect 25497 8256 26372 8258
rect 25497 8200 25502 8256
rect 25558 8200 26372 8256
rect 25497 8198 26372 8200
rect 25497 8195 25563 8198
rect 26366 8196 26372 8198
rect 26436 8258 26442 8260
rect 26969 8258 27035 8261
rect 26436 8256 27035 8258
rect 26436 8200 26974 8256
rect 27030 8200 27035 8256
rect 26436 8198 27035 8200
rect 26436 8196 26442 8198
rect 26969 8195 27035 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 14181 7988 14247 7989
rect 14181 7986 14228 7988
rect 14136 7984 14228 7986
rect 14136 7928 14186 7984
rect 14136 7926 14228 7928
rect 14181 7924 14228 7926
rect 14292 7924 14298 7988
rect 21081 7986 21147 7989
rect 26049 7986 26115 7989
rect 26785 7986 26851 7989
rect 21081 7984 22110 7986
rect 21081 7928 21086 7984
rect 21142 7928 22110 7984
rect 21081 7926 22110 7928
rect 14181 7923 14247 7924
rect 21081 7923 21147 7926
rect 19057 7850 19123 7853
rect 21173 7850 21239 7853
rect 19057 7848 21239 7850
rect 19057 7792 19062 7848
rect 19118 7792 21178 7848
rect 21234 7792 21239 7848
rect 19057 7790 21239 7792
rect 19057 7787 19123 7790
rect 21173 7787 21239 7790
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 8334 7516 8340 7580
rect 8404 7578 8410 7580
rect 8753 7578 8819 7581
rect 8404 7576 8819 7578
rect 8404 7520 8758 7576
rect 8814 7520 8819 7576
rect 8404 7518 8819 7520
rect 22050 7578 22110 7926
rect 26049 7984 26851 7986
rect 26049 7928 26054 7984
rect 26110 7928 26790 7984
rect 26846 7928 26851 7984
rect 26049 7926 26851 7928
rect 26049 7923 26115 7926
rect 26785 7923 26851 7926
rect 27797 7986 27863 7989
rect 28533 7988 28599 7989
rect 28022 7986 28028 7988
rect 27797 7984 28028 7986
rect 27797 7928 27802 7984
rect 27858 7928 28028 7984
rect 27797 7926 28028 7928
rect 27797 7923 27863 7926
rect 28022 7924 28028 7926
rect 28092 7924 28098 7988
rect 28533 7986 28580 7988
rect 28488 7984 28580 7986
rect 28488 7928 28538 7984
rect 28488 7926 28580 7928
rect 28533 7924 28580 7926
rect 28644 7924 28650 7988
rect 28533 7923 28599 7924
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 33041 7578 33107 7581
rect 33542 7578 33548 7580
rect 22050 7576 33548 7578
rect 22050 7520 33046 7576
rect 33102 7520 33548 7576
rect 22050 7518 33548 7520
rect 8404 7516 8410 7518
rect 8753 7515 8819 7518
rect 33041 7515 33107 7518
rect 33542 7516 33548 7518
rect 33612 7516 33618 7580
rect 4797 7442 4863 7445
rect 8661 7442 8727 7445
rect 4797 7440 8727 7442
rect 4797 7384 4802 7440
rect 4858 7384 8666 7440
rect 8722 7384 8727 7440
rect 4797 7382 8727 7384
rect 4797 7379 4863 7382
rect 8661 7379 8727 7382
rect 12249 7442 12315 7445
rect 28533 7442 28599 7445
rect 12249 7440 28599 7442
rect 12249 7384 12254 7440
rect 12310 7384 28538 7440
rect 28594 7384 28599 7440
rect 12249 7382 28599 7384
rect 12249 7379 12315 7382
rect 28533 7379 28599 7382
rect 5993 7306 6059 7309
rect 9029 7306 9095 7309
rect 5993 7304 9095 7306
rect 5993 7248 5998 7304
rect 6054 7248 9034 7304
rect 9090 7248 9095 7304
rect 5993 7246 9095 7248
rect 5993 7243 6059 7246
rect 9029 7243 9095 7246
rect 11789 7306 11855 7309
rect 13813 7306 13879 7309
rect 11789 7304 13879 7306
rect 11789 7248 11794 7304
rect 11850 7248 13818 7304
rect 13874 7248 13879 7304
rect 11789 7246 13879 7248
rect 11789 7243 11855 7246
rect 13813 7243 13879 7246
rect 16481 7306 16547 7309
rect 18965 7306 19031 7309
rect 16481 7304 19031 7306
rect 16481 7248 16486 7304
rect 16542 7248 18970 7304
rect 19026 7248 19031 7304
rect 16481 7246 19031 7248
rect 16481 7243 16547 7246
rect 18965 7243 19031 7246
rect 24945 7306 25011 7309
rect 29126 7306 29132 7308
rect 24945 7304 29132 7306
rect 24945 7248 24950 7304
rect 25006 7248 29132 7304
rect 24945 7246 29132 7248
rect 24945 7243 25011 7246
rect 29126 7244 29132 7246
rect 29196 7244 29202 7308
rect 21633 7170 21699 7173
rect 23974 7170 23980 7172
rect 21633 7168 23980 7170
rect 21633 7112 21638 7168
rect 21694 7112 23980 7168
rect 21633 7110 23980 7112
rect 21633 7107 21699 7110
rect 23974 7108 23980 7110
rect 24044 7170 24050 7172
rect 28165 7170 28231 7173
rect 24044 7168 28231 7170
rect 24044 7112 28170 7168
rect 28226 7112 28231 7168
rect 24044 7110 28231 7112
rect 24044 7108 24050 7110
rect 28165 7107 28231 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 3509 6898 3575 6901
rect 6545 6898 6611 6901
rect 3509 6896 6611 6898
rect 3509 6840 3514 6896
rect 3570 6840 6550 6896
rect 6606 6840 6611 6896
rect 3509 6838 6611 6840
rect 3509 6835 3575 6838
rect 6545 6835 6611 6838
rect 7230 6836 7236 6900
rect 7300 6898 7306 6900
rect 8569 6898 8635 6901
rect 7300 6896 8635 6898
rect 7300 6840 8574 6896
rect 8630 6840 8635 6896
rect 7300 6838 8635 6840
rect 7300 6836 7306 6838
rect 8569 6835 8635 6838
rect 9213 6900 9279 6901
rect 9213 6896 9260 6900
rect 9324 6898 9330 6900
rect 11513 6898 11579 6901
rect 11646 6898 11652 6900
rect 9213 6840 9218 6896
rect 9213 6836 9260 6840
rect 9324 6838 9370 6898
rect 11513 6896 11652 6898
rect 11513 6840 11518 6896
rect 11574 6840 11652 6896
rect 11513 6838 11652 6840
rect 9324 6836 9330 6838
rect 9213 6835 9279 6836
rect 11513 6835 11579 6838
rect 11646 6836 11652 6838
rect 11716 6836 11722 6900
rect 15193 6898 15259 6901
rect 15326 6898 15332 6900
rect 15193 6896 15332 6898
rect 15193 6840 15198 6896
rect 15254 6840 15332 6896
rect 15193 6838 15332 6840
rect 15193 6835 15259 6838
rect 15326 6836 15332 6838
rect 15396 6836 15402 6900
rect 21214 6836 21220 6900
rect 21284 6898 21290 6900
rect 21541 6898 21607 6901
rect 21284 6896 21607 6898
rect 21284 6840 21546 6896
rect 21602 6840 21607 6896
rect 21284 6838 21607 6840
rect 21284 6836 21290 6838
rect 21541 6835 21607 6838
rect 22829 6900 22895 6901
rect 22829 6896 22876 6900
rect 22940 6898 22946 6900
rect 22829 6840 22834 6896
rect 22829 6836 22876 6840
rect 22940 6838 22986 6898
rect 22940 6836 22946 6838
rect 22829 6835 22895 6836
rect 3969 6762 4035 6765
rect 7741 6762 7807 6765
rect 3969 6760 7807 6762
rect 3969 6704 3974 6760
rect 4030 6704 7746 6760
rect 7802 6704 7807 6760
rect 3969 6702 7807 6704
rect 3969 6699 4035 6702
rect 7741 6699 7807 6702
rect 18505 6762 18571 6765
rect 18873 6762 18939 6765
rect 18505 6760 18939 6762
rect 18505 6704 18510 6760
rect 18566 6704 18878 6760
rect 18934 6704 18939 6760
rect 18505 6702 18939 6704
rect 18505 6699 18571 6702
rect 18873 6699 18939 6702
rect 19977 6762 20043 6765
rect 27797 6762 27863 6765
rect 19977 6760 27863 6762
rect 19977 6704 19982 6760
rect 20038 6704 27802 6760
rect 27858 6704 27863 6760
rect 19977 6702 27863 6704
rect 19977 6699 20043 6702
rect 27797 6699 27863 6702
rect 6729 6626 6795 6629
rect 7465 6626 7531 6629
rect 6729 6624 7531 6626
rect 6729 6568 6734 6624
rect 6790 6568 7470 6624
rect 7526 6568 7531 6624
rect 6729 6566 7531 6568
rect 6729 6563 6795 6566
rect 7465 6563 7531 6566
rect 11605 6626 11671 6629
rect 13629 6626 13695 6629
rect 11605 6624 13695 6626
rect 11605 6568 11610 6624
rect 11666 6568 13634 6624
rect 13690 6568 13695 6624
rect 11605 6566 13695 6568
rect 11605 6563 11671 6566
rect 13629 6563 13695 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 11513 6492 11579 6493
rect 11462 6428 11468 6492
rect 11532 6490 11579 6492
rect 11532 6488 11624 6490
rect 11574 6432 11624 6488
rect 11532 6430 11624 6432
rect 11532 6428 11579 6430
rect 17534 6428 17540 6492
rect 17604 6490 17610 6492
rect 17677 6490 17743 6493
rect 17604 6488 17743 6490
rect 17604 6432 17682 6488
rect 17738 6432 17743 6488
rect 17604 6430 17743 6432
rect 17604 6428 17610 6430
rect 11513 6427 11579 6428
rect 17677 6427 17743 6430
rect 13813 6354 13879 6357
rect 27521 6354 27587 6357
rect 13813 6352 27587 6354
rect 13813 6296 13818 6352
rect 13874 6296 27526 6352
rect 27582 6296 27587 6352
rect 13813 6294 27587 6296
rect 13813 6291 13879 6294
rect 27521 6291 27587 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 31937 5946 32003 5949
rect 32070 5946 32076 5948
rect 31937 5944 32076 5946
rect 31937 5888 31942 5944
rect 31998 5888 32076 5944
rect 31937 5886 32076 5888
rect 31937 5883 32003 5886
rect 32070 5884 32076 5886
rect 32140 5884 32146 5948
rect 12893 5674 12959 5677
rect 13537 5676 13603 5677
rect 13486 5674 13492 5676
rect 12893 5672 13492 5674
rect 13556 5674 13603 5676
rect 26049 5674 26115 5677
rect 13556 5672 26115 5674
rect 12893 5616 12898 5672
rect 12954 5616 13492 5672
rect 13598 5616 26054 5672
rect 26110 5616 26115 5672
rect 12893 5614 13492 5616
rect 12893 5611 12959 5614
rect 13486 5612 13492 5614
rect 13556 5614 26115 5616
rect 13556 5612 13603 5614
rect 13537 5611 13603 5612
rect 26049 5611 26115 5614
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 21398 5340 21404 5404
rect 21468 5402 21474 5404
rect 21541 5402 21607 5405
rect 22001 5402 22067 5405
rect 21468 5400 22067 5402
rect 21468 5344 21546 5400
rect 21602 5344 22006 5400
rect 22062 5344 22067 5400
rect 21468 5342 22067 5344
rect 21468 5340 21474 5342
rect 21541 5339 21607 5342
rect 22001 5339 22067 5342
rect 17493 5266 17559 5269
rect 18638 5266 18644 5268
rect 17493 5264 18644 5266
rect 17493 5208 17498 5264
rect 17554 5208 18644 5264
rect 17493 5206 18644 5208
rect 17493 5203 17559 5206
rect 18638 5204 18644 5206
rect 18708 5204 18714 5268
rect 19742 5068 19748 5132
rect 19812 5130 19818 5132
rect 21081 5130 21147 5133
rect 30373 5132 30439 5133
rect 30373 5130 30420 5132
rect 19812 5128 21147 5130
rect 19812 5072 21086 5128
rect 21142 5072 21147 5128
rect 19812 5070 21147 5072
rect 30328 5128 30420 5130
rect 30328 5072 30378 5128
rect 30328 5070 30420 5072
rect 19812 5068 19818 5070
rect 21081 5067 21147 5070
rect 30373 5068 30420 5070
rect 30484 5068 30490 5132
rect 30373 5067 30439 5068
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 21950 4524 21956 4588
rect 22020 4586 22026 4588
rect 23841 4586 23907 4589
rect 22020 4584 23907 4586
rect 22020 4528 23846 4584
rect 23902 4528 23907 4584
rect 22020 4526 23907 4528
rect 22020 4524 22026 4526
rect 23841 4523 23907 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 18413 4316 18479 4317
rect 18413 4314 18460 4316
rect 18368 4312 18460 4314
rect 18368 4256 18418 4312
rect 18368 4254 18460 4256
rect 18413 4252 18460 4254
rect 18524 4252 18530 4316
rect 18413 4251 18479 4252
rect 15837 4178 15903 4181
rect 16246 4178 16252 4180
rect 15837 4176 16252 4178
rect 15837 4120 15842 4176
rect 15898 4120 16252 4176
rect 15837 4118 16252 4120
rect 15837 4115 15903 4118
rect 16246 4116 16252 4118
rect 16316 4116 16322 4180
rect 20989 4178 21055 4181
rect 23565 4178 23631 4181
rect 20989 4176 23631 4178
rect 20989 4120 20994 4176
rect 21050 4120 23570 4176
rect 23626 4120 23631 4176
rect 20989 4118 23631 4120
rect 20989 4115 21055 4118
rect 23565 4115 23631 4118
rect 11145 4044 11211 4045
rect 11094 4042 11100 4044
rect 11054 3982 11100 4042
rect 11164 4042 11211 4044
rect 18597 4042 18663 4045
rect 11164 4040 18663 4042
rect 11206 3984 18602 4040
rect 18658 3984 18663 4040
rect 11094 3980 11100 3982
rect 11164 3982 18663 3984
rect 11164 3980 11211 3982
rect 11145 3979 11211 3980
rect 18597 3979 18663 3982
rect 22185 4042 22251 4045
rect 22686 4042 22692 4044
rect 22185 4040 22692 4042
rect 22185 3984 22190 4040
rect 22246 3984 22692 4040
rect 22185 3982 22692 3984
rect 22185 3979 22251 3982
rect 22686 3980 22692 3982
rect 22756 3980 22762 4044
rect 23933 4042 23999 4045
rect 24894 4042 24900 4044
rect 23933 4040 24900 4042
rect 23933 3984 23938 4040
rect 23994 3984 24900 4040
rect 23933 3982 24900 3984
rect 23933 3979 23999 3982
rect 24894 3980 24900 3982
rect 24964 3980 24970 4044
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 21081 3636 21147 3637
rect 21030 3572 21036 3636
rect 21100 3634 21147 3636
rect 21100 3632 21192 3634
rect 21142 3576 21192 3632
rect 21100 3574 21192 3576
rect 21100 3572 21147 3574
rect 21081 3571 21147 3572
rect 36077 3498 36143 3501
rect 36782 3498 37582 3528
rect 36077 3496 37582 3498
rect 36077 3440 36082 3496
rect 36138 3440 37582 3496
rect 36077 3438 37582 3440
rect 36077 3435 36143 3438
rect 36782 3408 37582 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 20437 3228 20503 3229
rect 20437 3226 20484 3228
rect 20392 3224 20484 3226
rect 20548 3226 20554 3228
rect 21909 3226 21975 3229
rect 22277 3226 22343 3229
rect 20548 3224 22343 3226
rect 20392 3168 20442 3224
rect 20548 3168 21914 3224
rect 21970 3168 22282 3224
rect 22338 3168 22343 3224
rect 20392 3166 20484 3168
rect 20437 3164 20484 3166
rect 20548 3166 22343 3168
rect 20548 3164 20554 3166
rect 20437 3163 20503 3164
rect 21909 3163 21975 3166
rect 22277 3163 22343 3166
rect 14590 3028 14596 3092
rect 14660 3090 14666 3092
rect 16389 3090 16455 3093
rect 14660 3088 16455 3090
rect 14660 3032 16394 3088
rect 16450 3032 16455 3088
rect 14660 3030 16455 3032
rect 14660 3028 14666 3030
rect 16389 3027 16455 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 20300 34852 20364 34916
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 9628 33084 9692 33148
rect 4660 32948 4724 33012
rect 10916 32948 10980 33012
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4660 32268 4724 32332
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 13308 31996 13372 32060
rect 26372 32056 26436 32060
rect 26372 32000 26422 32056
rect 26422 32000 26436 32056
rect 26372 31996 26436 32000
rect 15516 31860 15580 31924
rect 5580 31724 5644 31788
rect 14964 31724 15028 31788
rect 27476 31724 27540 31788
rect 27660 31784 27724 31788
rect 27660 31728 27674 31784
rect 27674 31728 27724 31784
rect 27660 31724 27724 31728
rect 5580 31588 5644 31652
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 28212 31648 28276 31652
rect 28212 31592 28262 31648
rect 28262 31592 28276 31648
rect 28212 31588 28276 31592
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 27292 31512 27356 31516
rect 27292 31456 27306 31512
rect 27306 31456 27356 31512
rect 27292 31452 27356 31456
rect 15332 31240 15396 31244
rect 15332 31184 15382 31240
rect 15382 31184 15396 31240
rect 15332 31180 15396 31184
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 6316 30364 6380 30428
rect 9628 30228 9692 30292
rect 13124 30288 13188 30292
rect 13124 30232 13138 30288
rect 13138 30232 13188 30288
rect 13124 30228 13188 30232
rect 9076 30092 9140 30156
rect 12204 30092 12268 30156
rect 23796 30152 23860 30156
rect 23796 30096 23810 30152
rect 23810 30096 23860 30152
rect 23796 30092 23860 30096
rect 27476 30092 27540 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 26188 29684 26252 29748
rect 28212 29684 28276 29748
rect 24164 29548 24228 29612
rect 30972 29548 31036 29612
rect 9996 29412 10060 29476
rect 25268 29472 25332 29476
rect 25268 29416 25282 29472
rect 25282 29416 25332 29472
rect 25268 29412 25332 29416
rect 27292 29472 27356 29476
rect 27292 29416 27342 29472
rect 27342 29416 27356 29472
rect 27292 29412 27356 29416
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 11100 29140 11164 29204
rect 14044 29200 14108 29204
rect 14044 29144 14058 29200
rect 14058 29144 14108 29200
rect 14044 29140 14108 29144
rect 13860 29004 13924 29068
rect 15148 29004 15212 29068
rect 19196 29004 19260 29068
rect 30052 29064 30116 29068
rect 30052 29008 30066 29064
rect 30066 29008 30116 29064
rect 30052 29004 30116 29008
rect 33548 29004 33612 29068
rect 34284 29004 34348 29068
rect 27660 28868 27724 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 10916 28732 10980 28796
rect 27660 28732 27724 28796
rect 29132 28596 29196 28660
rect 15700 28460 15764 28524
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 26372 28188 26436 28252
rect 26004 28052 26068 28116
rect 12756 27840 12820 27844
rect 27660 27916 27724 27980
rect 12756 27784 12806 27840
rect 12806 27784 12820 27840
rect 12756 27780 12820 27784
rect 22876 27840 22940 27844
rect 22876 27784 22890 27840
rect 22890 27784 22940 27840
rect 22876 27780 22940 27784
rect 30420 27780 30484 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 18460 27644 18524 27708
rect 9812 27508 9876 27572
rect 26188 27508 26252 27572
rect 27292 27704 27356 27708
rect 27292 27648 27342 27704
rect 27342 27648 27356 27704
rect 27292 27644 27356 27648
rect 30972 27568 31036 27572
rect 30972 27512 31022 27568
rect 31022 27512 31036 27568
rect 30972 27508 31036 27512
rect 5764 27236 5828 27300
rect 7604 27236 7668 27300
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 31524 26828 31588 26892
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 21404 26556 21468 26620
rect 22140 26420 22204 26484
rect 8340 26344 8404 26348
rect 8340 26288 8390 26344
rect 8390 26288 8404 26344
rect 8340 26284 8404 26288
rect 16620 26284 16684 26348
rect 17172 26284 17236 26348
rect 17908 26284 17972 26348
rect 21036 26284 21100 26348
rect 22692 26284 22756 26348
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 32260 25936 32324 25940
rect 32260 25880 32310 25936
rect 32310 25880 32324 25936
rect 32260 25876 32324 25880
rect 24164 25740 24228 25804
rect 7788 25664 7852 25668
rect 7788 25608 7838 25664
rect 7838 25608 7852 25664
rect 7788 25604 7852 25608
rect 29316 25664 29380 25668
rect 29316 25608 29366 25664
rect 29366 25608 29380 25664
rect 29316 25604 29380 25608
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 5948 25060 6012 25124
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 18276 24924 18340 24988
rect 14044 24788 14108 24852
rect 12756 24516 12820 24580
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 12940 24380 13004 24444
rect 16804 24380 16868 24444
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 11100 24244 11164 24308
rect 13124 24304 13188 24308
rect 13124 24248 13138 24304
rect 13138 24248 13188 24304
rect 13124 24244 13188 24248
rect 20852 24168 20916 24172
rect 20852 24112 20866 24168
rect 20866 24112 20916 24168
rect 20852 24108 20916 24112
rect 27476 24168 27540 24172
rect 27476 24112 27526 24168
rect 27526 24112 27540 24168
rect 27476 24108 27540 24112
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 23612 23836 23676 23900
rect 14596 23700 14660 23764
rect 21220 23700 21284 23764
rect 30788 23700 30852 23764
rect 11468 23564 11532 23628
rect 14228 23564 14292 23628
rect 9628 23488 9692 23492
rect 9628 23432 9642 23488
rect 9642 23432 9692 23488
rect 9628 23428 9692 23432
rect 13492 23428 13556 23492
rect 31156 23428 31220 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 16988 23352 17052 23356
rect 16988 23296 17038 23352
rect 17038 23296 17052 23352
rect 16988 23292 17052 23296
rect 2636 23020 2700 23084
rect 16804 23020 16868 23084
rect 3924 22884 3988 22948
rect 6316 22944 6380 22948
rect 6316 22888 6366 22944
rect 6366 22888 6380 22944
rect 6316 22884 6380 22888
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 19196 22748 19260 22812
rect 29500 22748 29564 22812
rect 25452 22672 25516 22676
rect 25452 22616 25466 22672
rect 25466 22616 25516 22672
rect 25452 22612 25516 22616
rect 9076 22536 9140 22540
rect 9076 22480 9126 22536
rect 9126 22480 9140 22536
rect 9076 22476 9140 22480
rect 21588 22476 21652 22540
rect 28212 22536 28276 22540
rect 28212 22480 28226 22536
rect 28226 22480 28276 22536
rect 28212 22476 28276 22480
rect 8156 22400 8220 22404
rect 8156 22344 8170 22400
rect 8170 22344 8220 22400
rect 8156 22340 8220 22344
rect 24348 22400 24412 22404
rect 24348 22344 24398 22400
rect 24398 22344 24412 22400
rect 24348 22340 24412 22344
rect 24900 22340 24964 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 32812 22204 32876 22268
rect 11284 22068 11348 22132
rect 13860 22068 13924 22132
rect 23060 22128 23124 22132
rect 23060 22072 23074 22128
rect 23074 22072 23124 22128
rect 23060 22068 23124 22072
rect 32444 22068 32508 22132
rect 6684 21932 6748 21996
rect 10916 21932 10980 21996
rect 12204 21932 12268 21996
rect 20300 21932 20364 21996
rect 26372 21932 26436 21996
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 15516 21524 15580 21588
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 13308 21116 13372 21180
rect 5396 20844 5460 20908
rect 15332 20844 15396 20908
rect 20484 20708 20548 20772
rect 27660 20708 27724 20772
rect 34100 20708 34164 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 8340 20632 8404 20636
rect 8340 20576 8354 20632
rect 8354 20576 8404 20632
rect 8340 20572 8404 20576
rect 16252 20632 16316 20636
rect 16252 20576 16266 20632
rect 16266 20576 16316 20632
rect 16252 20572 16316 20576
rect 5948 20436 6012 20500
rect 11652 20164 11716 20228
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 5764 19892 5828 19956
rect 26004 19816 26068 19820
rect 26004 19760 26018 19816
rect 26018 19760 26068 19816
rect 26004 19756 26068 19760
rect 14780 19620 14844 19684
rect 20852 19620 20916 19684
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 16804 19484 16868 19548
rect 31156 19484 31220 19548
rect 7788 19408 7852 19412
rect 7788 19352 7838 19408
rect 7838 19352 7852 19408
rect 7788 19348 7852 19352
rect 8708 19348 8772 19412
rect 16620 19348 16684 19412
rect 15700 19272 15764 19276
rect 15700 19216 15750 19272
rect 15750 19216 15764 19272
rect 15700 19212 15764 19216
rect 22140 19348 22204 19412
rect 22876 19408 22940 19412
rect 22876 19352 22890 19408
rect 22890 19352 22940 19408
rect 22876 19348 22940 19352
rect 25268 19348 25332 19412
rect 30420 19408 30484 19412
rect 30420 19352 30434 19408
rect 30434 19352 30484 19408
rect 30420 19348 30484 19352
rect 21220 19076 21284 19140
rect 35388 19212 35452 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 16988 18940 17052 19004
rect 18644 18940 18708 19004
rect 21036 18940 21100 19004
rect 3924 18864 3988 18868
rect 3924 18808 3938 18864
rect 3938 18808 3988 18864
rect 3924 18804 3988 18808
rect 12756 18804 12820 18868
rect 24900 18804 24964 18868
rect 26740 18864 26804 18868
rect 26740 18808 26754 18864
rect 26754 18808 26804 18864
rect 26740 18804 26804 18808
rect 27660 18668 27724 18732
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 7604 18396 7668 18460
rect 25636 18260 25700 18324
rect 15332 18124 15396 18188
rect 18276 18124 18340 18188
rect 23612 18124 23676 18188
rect 28028 18260 28092 18324
rect 26188 18184 26252 18188
rect 26188 18128 26202 18184
rect 26202 18128 26252 18184
rect 26188 18124 26252 18128
rect 32076 18124 32140 18188
rect 32812 18124 32876 18188
rect 19380 17988 19444 18052
rect 21956 18048 22020 18052
rect 21956 17992 21970 18048
rect 21970 17992 22020 18048
rect 21956 17988 22020 17992
rect 23980 18048 24044 18052
rect 23980 17992 23994 18048
rect 23994 17992 24044 18048
rect 23980 17988 24044 17992
rect 24164 17988 24228 18052
rect 24900 17988 24964 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4660 17912 4724 17916
rect 4660 17856 4710 17912
rect 4710 17856 4724 17912
rect 4660 17852 4724 17856
rect 10364 17852 10428 17916
rect 10732 17852 10796 17916
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 10548 17716 10612 17780
rect 10180 17580 10244 17644
rect 28212 17580 28276 17644
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 9812 17308 9876 17372
rect 12940 17308 13004 17372
rect 15148 17308 15212 17372
rect 35388 17308 35452 17372
rect 10364 17172 10428 17236
rect 25636 17172 25700 17236
rect 10732 17036 10796 17100
rect 20484 17036 20548 17100
rect 28580 17036 28644 17100
rect 10548 16900 10612 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 25452 16764 25516 16828
rect 4660 16628 4724 16692
rect 14964 16628 15028 16692
rect 26372 16628 26436 16692
rect 22692 16416 22756 16420
rect 22692 16360 22706 16416
rect 22706 16360 22756 16416
rect 22692 16356 22756 16360
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 17172 16280 17236 16284
rect 17172 16224 17186 16280
rect 17186 16224 17236 16280
rect 17172 16220 17236 16224
rect 16620 15948 16684 16012
rect 23796 15948 23860 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 8340 15540 8404 15604
rect 10180 15540 10244 15604
rect 31524 15600 31588 15604
rect 31524 15544 31574 15600
rect 31574 15544 31588 15600
rect 31524 15540 31588 15544
rect 25084 15404 25148 15468
rect 21588 15268 21652 15332
rect 29316 15268 29380 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 2636 15132 2700 15196
rect 10916 15132 10980 15196
rect 19564 15132 19628 15196
rect 32260 15132 32324 15196
rect 21220 14996 21284 15060
rect 19748 14860 19812 14924
rect 21036 14860 21100 14924
rect 26188 14860 26252 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 8708 14512 8772 14516
rect 8708 14456 8722 14512
rect 8722 14456 8772 14512
rect 8708 14452 8772 14456
rect 9260 14452 9324 14516
rect 9996 14512 10060 14516
rect 9996 14456 10010 14512
rect 10010 14456 10060 14512
rect 9996 14452 10060 14456
rect 11284 14512 11348 14516
rect 11284 14456 11298 14512
rect 11298 14456 11348 14512
rect 11284 14452 11348 14456
rect 27292 14452 27356 14516
rect 35388 14452 35452 14516
rect 28212 14180 28276 14244
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 14780 13908 14844 13972
rect 4660 13832 4724 13836
rect 4660 13776 4674 13832
rect 4674 13776 4724 13832
rect 4660 13772 4724 13776
rect 9076 13636 9140 13700
rect 30604 13636 30668 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 30052 13364 30116 13428
rect 5580 13228 5644 13292
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 19380 13016 19444 13020
rect 19380 12960 19394 13016
rect 19394 12960 19444 13016
rect 19380 12956 19444 12960
rect 26004 12956 26068 13020
rect 3924 12820 3988 12884
rect 17540 12880 17604 12884
rect 17540 12824 17590 12880
rect 17590 12824 17604 12880
rect 17540 12820 17604 12824
rect 7236 12744 7300 12748
rect 7236 12688 7250 12744
rect 7250 12688 7300 12744
rect 7236 12684 7300 12688
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 5764 12412 5828 12476
rect 30788 12276 30852 12340
rect 32996 12276 33060 12340
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 16620 11928 16684 11932
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 16620 11872 16670 11928
rect 16670 11872 16684 11928
rect 16620 11868 16684 11872
rect 26740 11928 26804 11932
rect 26740 11872 26754 11928
rect 26754 11872 26804 11928
rect 26740 11868 26804 11872
rect 25084 11732 25148 11796
rect 26188 11732 26252 11796
rect 30052 11792 30116 11796
rect 30052 11736 30102 11792
rect 30102 11736 30116 11792
rect 30052 11732 30116 11736
rect 26372 11596 26436 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 25636 11324 25700 11388
rect 30420 11188 30484 11252
rect 32260 10916 32324 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 23060 10644 23124 10708
rect 25636 10644 25700 10708
rect 30604 10372 30668 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 24348 10236 24412 10300
rect 29500 10236 29564 10300
rect 31156 10296 31220 10300
rect 31156 10240 31206 10296
rect 31206 10240 31220 10296
rect 31156 10236 31220 10240
rect 3924 10100 3988 10164
rect 34284 10236 34348 10300
rect 32444 10024 32508 10028
rect 32444 9968 32494 10024
rect 32494 9968 32508 10024
rect 32444 9964 32508 9968
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 34100 9692 34164 9756
rect 5580 9556 5644 9620
rect 19564 9556 19628 9620
rect 12756 9420 12820 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 17908 9148 17972 9212
rect 26188 9208 26252 9212
rect 26188 9152 26202 9208
rect 26202 9152 26252 9208
rect 26188 9148 26252 9152
rect 5764 9012 5828 9076
rect 4660 8936 4724 8940
rect 4660 8880 4710 8936
rect 4710 8880 4724 8936
rect 4660 8876 4724 8880
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 6684 8604 6748 8668
rect 32996 8664 33060 8668
rect 32996 8608 33010 8664
rect 33010 8608 33060 8664
rect 32996 8604 33060 8608
rect 5396 8468 5460 8532
rect 9628 8528 9692 8532
rect 9628 8472 9678 8528
rect 9678 8472 9692 8528
rect 9628 8468 9692 8472
rect 11100 8392 11164 8396
rect 11100 8336 11114 8392
rect 11114 8336 11164 8392
rect 11100 8332 11164 8336
rect 26372 8196 26436 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 14228 7984 14292 7988
rect 14228 7928 14242 7984
rect 14242 7928 14292 7984
rect 14228 7924 14292 7928
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 8340 7516 8404 7580
rect 28028 7924 28092 7988
rect 28580 7984 28644 7988
rect 28580 7928 28594 7984
rect 28594 7928 28644 7984
rect 28580 7924 28644 7928
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 33548 7516 33612 7580
rect 29132 7244 29196 7308
rect 23980 7108 24044 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 7236 6836 7300 6900
rect 9260 6896 9324 6900
rect 9260 6840 9274 6896
rect 9274 6840 9324 6896
rect 9260 6836 9324 6840
rect 11652 6836 11716 6900
rect 15332 6836 15396 6900
rect 21220 6836 21284 6900
rect 22876 6896 22940 6900
rect 22876 6840 22890 6896
rect 22890 6840 22940 6896
rect 22876 6836 22940 6840
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 11468 6488 11532 6492
rect 11468 6432 11518 6488
rect 11518 6432 11532 6488
rect 11468 6428 11532 6432
rect 17540 6428 17604 6492
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 32076 5884 32140 5948
rect 13492 5672 13556 5676
rect 13492 5616 13542 5672
rect 13542 5616 13556 5672
rect 13492 5612 13556 5616
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 21404 5340 21468 5404
rect 18644 5204 18708 5268
rect 19748 5068 19812 5132
rect 30420 5128 30484 5132
rect 30420 5072 30434 5128
rect 30434 5072 30484 5128
rect 30420 5068 30484 5072
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 21956 4524 22020 4588
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 18460 4312 18524 4316
rect 18460 4256 18474 4312
rect 18474 4256 18524 4312
rect 18460 4252 18524 4256
rect 16252 4116 16316 4180
rect 11100 4040 11164 4044
rect 11100 3984 11150 4040
rect 11150 3984 11164 4040
rect 11100 3980 11164 3984
rect 22692 3980 22756 4044
rect 24900 3980 24964 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 21036 3632 21100 3636
rect 21036 3576 21086 3632
rect 21086 3576 21100 3632
rect 21036 3572 21100 3576
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 20484 3224 20548 3228
rect 20484 3168 20498 3224
rect 20498 3168 20548 3224
rect 20484 3164 20548 3168
rect 14596 3028 14660 3092
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 20299 34916 20365 34917
rect 20299 34852 20300 34916
rect 20364 34852 20365 34916
rect 20299 34851 20365 34852
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4659 33012 4725 33013
rect 4659 32948 4660 33012
rect 4724 32948 4725 33012
rect 4659 32947 4725 32948
rect 4662 32333 4722 32947
rect 4868 32672 5188 33696
rect 9627 33148 9693 33149
rect 9627 33084 9628 33148
rect 9692 33084 9693 33148
rect 9627 33083 9693 33084
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4659 32332 4725 32333
rect 4659 32268 4660 32332
rect 4724 32268 4725 32332
rect 4659 32267 4725 32268
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 2635 23084 2701 23085
rect 2635 23020 2636 23084
rect 2700 23020 2701 23084
rect 2635 23019 2701 23020
rect 2638 15197 2698 23019
rect 3923 22948 3989 22949
rect 3923 22884 3924 22948
rect 3988 22884 3989 22948
rect 3923 22883 3989 22884
rect 3926 18869 3986 22883
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 3923 18868 3989 18869
rect 3923 18804 3924 18868
rect 3988 18804 3989 18868
rect 3923 18803 3989 18804
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4868 31584 5188 32608
rect 5579 31788 5645 31789
rect 5579 31724 5580 31788
rect 5644 31724 5645 31788
rect 5579 31723 5645 31724
rect 5582 31653 5642 31723
rect 5579 31652 5645 31653
rect 5579 31588 5580 31652
rect 5644 31588 5645 31652
rect 5579 31587 5645 31588
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 6315 30428 6381 30429
rect 6315 30364 6316 30428
rect 6380 30364 6381 30428
rect 6315 30363 6381 30364
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 5763 27300 5829 27301
rect 5763 27236 5764 27300
rect 5828 27236 5829 27300
rect 5763 27235 5829 27236
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 5395 20908 5461 20909
rect 5395 20844 5396 20908
rect 5460 20844 5461 20908
rect 5395 20843 5461 20844
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4659 17916 4725 17917
rect 4659 17852 4660 17916
rect 4724 17852 4725 17916
rect 4659 17851 4725 17852
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4662 16693 4722 17851
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4659 16692 4725 16693
rect 4659 16628 4660 16692
rect 4724 16628 4725 16692
rect 4659 16627 4725 16628
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 2635 15196 2701 15197
rect 2635 15132 2636 15196
rect 2700 15132 2701 15196
rect 2635 15131 2701 15132
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4659 13836 4725 13837
rect 4659 13772 4660 13836
rect 4724 13772 4725 13836
rect 4659 13771 4725 13772
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 3926 10165 3986 12819
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3923 10164 3989 10165
rect 3923 10100 3924 10164
rect 3988 10100 3989 10164
rect 3923 10099 3989 10100
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4662 8941 4722 13771
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4659 8940 4725 8941
rect 4659 8876 4660 8940
rect 4724 8876 4725 8940
rect 4659 8875 4725 8876
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 5398 8533 5458 20843
rect 5766 19957 5826 27235
rect 5947 25124 6013 25125
rect 5947 25060 5948 25124
rect 6012 25060 6013 25124
rect 5947 25059 6013 25060
rect 5950 20501 6010 25059
rect 6318 22949 6378 30363
rect 9630 30293 9690 33083
rect 10915 33012 10981 33013
rect 10915 32948 10916 33012
rect 10980 32948 10981 33012
rect 10915 32947 10981 32948
rect 9627 30292 9693 30293
rect 9627 30228 9628 30292
rect 9692 30228 9693 30292
rect 9627 30227 9693 30228
rect 9075 30156 9141 30157
rect 9075 30092 9076 30156
rect 9140 30092 9141 30156
rect 9075 30091 9141 30092
rect 7603 27300 7669 27301
rect 7603 27236 7604 27300
rect 7668 27236 7669 27300
rect 7603 27235 7669 27236
rect 6315 22948 6381 22949
rect 6315 22884 6316 22948
rect 6380 22884 6381 22948
rect 6315 22883 6381 22884
rect 6683 21996 6749 21997
rect 6683 21932 6684 21996
rect 6748 21932 6749 21996
rect 6683 21931 6749 21932
rect 5947 20500 6013 20501
rect 5947 20436 5948 20500
rect 6012 20436 6013 20500
rect 5947 20435 6013 20436
rect 5763 19956 5829 19957
rect 5763 19892 5764 19956
rect 5828 19892 5829 19956
rect 5763 19891 5829 19892
rect 5579 13292 5645 13293
rect 5579 13228 5580 13292
rect 5644 13228 5645 13292
rect 5579 13227 5645 13228
rect 5582 9621 5642 13227
rect 5763 12476 5829 12477
rect 5763 12412 5764 12476
rect 5828 12412 5829 12476
rect 5763 12411 5829 12412
rect 5579 9620 5645 9621
rect 5579 9556 5580 9620
rect 5644 9556 5645 9620
rect 5579 9555 5645 9556
rect 5766 9077 5826 12411
rect 5763 9076 5829 9077
rect 5763 9012 5764 9076
rect 5828 9012 5829 9076
rect 5763 9011 5829 9012
rect 6686 8669 6746 21931
rect 7606 18461 7666 27235
rect 8339 26348 8405 26349
rect 8339 26284 8340 26348
rect 8404 26284 8405 26348
rect 8339 26283 8405 26284
rect 7787 25668 7853 25669
rect 7787 25604 7788 25668
rect 7852 25604 7853 25668
rect 7787 25603 7853 25604
rect 7790 19413 7850 25603
rect 8155 22404 8221 22405
rect 8155 22340 8156 22404
rect 8220 22340 8221 22404
rect 8155 22339 8221 22340
rect 7787 19412 7853 19413
rect 7787 19348 7788 19412
rect 7852 19348 7853 19412
rect 7787 19347 7853 19348
rect 7603 18460 7669 18461
rect 7603 18396 7604 18460
rect 7668 18396 7669 18460
rect 7603 18395 7669 18396
rect 8158 16690 8218 22339
rect 8342 20637 8402 26283
rect 9078 22541 9138 30091
rect 9995 29476 10061 29477
rect 9995 29412 9996 29476
rect 10060 29412 10061 29476
rect 9995 29411 10061 29412
rect 9811 27572 9877 27573
rect 9811 27508 9812 27572
rect 9876 27508 9877 27572
rect 9811 27507 9877 27508
rect 9627 23492 9693 23493
rect 9627 23428 9628 23492
rect 9692 23428 9693 23492
rect 9627 23427 9693 23428
rect 9075 22540 9141 22541
rect 9075 22476 9076 22540
rect 9140 22476 9141 22540
rect 9075 22475 9141 22476
rect 8339 20636 8405 20637
rect 8339 20572 8340 20636
rect 8404 20572 8405 20636
rect 8339 20571 8405 20572
rect 8707 19412 8773 19413
rect 8707 19348 8708 19412
rect 8772 19348 8773 19412
rect 8707 19347 8773 19348
rect 8158 16630 8402 16690
rect 8342 15605 8402 16630
rect 8339 15604 8405 15605
rect 8339 15540 8340 15604
rect 8404 15540 8405 15604
rect 8339 15539 8405 15540
rect 7235 12748 7301 12749
rect 7235 12684 7236 12748
rect 7300 12684 7301 12748
rect 7235 12683 7301 12684
rect 6683 8668 6749 8669
rect 6683 8604 6684 8668
rect 6748 8604 6749 8668
rect 6683 8603 6749 8604
rect 5395 8532 5461 8533
rect 5395 8468 5396 8532
rect 5460 8468 5461 8532
rect 5395 8467 5461 8468
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 7238 6901 7298 12683
rect 8342 7581 8402 15539
rect 8710 14517 8770 19347
rect 8707 14516 8773 14517
rect 8707 14452 8708 14516
rect 8772 14452 8773 14516
rect 8707 14451 8773 14452
rect 9078 13701 9138 22475
rect 9259 14516 9325 14517
rect 9259 14452 9260 14516
rect 9324 14452 9325 14516
rect 9259 14451 9325 14452
rect 9075 13700 9141 13701
rect 9075 13636 9076 13700
rect 9140 13636 9141 13700
rect 9075 13635 9141 13636
rect 8339 7580 8405 7581
rect 8339 7516 8340 7580
rect 8404 7516 8405 7580
rect 8339 7515 8405 7516
rect 9262 6901 9322 14451
rect 9630 8533 9690 23427
rect 9814 17373 9874 27507
rect 9811 17372 9877 17373
rect 9811 17308 9812 17372
rect 9876 17308 9877 17372
rect 9811 17307 9877 17308
rect 9998 14517 10058 29411
rect 10918 28797 10978 32947
rect 13307 32060 13373 32061
rect 13307 31996 13308 32060
rect 13372 31996 13373 32060
rect 13307 31995 13373 31996
rect 13123 30292 13189 30293
rect 13123 30228 13124 30292
rect 13188 30228 13189 30292
rect 13123 30227 13189 30228
rect 12203 30156 12269 30157
rect 12203 30092 12204 30156
rect 12268 30092 12269 30156
rect 12203 30091 12269 30092
rect 11099 29204 11165 29205
rect 11099 29140 11100 29204
rect 11164 29140 11165 29204
rect 11099 29139 11165 29140
rect 10915 28796 10981 28797
rect 10915 28732 10916 28796
rect 10980 28732 10981 28796
rect 10915 28731 10981 28732
rect 11102 24309 11162 29139
rect 11099 24308 11165 24309
rect 11099 24244 11100 24308
rect 11164 24244 11165 24308
rect 11099 24243 11165 24244
rect 11467 23628 11533 23629
rect 11467 23564 11468 23628
rect 11532 23564 11533 23628
rect 11467 23563 11533 23564
rect 11283 22132 11349 22133
rect 11283 22068 11284 22132
rect 11348 22068 11349 22132
rect 11283 22067 11349 22068
rect 10915 21996 10981 21997
rect 10915 21932 10916 21996
rect 10980 21932 10981 21996
rect 10915 21931 10981 21932
rect 10363 17916 10429 17917
rect 10363 17852 10364 17916
rect 10428 17852 10429 17916
rect 10363 17851 10429 17852
rect 10731 17916 10797 17917
rect 10731 17852 10732 17916
rect 10796 17852 10797 17916
rect 10731 17851 10797 17852
rect 10179 17644 10245 17645
rect 10179 17580 10180 17644
rect 10244 17580 10245 17644
rect 10179 17579 10245 17580
rect 10182 15605 10242 17579
rect 10366 17237 10426 17851
rect 10547 17780 10613 17781
rect 10547 17716 10548 17780
rect 10612 17716 10613 17780
rect 10547 17715 10613 17716
rect 10363 17236 10429 17237
rect 10363 17172 10364 17236
rect 10428 17172 10429 17236
rect 10363 17171 10429 17172
rect 10550 16965 10610 17715
rect 10734 17101 10794 17851
rect 10731 17100 10797 17101
rect 10731 17036 10732 17100
rect 10796 17036 10797 17100
rect 10731 17035 10797 17036
rect 10547 16964 10613 16965
rect 10547 16900 10548 16964
rect 10612 16900 10613 16964
rect 10547 16899 10613 16900
rect 10179 15604 10245 15605
rect 10179 15540 10180 15604
rect 10244 15540 10245 15604
rect 10179 15539 10245 15540
rect 10918 15197 10978 21931
rect 10915 15196 10981 15197
rect 10915 15132 10916 15196
rect 10980 15132 10981 15196
rect 10915 15131 10981 15132
rect 11286 14517 11346 22067
rect 9995 14516 10061 14517
rect 9995 14452 9996 14516
rect 10060 14452 10061 14516
rect 9995 14451 10061 14452
rect 11283 14516 11349 14517
rect 11283 14452 11284 14516
rect 11348 14452 11349 14516
rect 11283 14451 11349 14452
rect 9627 8532 9693 8533
rect 9627 8468 9628 8532
rect 9692 8468 9693 8532
rect 9627 8467 9693 8468
rect 11099 8396 11165 8397
rect 11099 8332 11100 8396
rect 11164 8332 11165 8396
rect 11099 8331 11165 8332
rect 7235 6900 7301 6901
rect 7235 6836 7236 6900
rect 7300 6836 7301 6900
rect 7235 6835 7301 6836
rect 9259 6900 9325 6901
rect 9259 6836 9260 6900
rect 9324 6836 9325 6900
rect 9259 6835 9325 6836
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 11102 4045 11162 8331
rect 11470 6493 11530 23563
rect 12206 21997 12266 30091
rect 12755 27844 12821 27845
rect 12755 27780 12756 27844
rect 12820 27780 12821 27844
rect 12755 27779 12821 27780
rect 12758 24581 12818 27779
rect 12755 24580 12821 24581
rect 12755 24516 12756 24580
rect 12820 24516 12821 24580
rect 12755 24515 12821 24516
rect 12939 24444 13005 24445
rect 12939 24380 12940 24444
rect 13004 24380 13005 24444
rect 12939 24379 13005 24380
rect 12203 21996 12269 21997
rect 12203 21932 12204 21996
rect 12268 21932 12269 21996
rect 12203 21931 12269 21932
rect 11651 20228 11717 20229
rect 11651 20164 11652 20228
rect 11716 20164 11717 20228
rect 11651 20163 11717 20164
rect 11654 6901 11714 20163
rect 12755 18868 12821 18869
rect 12755 18804 12756 18868
rect 12820 18804 12821 18868
rect 12755 18803 12821 18804
rect 12758 9485 12818 18803
rect 12942 17373 13002 24379
rect 13126 24309 13186 30227
rect 13123 24308 13189 24309
rect 13123 24244 13124 24308
rect 13188 24244 13189 24308
rect 13123 24243 13189 24244
rect 13310 21181 13370 31995
rect 15515 31924 15581 31925
rect 15515 31860 15516 31924
rect 15580 31860 15581 31924
rect 15515 31859 15581 31860
rect 14963 31788 15029 31789
rect 14963 31724 14964 31788
rect 15028 31724 15029 31788
rect 14963 31723 15029 31724
rect 14043 29204 14109 29205
rect 14043 29140 14044 29204
rect 14108 29140 14109 29204
rect 14043 29139 14109 29140
rect 13859 29068 13925 29069
rect 13859 29004 13860 29068
rect 13924 29004 13925 29068
rect 13859 29003 13925 29004
rect 13491 23492 13557 23493
rect 13491 23428 13492 23492
rect 13556 23428 13557 23492
rect 13491 23427 13557 23428
rect 13307 21180 13373 21181
rect 13307 21116 13308 21180
rect 13372 21116 13373 21180
rect 13307 21115 13373 21116
rect 12939 17372 13005 17373
rect 12939 17308 12940 17372
rect 13004 17308 13005 17372
rect 12939 17307 13005 17308
rect 12755 9484 12821 9485
rect 12755 9420 12756 9484
rect 12820 9420 12821 9484
rect 12755 9419 12821 9420
rect 11651 6900 11717 6901
rect 11651 6836 11652 6900
rect 11716 6836 11717 6900
rect 11651 6835 11717 6836
rect 11467 6492 11533 6493
rect 11467 6428 11468 6492
rect 11532 6428 11533 6492
rect 11467 6427 11533 6428
rect 13494 5677 13554 23427
rect 13862 22133 13922 29003
rect 14046 24853 14106 29139
rect 14043 24852 14109 24853
rect 14043 24788 14044 24852
rect 14108 24788 14109 24852
rect 14043 24787 14109 24788
rect 14595 23764 14661 23765
rect 14595 23700 14596 23764
rect 14660 23700 14661 23764
rect 14595 23699 14661 23700
rect 14227 23628 14293 23629
rect 14227 23564 14228 23628
rect 14292 23564 14293 23628
rect 14227 23563 14293 23564
rect 13859 22132 13925 22133
rect 13859 22068 13860 22132
rect 13924 22068 13925 22132
rect 13859 22067 13925 22068
rect 14230 7989 14290 23563
rect 14227 7988 14293 7989
rect 14227 7924 14228 7988
rect 14292 7924 14293 7988
rect 14227 7923 14293 7924
rect 13491 5676 13557 5677
rect 13491 5612 13492 5676
rect 13556 5612 13557 5676
rect 13491 5611 13557 5612
rect 11099 4044 11165 4045
rect 11099 3980 11100 4044
rect 11164 3980 11165 4044
rect 11099 3979 11165 3980
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 14598 3093 14658 23699
rect 14779 19684 14845 19685
rect 14779 19620 14780 19684
rect 14844 19620 14845 19684
rect 14779 19619 14845 19620
rect 14782 13973 14842 19619
rect 14966 16693 15026 31723
rect 15331 31244 15397 31245
rect 15331 31180 15332 31244
rect 15396 31180 15397 31244
rect 15331 31179 15397 31180
rect 15147 29068 15213 29069
rect 15147 29004 15148 29068
rect 15212 29004 15213 29068
rect 15147 29003 15213 29004
rect 15150 17373 15210 29003
rect 15334 20909 15394 31179
rect 15518 21589 15578 31859
rect 19195 29068 19261 29069
rect 19195 29004 19196 29068
rect 19260 29004 19261 29068
rect 19195 29003 19261 29004
rect 15699 28524 15765 28525
rect 15699 28460 15700 28524
rect 15764 28460 15765 28524
rect 15699 28459 15765 28460
rect 15515 21588 15581 21589
rect 15515 21524 15516 21588
rect 15580 21524 15581 21588
rect 15515 21523 15581 21524
rect 15331 20908 15397 20909
rect 15331 20844 15332 20908
rect 15396 20844 15397 20908
rect 15331 20843 15397 20844
rect 15702 19277 15762 28459
rect 18459 27708 18525 27709
rect 18459 27644 18460 27708
rect 18524 27644 18525 27708
rect 18459 27643 18525 27644
rect 16619 26348 16685 26349
rect 16619 26284 16620 26348
rect 16684 26284 16685 26348
rect 16619 26283 16685 26284
rect 17171 26348 17237 26349
rect 17171 26284 17172 26348
rect 17236 26284 17237 26348
rect 17171 26283 17237 26284
rect 17907 26348 17973 26349
rect 17907 26284 17908 26348
rect 17972 26284 17973 26348
rect 17907 26283 17973 26284
rect 16251 20636 16317 20637
rect 16251 20572 16252 20636
rect 16316 20572 16317 20636
rect 16251 20571 16317 20572
rect 15699 19276 15765 19277
rect 15699 19212 15700 19276
rect 15764 19212 15765 19276
rect 15699 19211 15765 19212
rect 15331 18188 15397 18189
rect 15331 18124 15332 18188
rect 15396 18124 15397 18188
rect 15331 18123 15397 18124
rect 15147 17372 15213 17373
rect 15147 17308 15148 17372
rect 15212 17308 15213 17372
rect 15147 17307 15213 17308
rect 14963 16692 15029 16693
rect 14963 16628 14964 16692
rect 15028 16628 15029 16692
rect 14963 16627 15029 16628
rect 14779 13972 14845 13973
rect 14779 13908 14780 13972
rect 14844 13908 14845 13972
rect 14779 13907 14845 13908
rect 15334 6901 15394 18123
rect 15331 6900 15397 6901
rect 15331 6836 15332 6900
rect 15396 6836 15397 6900
rect 15331 6835 15397 6836
rect 16254 4181 16314 20571
rect 16622 19413 16682 26283
rect 16803 24444 16869 24445
rect 16803 24380 16804 24444
rect 16868 24380 16869 24444
rect 16803 24379 16869 24380
rect 16806 23085 16866 24379
rect 16987 23356 17053 23357
rect 16987 23292 16988 23356
rect 17052 23292 17053 23356
rect 16987 23291 17053 23292
rect 16803 23084 16869 23085
rect 16803 23020 16804 23084
rect 16868 23020 16869 23084
rect 16803 23019 16869 23020
rect 16806 19549 16866 23019
rect 16803 19548 16869 19549
rect 16803 19484 16804 19548
rect 16868 19484 16869 19548
rect 16803 19483 16869 19484
rect 16619 19412 16685 19413
rect 16619 19348 16620 19412
rect 16684 19348 16685 19412
rect 16619 19347 16685 19348
rect 16990 19005 17050 23291
rect 16987 19004 17053 19005
rect 16987 18940 16988 19004
rect 17052 18940 17053 19004
rect 16987 18939 17053 18940
rect 17174 16285 17234 26283
rect 17171 16284 17237 16285
rect 17171 16220 17172 16284
rect 17236 16220 17237 16284
rect 17171 16219 17237 16220
rect 16619 16012 16685 16013
rect 16619 15948 16620 16012
rect 16684 15948 16685 16012
rect 16619 15947 16685 15948
rect 16622 11933 16682 15947
rect 17539 12884 17605 12885
rect 17539 12820 17540 12884
rect 17604 12820 17605 12884
rect 17539 12819 17605 12820
rect 16619 11932 16685 11933
rect 16619 11868 16620 11932
rect 16684 11868 16685 11932
rect 16619 11867 16685 11868
rect 17542 6493 17602 12819
rect 17910 9213 17970 26283
rect 18275 24988 18341 24989
rect 18275 24924 18276 24988
rect 18340 24924 18341 24988
rect 18275 24923 18341 24924
rect 18278 18189 18338 24923
rect 18275 18188 18341 18189
rect 18275 18124 18276 18188
rect 18340 18124 18341 18188
rect 18275 18123 18341 18124
rect 17907 9212 17973 9213
rect 17907 9148 17908 9212
rect 17972 9148 17973 9212
rect 17907 9147 17973 9148
rect 17539 6492 17605 6493
rect 17539 6428 17540 6492
rect 17604 6428 17605 6492
rect 17539 6427 17605 6428
rect 18462 4317 18522 27643
rect 19198 22813 19258 29003
rect 19195 22812 19261 22813
rect 19195 22748 19196 22812
rect 19260 22748 19261 22812
rect 19195 22747 19261 22748
rect 20302 21997 20362 34851
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 26371 32060 26437 32061
rect 26371 31996 26372 32060
rect 26436 31996 26437 32060
rect 26371 31995 26437 31996
rect 23795 30156 23861 30157
rect 23795 30092 23796 30156
rect 23860 30092 23861 30156
rect 23795 30091 23861 30092
rect 22875 27844 22941 27845
rect 22875 27780 22876 27844
rect 22940 27780 22941 27844
rect 22875 27779 22941 27780
rect 21403 26620 21469 26621
rect 21403 26556 21404 26620
rect 21468 26556 21469 26620
rect 21403 26555 21469 26556
rect 21035 26348 21101 26349
rect 21035 26284 21036 26348
rect 21100 26284 21101 26348
rect 21035 26283 21101 26284
rect 20851 24172 20917 24173
rect 20851 24108 20852 24172
rect 20916 24108 20917 24172
rect 20851 24107 20917 24108
rect 20299 21996 20365 21997
rect 20299 21932 20300 21996
rect 20364 21932 20365 21996
rect 20299 21931 20365 21932
rect 20483 20772 20549 20773
rect 20483 20708 20484 20772
rect 20548 20708 20549 20772
rect 20483 20707 20549 20708
rect 18643 19004 18709 19005
rect 18643 18940 18644 19004
rect 18708 18940 18709 19004
rect 18643 18939 18709 18940
rect 18646 5269 18706 18939
rect 19379 18052 19445 18053
rect 19379 17988 19380 18052
rect 19444 17988 19445 18052
rect 19379 17987 19445 17988
rect 19382 13021 19442 17987
rect 20486 17101 20546 20707
rect 20854 19685 20914 24107
rect 20851 19684 20917 19685
rect 20851 19620 20852 19684
rect 20916 19620 20917 19684
rect 20851 19619 20917 19620
rect 21038 19005 21098 26283
rect 21219 23764 21285 23765
rect 21219 23700 21220 23764
rect 21284 23700 21285 23764
rect 21219 23699 21285 23700
rect 21222 19141 21282 23699
rect 21219 19140 21285 19141
rect 21219 19076 21220 19140
rect 21284 19076 21285 19140
rect 21219 19075 21285 19076
rect 21035 19004 21101 19005
rect 21035 18940 21036 19004
rect 21100 18940 21101 19004
rect 21035 18939 21101 18940
rect 20483 17100 20549 17101
rect 20483 17036 20484 17100
rect 20548 17036 20549 17100
rect 20483 17035 20549 17036
rect 19563 15196 19629 15197
rect 19563 15132 19564 15196
rect 19628 15132 19629 15196
rect 19563 15131 19629 15132
rect 19379 13020 19445 13021
rect 19379 12956 19380 13020
rect 19444 12956 19445 13020
rect 19379 12955 19445 12956
rect 19566 9621 19626 15131
rect 19747 14924 19813 14925
rect 19747 14860 19748 14924
rect 19812 14860 19813 14924
rect 19747 14859 19813 14860
rect 19563 9620 19629 9621
rect 19563 9556 19564 9620
rect 19628 9556 19629 9620
rect 19563 9555 19629 9556
rect 18643 5268 18709 5269
rect 18643 5204 18644 5268
rect 18708 5204 18709 5268
rect 18643 5203 18709 5204
rect 19750 5133 19810 14859
rect 19747 5132 19813 5133
rect 19747 5068 19748 5132
rect 19812 5068 19813 5132
rect 19747 5067 19813 5068
rect 18459 4316 18525 4317
rect 18459 4252 18460 4316
rect 18524 4252 18525 4316
rect 18459 4251 18525 4252
rect 16251 4180 16317 4181
rect 16251 4116 16252 4180
rect 16316 4116 16317 4180
rect 16251 4115 16317 4116
rect 20486 3229 20546 17035
rect 21219 15060 21285 15061
rect 21219 14996 21220 15060
rect 21284 14996 21285 15060
rect 21219 14995 21285 14996
rect 21035 14924 21101 14925
rect 21035 14860 21036 14924
rect 21100 14860 21101 14924
rect 21035 14859 21101 14860
rect 21038 3637 21098 14859
rect 21222 6901 21282 14995
rect 21219 6900 21285 6901
rect 21219 6836 21220 6900
rect 21284 6836 21285 6900
rect 21219 6835 21285 6836
rect 21406 5405 21466 26555
rect 22139 26484 22205 26485
rect 22139 26420 22140 26484
rect 22204 26420 22205 26484
rect 22139 26419 22205 26420
rect 21587 22540 21653 22541
rect 21587 22476 21588 22540
rect 21652 22476 21653 22540
rect 21587 22475 21653 22476
rect 21590 15333 21650 22475
rect 22142 19413 22202 26419
rect 22691 26348 22757 26349
rect 22691 26284 22692 26348
rect 22756 26284 22757 26348
rect 22691 26283 22757 26284
rect 22139 19412 22205 19413
rect 22139 19348 22140 19412
rect 22204 19348 22205 19412
rect 22139 19347 22205 19348
rect 21955 18052 22021 18053
rect 21955 17988 21956 18052
rect 22020 17988 22021 18052
rect 21955 17987 22021 17988
rect 21587 15332 21653 15333
rect 21587 15268 21588 15332
rect 21652 15268 21653 15332
rect 21587 15267 21653 15268
rect 21403 5404 21469 5405
rect 21403 5340 21404 5404
rect 21468 5340 21469 5404
rect 21403 5339 21469 5340
rect 21958 4589 22018 17987
rect 22694 16421 22754 26283
rect 22878 19413 22938 27779
rect 23611 23900 23677 23901
rect 23611 23836 23612 23900
rect 23676 23836 23677 23900
rect 23611 23835 23677 23836
rect 23059 22132 23125 22133
rect 23059 22068 23060 22132
rect 23124 22068 23125 22132
rect 23059 22067 23125 22068
rect 22875 19412 22941 19413
rect 22875 19348 22876 19412
rect 22940 19348 22941 19412
rect 22875 19347 22941 19348
rect 22691 16420 22757 16421
rect 22691 16356 22692 16420
rect 22756 16356 22757 16420
rect 22691 16355 22757 16356
rect 21955 4588 22021 4589
rect 21955 4524 21956 4588
rect 22020 4524 22021 4588
rect 21955 4523 22021 4524
rect 22694 4045 22754 16355
rect 22878 6901 22938 19347
rect 23062 10709 23122 22067
rect 23614 18189 23674 23835
rect 23611 18188 23677 18189
rect 23611 18124 23612 18188
rect 23676 18124 23677 18188
rect 23611 18123 23677 18124
rect 23798 16013 23858 30091
rect 26187 29748 26253 29749
rect 26187 29684 26188 29748
rect 26252 29684 26253 29748
rect 26187 29683 26253 29684
rect 24163 29612 24229 29613
rect 24163 29548 24164 29612
rect 24228 29548 24229 29612
rect 24163 29547 24229 29548
rect 24166 25805 24226 29547
rect 25267 29476 25333 29477
rect 25267 29412 25268 29476
rect 25332 29412 25333 29476
rect 25267 29411 25333 29412
rect 24163 25804 24229 25805
rect 24163 25740 24164 25804
rect 24228 25740 24229 25804
rect 24163 25739 24229 25740
rect 24166 18053 24226 25739
rect 24347 22404 24413 22405
rect 24347 22340 24348 22404
rect 24412 22340 24413 22404
rect 24347 22339 24413 22340
rect 24899 22404 24965 22405
rect 24899 22340 24900 22404
rect 24964 22340 24965 22404
rect 24899 22339 24965 22340
rect 23979 18052 24045 18053
rect 23979 17988 23980 18052
rect 24044 17988 24045 18052
rect 23979 17987 24045 17988
rect 24163 18052 24229 18053
rect 24163 17988 24164 18052
rect 24228 17988 24229 18052
rect 24163 17987 24229 17988
rect 23795 16012 23861 16013
rect 23795 15948 23796 16012
rect 23860 15948 23861 16012
rect 23795 15947 23861 15948
rect 23059 10708 23125 10709
rect 23059 10644 23060 10708
rect 23124 10644 23125 10708
rect 23059 10643 23125 10644
rect 23982 7173 24042 17987
rect 24350 10301 24410 22339
rect 24902 18869 24962 22339
rect 25270 19413 25330 29411
rect 26003 28116 26069 28117
rect 26003 28052 26004 28116
rect 26068 28052 26069 28116
rect 26003 28051 26069 28052
rect 25451 22676 25517 22677
rect 25451 22612 25452 22676
rect 25516 22612 25517 22676
rect 25451 22611 25517 22612
rect 25267 19412 25333 19413
rect 25267 19348 25268 19412
rect 25332 19348 25333 19412
rect 25267 19347 25333 19348
rect 24899 18868 24965 18869
rect 24899 18804 24900 18868
rect 24964 18804 24965 18868
rect 24899 18803 24965 18804
rect 24899 18052 24965 18053
rect 24899 17988 24900 18052
rect 24964 17988 24965 18052
rect 24899 17987 24965 17988
rect 24347 10300 24413 10301
rect 24347 10236 24348 10300
rect 24412 10236 24413 10300
rect 24347 10235 24413 10236
rect 23979 7172 24045 7173
rect 23979 7108 23980 7172
rect 24044 7108 24045 7172
rect 23979 7107 24045 7108
rect 22875 6900 22941 6901
rect 22875 6836 22876 6900
rect 22940 6836 22941 6900
rect 22875 6835 22941 6836
rect 24902 4045 24962 17987
rect 25454 16829 25514 22611
rect 26006 19821 26066 28051
rect 26190 27573 26250 29683
rect 26374 28253 26434 31995
rect 27475 31788 27541 31789
rect 27475 31724 27476 31788
rect 27540 31724 27541 31788
rect 27475 31723 27541 31724
rect 27659 31788 27725 31789
rect 27659 31724 27660 31788
rect 27724 31724 27725 31788
rect 27659 31723 27725 31724
rect 27291 31516 27357 31517
rect 27291 31452 27292 31516
rect 27356 31452 27357 31516
rect 27291 31451 27357 31452
rect 27294 29477 27354 31451
rect 27478 30157 27538 31723
rect 27475 30156 27541 30157
rect 27475 30092 27476 30156
rect 27540 30092 27541 30156
rect 27475 30091 27541 30092
rect 27291 29476 27357 29477
rect 27291 29412 27292 29476
rect 27356 29412 27357 29476
rect 27291 29411 27357 29412
rect 26371 28252 26437 28253
rect 26371 28188 26372 28252
rect 26436 28188 26437 28252
rect 26371 28187 26437 28188
rect 27291 27708 27357 27709
rect 27291 27644 27292 27708
rect 27356 27644 27357 27708
rect 27291 27643 27357 27644
rect 26187 27572 26253 27573
rect 26187 27508 26188 27572
rect 26252 27508 26253 27572
rect 26187 27507 26253 27508
rect 26371 21996 26437 21997
rect 26371 21932 26372 21996
rect 26436 21932 26437 21996
rect 26371 21931 26437 21932
rect 26003 19820 26069 19821
rect 26003 19756 26004 19820
rect 26068 19756 26069 19820
rect 26003 19755 26069 19756
rect 25635 18324 25701 18325
rect 25635 18260 25636 18324
rect 25700 18260 25701 18324
rect 25635 18259 25701 18260
rect 25638 17237 25698 18259
rect 25635 17236 25701 17237
rect 25635 17172 25636 17236
rect 25700 17172 25701 17236
rect 25635 17171 25701 17172
rect 25451 16828 25517 16829
rect 25451 16764 25452 16828
rect 25516 16764 25517 16828
rect 25451 16763 25517 16764
rect 25083 15468 25149 15469
rect 25083 15404 25084 15468
rect 25148 15404 25149 15468
rect 25083 15403 25149 15404
rect 25086 11797 25146 15403
rect 25083 11796 25149 11797
rect 25083 11732 25084 11796
rect 25148 11732 25149 11796
rect 25083 11731 25149 11732
rect 25638 11389 25698 17171
rect 26006 13021 26066 19755
rect 26187 18188 26253 18189
rect 26187 18124 26188 18188
rect 26252 18124 26253 18188
rect 26187 18123 26253 18124
rect 26190 14925 26250 18123
rect 26374 16693 26434 21931
rect 26739 18868 26805 18869
rect 26739 18804 26740 18868
rect 26804 18804 26805 18868
rect 26739 18803 26805 18804
rect 26371 16692 26437 16693
rect 26371 16628 26372 16692
rect 26436 16628 26437 16692
rect 26371 16627 26437 16628
rect 26187 14924 26253 14925
rect 26187 14860 26188 14924
rect 26252 14860 26253 14924
rect 26187 14859 26253 14860
rect 26003 13020 26069 13021
rect 26003 12956 26004 13020
rect 26068 12956 26069 13020
rect 26003 12955 26069 12956
rect 26742 11933 26802 18803
rect 27294 14517 27354 27643
rect 27478 24173 27538 30091
rect 27662 28933 27722 31723
rect 28211 31652 28277 31653
rect 28211 31588 28212 31652
rect 28276 31588 28277 31652
rect 28211 31587 28277 31588
rect 28214 29749 28274 31587
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 28211 29748 28277 29749
rect 28211 29684 28212 29748
rect 28276 29684 28277 29748
rect 28211 29683 28277 29684
rect 30971 29612 31037 29613
rect 30971 29548 30972 29612
rect 31036 29548 31037 29612
rect 30971 29547 31037 29548
rect 30051 29068 30117 29069
rect 30051 29004 30052 29068
rect 30116 29004 30117 29068
rect 30051 29003 30117 29004
rect 27659 28932 27725 28933
rect 27659 28868 27660 28932
rect 27724 28868 27725 28932
rect 27659 28867 27725 28868
rect 27659 28796 27725 28797
rect 27659 28732 27660 28796
rect 27724 28732 27725 28796
rect 27659 28731 27725 28732
rect 27662 27981 27722 28731
rect 29131 28660 29197 28661
rect 29131 28596 29132 28660
rect 29196 28596 29197 28660
rect 29131 28595 29197 28596
rect 27659 27980 27725 27981
rect 27659 27916 27660 27980
rect 27724 27916 27725 27980
rect 27659 27915 27725 27916
rect 27475 24172 27541 24173
rect 27475 24108 27476 24172
rect 27540 24108 27541 24172
rect 27475 24107 27541 24108
rect 28211 22540 28277 22541
rect 28211 22476 28212 22540
rect 28276 22476 28277 22540
rect 28211 22475 28277 22476
rect 27659 20772 27725 20773
rect 27659 20708 27660 20772
rect 27724 20708 27725 20772
rect 27659 20707 27725 20708
rect 27662 18733 27722 20707
rect 27659 18732 27725 18733
rect 27659 18668 27660 18732
rect 27724 18668 27725 18732
rect 27659 18667 27725 18668
rect 28027 18324 28093 18325
rect 28027 18260 28028 18324
rect 28092 18260 28093 18324
rect 28027 18259 28093 18260
rect 27291 14516 27357 14517
rect 27291 14452 27292 14516
rect 27356 14452 27357 14516
rect 27291 14451 27357 14452
rect 26739 11932 26805 11933
rect 26739 11868 26740 11932
rect 26804 11868 26805 11932
rect 26739 11867 26805 11868
rect 26187 11796 26253 11797
rect 26187 11732 26188 11796
rect 26252 11732 26253 11796
rect 26187 11731 26253 11732
rect 25635 11388 25701 11389
rect 25635 11324 25636 11388
rect 25700 11324 25701 11388
rect 25635 11323 25701 11324
rect 25638 10709 25698 11323
rect 25635 10708 25701 10709
rect 25635 10644 25636 10708
rect 25700 10644 25701 10708
rect 25635 10643 25701 10644
rect 26190 9213 26250 11731
rect 26371 11660 26437 11661
rect 26371 11596 26372 11660
rect 26436 11596 26437 11660
rect 26371 11595 26437 11596
rect 26187 9212 26253 9213
rect 26187 9148 26188 9212
rect 26252 9148 26253 9212
rect 26187 9147 26253 9148
rect 26374 8261 26434 11595
rect 26371 8260 26437 8261
rect 26371 8196 26372 8260
rect 26436 8196 26437 8260
rect 26371 8195 26437 8196
rect 28030 7989 28090 18259
rect 28214 17645 28274 22475
rect 28211 17644 28277 17645
rect 28211 17580 28212 17644
rect 28276 17580 28277 17644
rect 28211 17579 28277 17580
rect 28214 14245 28274 17579
rect 28579 17100 28645 17101
rect 28579 17036 28580 17100
rect 28644 17036 28645 17100
rect 28579 17035 28645 17036
rect 28211 14244 28277 14245
rect 28211 14180 28212 14244
rect 28276 14180 28277 14244
rect 28211 14179 28277 14180
rect 28582 7989 28642 17035
rect 28027 7988 28093 7989
rect 28027 7924 28028 7988
rect 28092 7924 28093 7988
rect 28027 7923 28093 7924
rect 28579 7988 28645 7989
rect 28579 7924 28580 7988
rect 28644 7924 28645 7988
rect 28579 7923 28645 7924
rect 29134 7309 29194 28595
rect 29315 25668 29381 25669
rect 29315 25604 29316 25668
rect 29380 25604 29381 25668
rect 29315 25603 29381 25604
rect 29318 15333 29378 25603
rect 29499 22812 29565 22813
rect 29499 22748 29500 22812
rect 29564 22748 29565 22812
rect 29499 22747 29565 22748
rect 29315 15332 29381 15333
rect 29315 15268 29316 15332
rect 29380 15268 29381 15332
rect 29315 15267 29381 15268
rect 29502 10301 29562 22747
rect 30054 13429 30114 29003
rect 30419 27844 30485 27845
rect 30419 27780 30420 27844
rect 30484 27780 30485 27844
rect 30419 27779 30485 27780
rect 30422 19413 30482 27779
rect 30974 27573 31034 29547
rect 33547 29068 33613 29069
rect 33547 29004 33548 29068
rect 33612 29004 33613 29068
rect 33547 29003 33613 29004
rect 34283 29068 34349 29069
rect 34283 29004 34284 29068
rect 34348 29004 34349 29068
rect 34283 29003 34349 29004
rect 30971 27572 31037 27573
rect 30971 27508 30972 27572
rect 31036 27508 31037 27572
rect 30971 27507 31037 27508
rect 31523 26892 31589 26893
rect 31523 26828 31524 26892
rect 31588 26828 31589 26892
rect 31523 26827 31589 26828
rect 30787 23764 30853 23765
rect 30787 23700 30788 23764
rect 30852 23700 30853 23764
rect 30787 23699 30853 23700
rect 30419 19412 30485 19413
rect 30419 19348 30420 19412
rect 30484 19348 30485 19412
rect 30419 19347 30485 19348
rect 30603 13700 30669 13701
rect 30603 13636 30604 13700
rect 30668 13636 30669 13700
rect 30603 13635 30669 13636
rect 30051 13428 30117 13429
rect 30051 13364 30052 13428
rect 30116 13364 30117 13428
rect 30051 13363 30117 13364
rect 30054 11797 30114 13363
rect 30051 11796 30117 11797
rect 30051 11732 30052 11796
rect 30116 11732 30117 11796
rect 30051 11731 30117 11732
rect 30419 11252 30485 11253
rect 30419 11188 30420 11252
rect 30484 11188 30485 11252
rect 30419 11187 30485 11188
rect 29499 10300 29565 10301
rect 29499 10236 29500 10300
rect 29564 10236 29565 10300
rect 29499 10235 29565 10236
rect 29131 7308 29197 7309
rect 29131 7244 29132 7308
rect 29196 7244 29197 7308
rect 29131 7243 29197 7244
rect 30422 5133 30482 11187
rect 30606 10437 30666 13635
rect 30790 12341 30850 23699
rect 31155 23492 31221 23493
rect 31155 23428 31156 23492
rect 31220 23428 31221 23492
rect 31155 23427 31221 23428
rect 31158 19549 31218 23427
rect 31155 19548 31221 19549
rect 31155 19484 31156 19548
rect 31220 19484 31221 19548
rect 31155 19483 31221 19484
rect 30787 12340 30853 12341
rect 30787 12276 30788 12340
rect 30852 12276 30853 12340
rect 30787 12275 30853 12276
rect 30603 10436 30669 10437
rect 30603 10372 30604 10436
rect 30668 10372 30669 10436
rect 30603 10371 30669 10372
rect 31158 10301 31218 19483
rect 31526 15605 31586 26827
rect 32259 25940 32325 25941
rect 32259 25876 32260 25940
rect 32324 25876 32325 25940
rect 32259 25875 32325 25876
rect 32075 18188 32141 18189
rect 32075 18124 32076 18188
rect 32140 18124 32141 18188
rect 32075 18123 32141 18124
rect 31523 15604 31589 15605
rect 31523 15540 31524 15604
rect 31588 15540 31589 15604
rect 31523 15539 31589 15540
rect 31155 10300 31221 10301
rect 31155 10236 31156 10300
rect 31220 10236 31221 10300
rect 31155 10235 31221 10236
rect 32078 5949 32138 18123
rect 32262 15197 32322 25875
rect 32811 22268 32877 22269
rect 32811 22204 32812 22268
rect 32876 22204 32877 22268
rect 32811 22203 32877 22204
rect 32443 22132 32509 22133
rect 32443 22068 32444 22132
rect 32508 22068 32509 22132
rect 32443 22067 32509 22068
rect 32259 15196 32325 15197
rect 32259 15132 32260 15196
rect 32324 15132 32325 15196
rect 32259 15131 32325 15132
rect 32262 10981 32322 15131
rect 32259 10980 32325 10981
rect 32259 10916 32260 10980
rect 32324 10916 32325 10980
rect 32259 10915 32325 10916
rect 32446 10029 32506 22067
rect 32814 18189 32874 22203
rect 32811 18188 32877 18189
rect 32811 18124 32812 18188
rect 32876 18124 32877 18188
rect 32811 18123 32877 18124
rect 32995 12340 33061 12341
rect 32995 12276 32996 12340
rect 33060 12276 33061 12340
rect 32995 12275 33061 12276
rect 32443 10028 32509 10029
rect 32443 9964 32444 10028
rect 32508 9964 32509 10028
rect 32443 9963 32509 9964
rect 32998 8669 33058 12275
rect 32995 8668 33061 8669
rect 32995 8604 32996 8668
rect 33060 8604 33061 8668
rect 32995 8603 33061 8604
rect 33550 7581 33610 29003
rect 34099 20772 34165 20773
rect 34099 20708 34100 20772
rect 34164 20708 34165 20772
rect 34099 20707 34165 20708
rect 34102 9757 34162 20707
rect 34286 10301 34346 29003
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35387 19276 35453 19277
rect 35387 19212 35388 19276
rect 35452 19212 35453 19276
rect 35387 19211 35453 19212
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 35390 17373 35450 19211
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35387 17372 35453 17373
rect 35387 17308 35388 17372
rect 35452 17308 35453 17372
rect 35387 17307 35453 17308
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 35390 14517 35450 17307
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35387 14516 35453 14517
rect 35387 14452 35388 14516
rect 35452 14452 35453 14516
rect 35387 14451 35453 14452
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34283 10300 34349 10301
rect 34283 10236 34284 10300
rect 34348 10236 34349 10300
rect 34283 10235 34349 10236
rect 34099 9756 34165 9757
rect 34099 9692 34100 9756
rect 34164 9692 34165 9756
rect 34099 9691 34165 9692
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 33547 7580 33613 7581
rect 33547 7516 33548 7580
rect 33612 7516 33613 7580
rect 33547 7515 33613 7516
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 32075 5948 32141 5949
rect 32075 5884 32076 5948
rect 32140 5884 32141 5948
rect 32075 5883 32141 5884
rect 30419 5132 30485 5133
rect 30419 5068 30420 5132
rect 30484 5068 30485 5132
rect 30419 5067 30485 5068
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 22691 4044 22757 4045
rect 22691 3980 22692 4044
rect 22756 3980 22757 4044
rect 22691 3979 22757 3980
rect 24899 4044 24965 4045
rect 24899 3980 24900 4044
rect 24964 3980 24965 4044
rect 24899 3979 24965 3980
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 21035 3636 21101 3637
rect 21035 3572 21036 3636
rect 21100 3572 21101 3636
rect 21035 3571 21101 3572
rect 20483 3228 20549 3229
rect 20483 3164 20484 3228
rect 20548 3164 20549 3228
rect 20483 3163 20549 3164
rect 14595 3092 14661 3093
rect 14595 3028 14596 3092
rect 14660 3028 14661 3092
rect 14595 3027 14661 3028
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
use sky130_fd_sc_hd__inv_2  _1336_
timestamp 18001
transform -1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1337_
timestamp 18001
transform -1 0 28980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1338_
timestamp 18001
transform -1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 18001
transform -1 0 19504 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1340_
timestamp 18001
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1341_
timestamp 18001
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1342_
timestamp 18001
transform -1 0 16192 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1343_
timestamp 18001
transform 1 0 13616 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1344_
timestamp 18001
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1345_
timestamp 18001
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1346_
timestamp 18001
transform -1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1347_
timestamp 18001
transform -1 0 27416 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _1348_
timestamp 18001
transform -1 0 26864 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1349_
timestamp 18001
transform 1 0 24748 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1350_
timestamp 18001
transform -1 0 23276 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1351_
timestamp 18001
transform 1 0 21252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1352_
timestamp 18001
transform -1 0 31280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _1353_
timestamp 18001
transform -1 0 34224 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__and2b_2  _1354_
timestamp 18001
transform -1 0 25760 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _1355_
timestamp 18001
transform 1 0 29256 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_2  _1356_
timestamp 18001
transform -1 0 31648 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1357_
timestamp 18001
transform -1 0 28244 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1358_
timestamp 18001
transform -1 0 31924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_1  _1359_
timestamp 18001
transform 1 0 24472 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _1360_
timestamp 18001
transform 1 0 27416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1361_
timestamp 18001
transform -1 0 26864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1362_
timestamp 18001
transform -1 0 23736 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _1363_
timestamp 18001
transform -1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_2  _1364_
timestamp 18001
transform 1 0 33764 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1365_
timestamp 18001
transform -1 0 25392 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1366_
timestamp 18001
transform 1 0 32844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1367_
timestamp 18001
transform -1 0 30360 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1368_
timestamp 18001
transform -1 0 28060 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1369_
timestamp 18001
transform -1 0 24196 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1370_
timestamp 18001
transform 1 0 33764 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _1371_
timestamp 18001
transform 1 0 31832 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__and4b_4  _1372_
timestamp 18001
transform 1 0 26312 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _1373_
timestamp 18001
transform -1 0 25392 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1374_
timestamp 18001
transform -1 0 23460 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1375_
timestamp 18001
transform -1 0 19596 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1376_
timestamp 18001
transform 1 0 15548 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1377_
timestamp 18001
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 18001
transform 1 0 18216 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _1379_
timestamp 18001
transform -1 0 20884 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_2  _1380_
timestamp 18001
transform 1 0 29532 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_4  _1381_
timestamp 18001
transform -1 0 33396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _1382_
timestamp 18001
transform 1 0 32292 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1383_
timestamp 18001
transform -1 0 31924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1384_
timestamp 18001
transform -1 0 31188 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_2  _1385_
timestamp 18001
transform -1 0 26036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_4  _1386_
timestamp 18001
transform 1 0 34684 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1387_
timestamp 18001
transform -1 0 33488 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1388_
timestamp 18001
transform -1 0 33212 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1389_
timestamp 18001
transform 1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1390_
timestamp 18001
transform -1 0 24932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _1391_
timestamp 18001
transform -1 0 30544 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _1392_
timestamp 18001
transform 1 0 29256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_4  _1393_
timestamp 18001
transform 1 0 32108 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__or4bb_4  _1394_
timestamp 18001
transform 1 0 26220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1395_
timestamp 18001
transform -1 0 27784 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1396_
timestamp 18001
transform -1 0 23736 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1397_
timestamp 18001
transform -1 0 23184 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1398_
timestamp 18001
transform -1 0 31832 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1399_
timestamp 18001
transform -1 0 26128 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_2  _1400_
timestamp 18001
transform -1 0 33028 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _1401_
timestamp 18001
transform -1 0 25852 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1402_
timestamp 18001
transform 1 0 24932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_2  _1403_
timestamp 18001
transform -1 0 31280 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_4  _1404_
timestamp 18001
transform -1 0 31556 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1405_
timestamp 18001
transform -1 0 31280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1406_
timestamp 18001
transform -1 0 25024 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _1407_
timestamp 18001
transform 1 0 22724 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _1408_
timestamp 18001
transform 1 0 25116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _1409_
timestamp 18001
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1410_
timestamp 18001
transform -1 0 22632 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1411_
timestamp 18001
transform 1 0 21712 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1412_
timestamp 18001
transform -1 0 19044 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1413_
timestamp 18001
transform 1 0 17112 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1414_
timestamp 18001
transform 1 0 21528 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1415_
timestamp 18001
transform -1 0 14996 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_2  _1416_
timestamp 18001
transform 1 0 32200 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _1417_
timestamp 18001
transform -1 0 34224 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1418_
timestamp 18001
transform 1 0 28704 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _1419_
timestamp 18001
transform 1 0 29624 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1420_
timestamp 18001
transform -1 0 31832 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1421_
timestamp 18001
transform -1 0 28704 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1422_
timestamp 18001
transform -1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1423_
timestamp 18001
transform -1 0 29072 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1424_
timestamp 18001
transform 1 0 26036 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1425_
timestamp 18001
transform -1 0 27416 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1426_
timestamp 18001
transform 1 0 26864 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1427_
timestamp 18001
transform 1 0 25300 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1428_
timestamp 18001
transform -1 0 29072 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1429_
timestamp 18001
transform -1 0 27784 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1430_
timestamp 18001
transform -1 0 27876 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_4  _1431_
timestamp 18001
transform 1 0 27232 0 -1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_2  _1432_
timestamp 18001
transform -1 0 27232 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1433_
timestamp 18001
transform -1 0 21620 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1434_
timestamp 18001
transform 1 0 13432 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1435_
timestamp 18001
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1436_
timestamp 18001
transform -1 0 20700 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1437_
timestamp 18001
transform -1 0 24932 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1438_
timestamp 18001
transform 1 0 31556 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 18001
transform 1 0 22264 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1440_
timestamp 18001
transform -1 0 22080 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1441_
timestamp 18001
transform -1 0 30728 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1442_
timestamp 18001
transform -1 0 28888 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1443_
timestamp 18001
transform 1 0 24932 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1444_
timestamp 18001
transform 1 0 20976 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1445_
timestamp 18001
transform 1 0 19688 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1446_
timestamp 18001
transform -1 0 23000 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1447_
timestamp 18001
transform 1 0 20608 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1448_
timestamp 18001
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1449_
timestamp 18001
transform 1 0 32384 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1450_
timestamp 18001
transform -1 0 32568 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1451_
timestamp 18001
transform 1 0 22816 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1452_
timestamp 18001
transform 1 0 21896 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1453_
timestamp 18001
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_2  _1454_
timestamp 18001
transform 1 0 27140 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1455_
timestamp 18001
transform -1 0 28520 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 18001
transform -1 0 21252 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1457_
timestamp 18001
transform -1 0 24748 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1458_
timestamp 18001
transform -1 0 22264 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1459_
timestamp 18001
transform -1 0 21620 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 18001
transform 1 0 20884 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1461_
timestamp 18001
transform -1 0 21804 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1462_
timestamp 18001
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1463_
timestamp 18001
transform 1 0 22172 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1464_
timestamp 18001
transform -1 0 28888 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _1465_
timestamp 18001
transform 1 0 29072 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1466_
timestamp 18001
transform 1 0 26036 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1467_
timestamp 18001
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1468_
timestamp 18001
transform -1 0 31832 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1469_
timestamp 18001
transform 1 0 23644 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1470_
timestamp 18001
transform 1 0 29624 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1471_
timestamp 18001
transform 1 0 23920 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1472_
timestamp 18001
transform 1 0 24656 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1473_
timestamp 18001
transform 1 0 18124 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_2  _1474_
timestamp 18001
transform 1 0 24932 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _1475_
timestamp 18001
transform -1 0 29716 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1476_
timestamp 18001
transform 1 0 26496 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1477_
timestamp 18001
transform 1 0 27692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1478_
timestamp 18001
transform -1 0 28428 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1479_
timestamp 18001
transform -1 0 26036 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1480_
timestamp 18001
transform 1 0 25668 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1481_
timestamp 18001
transform -1 0 27692 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1482_
timestamp 18001
transform -1 0 25852 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1483_
timestamp 18001
transform 1 0 25208 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1484_
timestamp 18001
transform 1 0 25024 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1485_
timestamp 18001
transform 1 0 25116 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1486_
timestamp 18001
transform -1 0 24472 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1487_
timestamp 18001
transform -1 0 21712 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1488_
timestamp 18001
transform 1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1489_
timestamp 18001
transform -1 0 27600 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1490_
timestamp 18001
transform 1 0 26680 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1491_
timestamp 18001
transform -1 0 26128 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1492_
timestamp 18001
transform -1 0 29440 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1493_
timestamp 18001
transform -1 0 30452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1494_
timestamp 18001
transform 1 0 28428 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1495_
timestamp 18001
transform -1 0 28704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1496_
timestamp 18001
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1497_
timestamp 18001
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1498_
timestamp 18001
transform 1 0 25392 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1499_
timestamp 18001
transform 1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1500_
timestamp 18001
transform -1 0 26312 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1501_
timestamp 18001
transform -1 0 22356 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1502_
timestamp 18001
transform -1 0 23460 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1503_
timestamp 18001
transform 1 0 23552 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1504_
timestamp 18001
transform 1 0 24196 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1505_
timestamp 18001
transform 1 0 23368 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1506_
timestamp 18001
transform 1 0 23828 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 18001
transform 1 0 21160 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 18001
transform -1 0 17296 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1509_
timestamp 18001
transform -1 0 17388 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_2  _1510_
timestamp 18001
transform 1 0 22540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1511_
timestamp 18001
transform -1 0 23736 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a32oi_4  _1512_
timestamp 18001
transform 1 0 22080 0 1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__a32o_1  _1513_
timestamp 18001
transform 1 0 22356 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _1514_
timestamp 18001
transform -1 0 22080 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1515_
timestamp 18001
transform -1 0 21804 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1516_
timestamp 18001
transform -1 0 23092 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_4  _1517_
timestamp 18001
transform -1 0 23368 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _1518_
timestamp 18001
transform -1 0 23552 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_2  _1519_
timestamp 18001
transform 1 0 21896 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a211oi_4  _1520_
timestamp 18001
transform 1 0 22816 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1521_
timestamp 18001
transform 1 0 20608 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1522_
timestamp 18001
transform 1 0 21896 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1523_
timestamp 18001
transform -1 0 22632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1524_
timestamp 18001
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 18001
transform -1 0 26036 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _1526_
timestamp 18001
transform 1 0 25852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1527_
timestamp 18001
transform -1 0 24012 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1528_
timestamp 18001
transform 1 0 24104 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1529_
timestamp 18001
transform 1 0 21988 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1530_
timestamp 18001
transform 1 0 21068 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1531_
timestamp 18001
transform 1 0 18124 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1532_
timestamp 18001
transform -1 0 19596 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1533_
timestamp 18001
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1534_
timestamp 18001
transform -1 0 26864 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1535_
timestamp 18001
transform -1 0 31188 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1536_
timestamp 18001
transform 1 0 27600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1537_
timestamp 18001
transform -1 0 30912 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _1538_
timestamp 18001
transform 1 0 28060 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1539_
timestamp 18001
transform 1 0 31096 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1540_
timestamp 18001
transform 1 0 26220 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1541_
timestamp 18001
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1542_
timestamp 18001
transform 1 0 26864 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1543_
timestamp 18001
transform 1 0 27692 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 18001
transform -1 0 26772 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1545_
timestamp 18001
transform 1 0 30360 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1546_
timestamp 18001
transform 1 0 31004 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1547_
timestamp 18001
transform -1 0 31556 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1548_
timestamp 18001
transform -1 0 31464 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1549_
timestamp 18001
transform -1 0 32292 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1550_
timestamp 18001
transform -1 0 31372 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1551_
timestamp 18001
transform 1 0 31372 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _1552_
timestamp 18001
transform -1 0 30820 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1553_
timestamp 18001
transform -1 0 30544 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1554_
timestamp 18001
transform 1 0 32384 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1555_
timestamp 18001
transform -1 0 33028 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1556_
timestamp 18001
transform 1 0 33028 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1557_
timestamp 18001
transform -1 0 28980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1558_
timestamp 18001
transform 1 0 32016 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1559_
timestamp 18001
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1560_
timestamp 18001
transform -1 0 28244 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1561_
timestamp 18001
transform 1 0 27048 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1562_
timestamp 18001
transform 1 0 27416 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1563_
timestamp 18001
transform -1 0 28336 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1564_
timestamp 18001
transform -1 0 27784 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1565_
timestamp 18001
transform -1 0 26220 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1566_
timestamp 18001
transform 1 0 28152 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1567_
timestamp 18001
transform -1 0 25760 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1568_
timestamp 18001
transform -1 0 27600 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1569_
timestamp 18001
transform -1 0 24656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1570_
timestamp 18001
transform -1 0 21712 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1571_
timestamp 18001
transform 1 0 22724 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 18001
transform -1 0 28244 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _1573_
timestamp 18001
transform 1 0 28428 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1574_
timestamp 18001
transform 1 0 29992 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1575_
timestamp 18001
transform -1 0 29992 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1576_
timestamp 18001
transform 1 0 29808 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1577_
timestamp 18001
transform 1 0 28980 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1578_
timestamp 18001
transform 1 0 26772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1579_
timestamp 18001
transform -1 0 28244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1580_
timestamp 18001
transform 1 0 26036 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1581_
timestamp 18001
transform 1 0 29072 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1582_
timestamp 18001
transform 1 0 28980 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1583_
timestamp 18001
transform 1 0 29624 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1584_
timestamp 18001
transform 1 0 30360 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1585_
timestamp 18001
transform -1 0 32016 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1586_
timestamp 18001
transform 1 0 21620 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1587_
timestamp 18001
transform -1 0 29348 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1588_
timestamp 18001
transform -1 0 28888 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1589_
timestamp 18001
transform -1 0 27416 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1590_
timestamp 18001
transform -1 0 29992 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1591_
timestamp 18001
transform 1 0 27876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1592_
timestamp 18001
transform 1 0 28244 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1593_
timestamp 18001
transform 1 0 25392 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1594_
timestamp 18001
transform -1 0 32016 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _1595_
timestamp 18001
transform -1 0 33580 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1596_
timestamp 18001
transform 1 0 26036 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1597_
timestamp 18001
transform 1 0 27048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1598_
timestamp 18001
transform -1 0 27784 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1599_
timestamp 18001
transform -1 0 30176 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1600_
timestamp 18001
transform -1 0 30176 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1601_
timestamp 18001
transform 1 0 30544 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1602_
timestamp 18001
transform 1 0 26680 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _1603_
timestamp 18001
transform 1 0 30360 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1604_
timestamp 18001
transform 1 0 31188 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1605_
timestamp 18001
transform 1 0 34500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1606_
timestamp 18001
transform 1 0 35144 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_4  _1607_
timestamp 18001
transform -1 0 27692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 18001
transform 1 0 27324 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1609_
timestamp 18001
transform -1 0 29440 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _1610_
timestamp 18001
transform 1 0 28704 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1611_
timestamp 18001
transform -1 0 28704 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1612_
timestamp 18001
transform -1 0 25668 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1613_
timestamp 18001
transform 1 0 25668 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1614_
timestamp 18001
transform 1 0 26036 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1615_
timestamp 18001
transform 1 0 27876 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1616_
timestamp 18001
transform 1 0 25944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1617_
timestamp 18001
transform 1 0 25944 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1618_
timestamp 18001
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1619_
timestamp 18001
transform 1 0 25668 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1620_
timestamp 18001
transform 1 0 33856 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1621_
timestamp 18001
transform 1 0 25668 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1622_
timestamp 18001
transform -1 0 35420 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1623_
timestamp 18001
transform 1 0 28060 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1624_
timestamp 18001
transform 1 0 28428 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 18001
transform 1 0 27876 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1626_
timestamp 18001
transform 1 0 29164 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1627_
timestamp 18001
transform -1 0 29164 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1628_
timestamp 18001
transform 1 0 33764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1629_
timestamp 18001
transform -1 0 34316 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1630_
timestamp 18001
transform 1 0 32384 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1631_
timestamp 18001
transform -1 0 32384 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1632_
timestamp 18001
transform -1 0 32016 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1633_
timestamp 18001
transform 1 0 27508 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1634_
timestamp 18001
transform 1 0 27692 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1635_
timestamp 18001
transform -1 0 29624 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1636_
timestamp 18001
transform 1 0 31556 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1637_
timestamp 18001
transform 1 0 28704 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1638_
timestamp 18001
transform 1 0 26864 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1639_
timestamp 18001
transform 1 0 27048 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1640_
timestamp 18001
transform 1 0 28428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1641_
timestamp 18001
transform 1 0 31648 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1642_
timestamp 18001
transform -1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1643_
timestamp 18001
transform -1 0 31188 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1644_
timestamp 18001
transform 1 0 31188 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1645_
timestamp 18001
transform 1 0 34408 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1646_
timestamp 18001
transform 1 0 26680 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1647_
timestamp 18001
transform 1 0 26956 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 18001
transform 1 0 25484 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1649_
timestamp 18001
transform 1 0 28060 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1650_
timestamp 18001
transform -1 0 26864 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1651_
timestamp 18001
transform 1 0 27232 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1652_
timestamp 18001
transform 1 0 27416 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1653_
timestamp 18001
transform 1 0 27600 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1654_
timestamp 18001
transform 1 0 27508 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1655_
timestamp 18001
transform 1 0 28980 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1656_
timestamp 18001
transform 1 0 29624 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1657_
timestamp 18001
transform 1 0 32292 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1658_
timestamp 18001
transform 1 0 29716 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1659_
timestamp 18001
transform 1 0 33028 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1660_
timestamp 18001
transform -1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1661_
timestamp 18001
transform 1 0 33764 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 18001
transform -1 0 30912 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1663_
timestamp 18001
transform -1 0 27600 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1664_
timestamp 18001
transform 1 0 27232 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1665_
timestamp 18001
transform 1 0 27508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1666_
timestamp 18001
transform 1 0 29532 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1667_
timestamp 18001
transform 1 0 28336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1668_
timestamp 18001
transform 1 0 34592 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1669_
timestamp 18001
transform 1 0 27324 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1670_
timestamp 18001
transform -1 0 30268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1671_
timestamp 18001
transform 1 0 34868 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1672_
timestamp 18001
transform 1 0 35420 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1673_
timestamp 18001
transform -1 0 32844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1674_
timestamp 18001
transform -1 0 33212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 18001
transform 1 0 30636 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1676_
timestamp 18001
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1677_
timestamp 18001
transform -1 0 34500 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1678_
timestamp 18001
transform 1 0 33488 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1679_
timestamp 18001
transform -1 0 32660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1680_
timestamp 18001
transform -1 0 32844 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1681_
timestamp 18001
transform 1 0 34868 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1682_
timestamp 18001
transform 1 0 28520 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1683_
timestamp 18001
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1684_
timestamp 18001
transform -1 0 27968 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1685_
timestamp 18001
transform -1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1686_
timestamp 18001
transform 1 0 33304 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1687_
timestamp 18001
transform -1 0 30820 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1688_
timestamp 18001
transform 1 0 30544 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1689_
timestamp 18001
transform -1 0 30176 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1690_
timestamp 18001
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1691_
timestamp 18001
transform 1 0 32384 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1692_
timestamp 18001
transform 1 0 34684 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1693_
timestamp 18001
transform 1 0 35328 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1694_
timestamp 18001
transform -1 0 30636 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1695_
timestamp 18001
transform -1 0 31280 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1696_
timestamp 18001
transform 1 0 31280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1697_
timestamp 18001
transform -1 0 30360 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1698_
timestamp 18001
transform 1 0 30360 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1699_
timestamp 18001
transform 1 0 29532 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1700_
timestamp 18001
transform 1 0 27784 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1701_
timestamp 18001
transform 1 0 27416 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1702_
timestamp 18001
transform 1 0 28796 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1703_
timestamp 18001
transform -1 0 31740 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1704_
timestamp 18001
transform 1 0 32752 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1705_
timestamp 18001
transform 1 0 33856 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1706_
timestamp 18001
transform -1 0 34132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1707_
timestamp 18001
transform -1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1708_
timestamp 18001
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1709_
timestamp 18001
transform 1 0 32660 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1710_
timestamp 18001
transform -1 0 33580 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1711_
timestamp 18001
transform 1 0 33948 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1712_
timestamp 18001
transform 1 0 34500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1713_
timestamp 18001
transform 1 0 35144 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1714_
timestamp 18001
transform 1 0 33120 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1715_
timestamp 18001
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1716_
timestamp 18001
transform 1 0 32016 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1717_
timestamp 18001
transform 1 0 34132 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1718_
timestamp 18001
transform 1 0 32752 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1719_
timestamp 18001
transform 1 0 27876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1720_
timestamp 18001
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1721_
timestamp 18001
transform 1 0 34500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1722_
timestamp 18001
transform -1 0 32844 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1723_
timestamp 18001
transform 1 0 33304 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1724_
timestamp 18001
transform 1 0 33488 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1725_
timestamp 18001
transform 1 0 31280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1726_
timestamp 18001
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1727_
timestamp 18001
transform 1 0 27508 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1728_
timestamp 18001
transform 1 0 27232 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1729_
timestamp 18001
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1730_
timestamp 18001
transform 1 0 31464 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1731_
timestamp 18001
transform 1 0 30268 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1732_
timestamp 18001
transform -1 0 35236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1733_
timestamp 18001
transform -1 0 30728 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1734_
timestamp 18001
transform 1 0 30268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1735_
timestamp 18001
transform 1 0 32108 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1736_
timestamp 18001
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1737_
timestamp 18001
transform 1 0 16744 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1738_
timestamp 18001
transform 1 0 17296 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1739_
timestamp 18001
transform -1 0 15640 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1740_
timestamp 18001
transform 1 0 17388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_2  _1741_
timestamp 18001
transform 1 0 21068 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1742_
timestamp 18001
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1743_
timestamp 18001
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1744_
timestamp 18001
transform 1 0 14444 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1745_
timestamp 18001
transform 1 0 20884 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1746_
timestamp 18001
transform -1 0 17204 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1747_
timestamp 18001
transform 1 0 16928 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1748_
timestamp 18001
transform 1 0 15824 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1749_
timestamp 18001
transform -1 0 17204 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1750_
timestamp 18001
transform 1 0 15732 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1751_
timestamp 18001
transform -1 0 15364 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1752_
timestamp 18001
transform -1 0 14812 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1753_
timestamp 18001
transform 1 0 17756 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1754_
timestamp 18001
transform -1 0 26588 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1755_
timestamp 18001
transform 1 0 17572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1756_
timestamp 18001
transform 1 0 16560 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1757_
timestamp 18001
transform 1 0 16008 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1758_
timestamp 18001
transform -1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1759_
timestamp 18001
transform 1 0 14260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1760_
timestamp 18001
transform 1 0 14444 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_4  _1761_
timestamp 18001
transform 1 0 19872 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__nand2_2  _1762_
timestamp 18001
transform -1 0 15272 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1763_
timestamp 18001
transform -1 0 17756 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1764_
timestamp 18001
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1765_
timestamp 18001
transform 1 0 14720 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1766_
timestamp 18001
transform -1 0 27140 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1767_
timestamp 18001
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1768_
timestamp 18001
transform 1 0 18308 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1769_
timestamp 18001
transform -1 0 18308 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1770_
timestamp 18001
transform 1 0 17388 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1771_
timestamp 18001
transform -1 0 19044 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1772_
timestamp 18001
transform 1 0 14720 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1773_
timestamp 18001
transform -1 0 15548 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1774_
timestamp 18001
transform -1 0 12512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1775_
timestamp 18001
transform -1 0 11408 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1776_
timestamp 18001
transform -1 0 18492 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1777_
timestamp 18001
transform 1 0 17664 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1778_
timestamp 18001
transform -1 0 20424 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1779_
timestamp 18001
transform -1 0 19964 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1780_
timestamp 18001
transform 1 0 17572 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1781_
timestamp 18001
transform 1 0 17204 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1782_
timestamp 18001
transform 1 0 14076 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1783_
timestamp 18001
transform -1 0 14076 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1784_
timestamp 18001
transform 1 0 17480 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1785_
timestamp 18001
transform 1 0 13892 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1786_
timestamp 18001
transform 1 0 23552 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1787_
timestamp 18001
transform 1 0 12880 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1788_
timestamp 18001
transform -1 0 13156 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1789_
timestamp 18001
transform -1 0 18216 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1790_
timestamp 18001
transform 1 0 14352 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1791_
timestamp 18001
transform -1 0 23460 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1792_
timestamp 18001
transform 1 0 13984 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1793_
timestamp 18001
transform -1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1794_
timestamp 18001
transform -1 0 13064 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1795_
timestamp 18001
transform -1 0 16560 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1796_
timestamp 18001
transform 1 0 15364 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1797_
timestamp 18001
transform 1 0 15088 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1798_
timestamp 18001
transform 1 0 12420 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1799_
timestamp 18001
transform -1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1800_
timestamp 18001
transform 1 0 17756 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1801_
timestamp 18001
transform 1 0 17572 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1802_
timestamp 18001
transform 1 0 17112 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1803_
timestamp 18001
transform 1 0 17296 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1804_
timestamp 18001
transform -1 0 13800 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1805_
timestamp 18001
transform -1 0 26772 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _1806_
timestamp 18001
transform 1 0 25300 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1807_
timestamp 18001
transform 1 0 23184 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1808_
timestamp 18001
transform -1 0 21252 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1809_
timestamp 18001
transform -1 0 21068 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1810_
timestamp 18001
transform 1 0 19412 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1811_
timestamp 18001
transform 1 0 19964 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1812_
timestamp 18001
transform -1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1813_
timestamp 18001
transform 1 0 18676 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1814_
timestamp 18001
transform 1 0 20332 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_2  _1815_
timestamp 18001
transform -1 0 20792 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1816_
timestamp 18001
transform -1 0 15916 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _1817_
timestamp 18001
transform 1 0 22724 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__a211oi_4  _1818_
timestamp 18001
transform 1 0 15088 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1819_
timestamp 18001
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _1820_
timestamp 18001
transform 1 0 18768 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1821_
timestamp 18001
transform -1 0 18032 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1822_
timestamp 18001
transform -1 0 17848 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1823_
timestamp 18001
transform -1 0 15456 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1824_
timestamp 18001
transform -1 0 17664 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1825_
timestamp 18001
transform -1 0 16560 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1826_
timestamp 18001
transform 1 0 17572 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1827_
timestamp 18001
transform 1 0 18400 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1828_
timestamp 18001
transform -1 0 21896 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1829_
timestamp 18001
transform -1 0 20976 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1830_
timestamp 18001
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1831_
timestamp 18001
transform 1 0 20700 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1832_
timestamp 18001
transform -1 0 18400 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1833_
timestamp 18001
transform 1 0 16652 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1834_
timestamp 18001
transform 1 0 17388 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1835_
timestamp 18001
transform 1 0 18308 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1836_
timestamp 18001
transform -1 0 17204 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1837_
timestamp 18001
transform 1 0 16652 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1838_
timestamp 18001
transform 1 0 17388 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1839_
timestamp 18001
transform -1 0 19964 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1840_
timestamp 18001
transform 1 0 18124 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1841_
timestamp 18001
transform -1 0 16560 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1842_
timestamp 18001
transform 1 0 16652 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1843_
timestamp 18001
transform 1 0 17388 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1844_
timestamp 18001
transform -1 0 15272 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1845_
timestamp 18001
transform 1 0 15824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1846_
timestamp 18001
transform -1 0 16376 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _1847_
timestamp 18001
transform -1 0 14536 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_1  _1848_
timestamp 18001
transform 1 0 14352 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1849_
timestamp 18001
transform -1 0 15272 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1850_
timestamp 18001
transform -1 0 26680 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1851_
timestamp 18001
transform -1 0 17756 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1852_
timestamp 18001
transform -1 0 16376 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1853_
timestamp 18001
transform 1 0 12512 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1854_
timestamp 18001
transform -1 0 12696 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1855_
timestamp 18001
transform 1 0 6348 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1856_
timestamp 18001
transform -1 0 14536 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1857_
timestamp 18001
transform -1 0 17296 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1858_
timestamp 18001
transform 1 0 12604 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1859_
timestamp 18001
transform -1 0 15456 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _1860_
timestamp 18001
transform -1 0 16468 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1861_
timestamp 18001
transform -1 0 13708 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1862_
timestamp 18001
transform 1 0 12788 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1863_
timestamp 18001
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1864_
timestamp 18001
transform 1 0 8924 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1865_
timestamp 18001
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1866_
timestamp 18001
transform -1 0 14536 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1867_
timestamp 18001
transform -1 0 16652 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1868_
timestamp 18001
transform -1 0 15640 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1869_
timestamp 18001
transform -1 0 15640 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _1870_
timestamp 18001
transform -1 0 11040 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1871_
timestamp 18001
transform -1 0 10856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1872_
timestamp 18001
transform 1 0 19320 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1873_
timestamp 18001
transform -1 0 12880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1874_
timestamp 18001
transform -1 0 12788 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1875_
timestamp 18001
transform -1 0 12880 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1876_
timestamp 18001
transform 1 0 20608 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1877_
timestamp 18001
transform -1 0 20700 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1878_
timestamp 18001
transform 1 0 19412 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1879_
timestamp 18001
transform 1 0 17940 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1880_
timestamp 18001
transform 1 0 19044 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1881_
timestamp 18001
transform 1 0 19872 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1882_
timestamp 18001
transform 1 0 20976 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1883_
timestamp 18001
transform -1 0 20608 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1884_
timestamp 18001
transform -1 0 19964 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1885_
timestamp 18001
transform 1 0 15548 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1886_
timestamp 18001
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1887_
timestamp 18001
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1888_
timestamp 18001
transform 1 0 24380 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1889_
timestamp 18001
transform 1 0 23000 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1890_
timestamp 18001
transform 1 0 25024 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1891_
timestamp 18001
transform 1 0 24380 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1892_
timestamp 18001
transform -1 0 24564 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1893_
timestamp 18001
transform -1 0 23000 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1894_
timestamp 18001
transform 1 0 17204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1895_
timestamp 18001
transform 1 0 26956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1896_
timestamp 18001
transform -1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1897_
timestamp 18001
transform -1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1898_
timestamp 18001
transform 1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1899_
timestamp 18001
transform -1 0 12420 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1900_
timestamp 18001
transform -1 0 22080 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1901_
timestamp 18001
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1902_
timestamp 18001
transform 1 0 22632 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1903_
timestamp 18001
transform 1 0 26128 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1904_
timestamp 18001
transform 1 0 17756 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1905_
timestamp 18001
transform -1 0 17480 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1906_
timestamp 18001
transform -1 0 12328 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1907_
timestamp 18001
transform -1 0 13248 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1908_
timestamp 18001
transform -1 0 13524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1909_
timestamp 18001
transform 1 0 12328 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _1910_
timestamp 18001
transform 1 0 11500 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_1  _1911_
timestamp 18001
transform 1 0 10304 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1912_
timestamp 18001
transform -1 0 12052 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _1913_
timestamp 18001
transform -1 0 11132 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1914_
timestamp 18001
transform 1 0 12788 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1915_
timestamp 18001
transform 1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1916_
timestamp 18001
transform -1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1917_
timestamp 18001
transform -1 0 8648 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1918_
timestamp 18001
transform 1 0 8188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1919_
timestamp 18001
transform 1 0 8188 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1920_
timestamp 18001
transform 1 0 8464 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1921_
timestamp 18001
transform 1 0 24748 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1922_
timestamp 18001
transform 1 0 24288 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1923_
timestamp 18001
transform 1 0 24012 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1924_
timestamp 18001
transform 1 0 23736 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1925_
timestamp 18001
transform 1 0 23000 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1926_
timestamp 18001
transform -1 0 24380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1927_
timestamp 18001
transform 1 0 25024 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1928_
timestamp 18001
transform 1 0 22540 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1929_
timestamp 18001
transform -1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1930_
timestamp 18001
transform -1 0 25116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1931_
timestamp 18001
transform -1 0 24104 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1932_
timestamp 18001
transform -1 0 23920 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1933_
timestamp 18001
transform 1 0 23828 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1934_
timestamp 18001
transform -1 0 25024 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1935_
timestamp 18001
transform -1 0 24288 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1936_
timestamp 18001
transform -1 0 23276 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1937_
timestamp 18001
transform 1 0 23092 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1938_
timestamp 18001
transform -1 0 23184 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1939_
timestamp 18001
transform 1 0 19872 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1940_
timestamp 18001
transform 1 0 19228 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1941_
timestamp 18001
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1942_
timestamp 18001
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1943_
timestamp 18001
transform -1 0 16652 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1944_
timestamp 18001
transform 1 0 16836 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _1945_
timestamp 18001
transform 1 0 17940 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1946_
timestamp 18001
transform 1 0 19780 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1947_
timestamp 18001
transform 1 0 20240 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1948_
timestamp 18001
transform -1 0 21528 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1949_
timestamp 18001
transform 1 0 20608 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1950_
timestamp 18001
transform 1 0 20608 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1951_
timestamp 18001
transform 1 0 20884 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1952_
timestamp 18001
transform -1 0 22356 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1953_
timestamp 18001
transform -1 0 21252 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_8  _1954_
timestamp 18001
transform -1 0 16284 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_4  _1955_
timestamp 18001
transform -1 0 14812 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1956_
timestamp 18001
transform -1 0 15916 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1957_
timestamp 18001
transform -1 0 23368 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1958_
timestamp 18001
transform -1 0 16192 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1959_
timestamp 18001
transform 1 0 17204 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1960_
timestamp 18001
transform 1 0 16836 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_4  _1961_
timestamp 18001
transform 1 0 13064 0 -1 28288
box -38 -48 1786 592
use sky130_fd_sc_hd__a221oi_2  _1962_
timestamp 18001
transform 1 0 12880 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _1963_
timestamp 18001
transform -1 0 8832 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1964_
timestamp 18001
transform 1 0 8924 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1965_
timestamp 18001
transform 1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1966_
timestamp 18001
transform -1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1967_
timestamp 18001
transform -1 0 13708 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1968_
timestamp 18001
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1969_
timestamp 18001
transform 1 0 12328 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1970_
timestamp 18001
transform 1 0 15364 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1971_
timestamp 18001
transform -1 0 15364 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1972_
timestamp 18001
transform 1 0 14076 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1973_
timestamp 18001
transform 1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1974_
timestamp 18001
transform 1 0 12236 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1975_
timestamp 18001
transform 1 0 14076 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1976_
timestamp 18001
transform -1 0 14168 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1977_
timestamp 18001
transform 1 0 16652 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1978_
timestamp 18001
transform -1 0 14444 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1979_
timestamp 18001
transform 1 0 13064 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1980_
timestamp 18001
transform -1 0 11592 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1981_
timestamp 18001
transform 1 0 8924 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1982_
timestamp 18001
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1983_
timestamp 18001
transform -1 0 16008 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _1984_
timestamp 18001
transform 1 0 8004 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1985_
timestamp 18001
transform 1 0 15364 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1986_
timestamp 18001
transform 1 0 14812 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1987_
timestamp 18001
transform 1 0 19688 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1988_
timestamp 18001
transform -1 0 19688 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1989_
timestamp 18001
transform 1 0 19228 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1990_
timestamp 18001
transform 1 0 15456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1991_
timestamp 18001
transform 1 0 19228 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1992_
timestamp 18001
transform 1 0 18216 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1993_
timestamp 18001
transform 1 0 19780 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1994_
timestamp 18001
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1995_
timestamp 18001
transform -1 0 18676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1996_
timestamp 18001
transform -1 0 19780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1997_
timestamp 18001
transform -1 0 19228 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1998_
timestamp 18001
transform -1 0 13800 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1999_
timestamp 18001
transform 1 0 14352 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2000_
timestamp 18001
transform -1 0 21160 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2001_
timestamp 18001
transform -1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _2002_
timestamp 18001
transform 1 0 19320 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2003_
timestamp 18001
transform 1 0 12972 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _2004_
timestamp 18001
transform -1 0 13892 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _2005_
timestamp 18001
transform -1 0 13892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2006_
timestamp 18001
transform -1 0 13340 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2007_
timestamp 18001
transform -1 0 14352 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _2008_
timestamp 18001
transform -1 0 12880 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _2009_
timestamp 18001
transform -1 0 11500 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2010_
timestamp 18001
transform -1 0 8832 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _2011_
timestamp 18001
transform -1 0 12972 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2012_
timestamp 18001
transform 1 0 7820 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2013_
timestamp 18001
transform 1 0 9384 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2014_
timestamp 18001
transform -1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2015_
timestamp 18001
transform 1 0 7912 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2016_
timestamp 18001
transform -1 0 8004 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2017_
timestamp 18001
transform 1 0 7636 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2018_
timestamp 18001
transform -1 0 8832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2019_
timestamp 18001
transform -1 0 7176 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2020_
timestamp 18001
transform 1 0 9476 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2021_
timestamp 18001
transform -1 0 10764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2022_
timestamp 18001
transform 1 0 6624 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2023_
timestamp 18001
transform -1 0 6348 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2024_
timestamp 18001
transform 1 0 5428 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2025_
timestamp 18001
transform 1 0 4600 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2026_
timestamp 18001
transform 1 0 2576 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2027_
timestamp 18001
transform -1 0 5428 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _2028_
timestamp 18001
transform 1 0 12052 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _2029_
timestamp 18001
transform 1 0 4140 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _2030_
timestamp 18001
transform 1 0 4232 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2031_
timestamp 18001
transform 1 0 5612 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2032_
timestamp 18001
transform 1 0 4876 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2033_
timestamp 18001
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2034_
timestamp 18001
transform -1 0 6256 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _2035_
timestamp 18001
transform -1 0 6624 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2036_
timestamp 18001
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2037_
timestamp 18001
transform -1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2038_
timestamp 18001
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2039_
timestamp 18001
transform 1 0 6164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _2040_
timestamp 18001
transform 1 0 6716 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _2041_
timestamp 18001
transform -1 0 7268 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2042_
timestamp 18001
transform -1 0 7268 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2043_
timestamp 18001
transform 1 0 6716 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2044_
timestamp 18001
transform 1 0 5428 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2045_
timestamp 18001
transform 1 0 8924 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _2046_
timestamp 18001
transform 1 0 12144 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _2047_
timestamp 18001
transform 1 0 7176 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2048_
timestamp 18001
transform 1 0 8372 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2049_
timestamp 18001
transform 1 0 9200 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2050_
timestamp 18001
transform 1 0 9844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2051_
timestamp 18001
transform -1 0 8556 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2052_
timestamp 18001
transform -1 0 8004 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2053_
timestamp 18001
transform 1 0 7360 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _2054_
timestamp 18001
transform 1 0 6900 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2055_
timestamp 18001
transform -1 0 6072 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2056_
timestamp 18001
transform 1 0 7360 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2057_
timestamp 18001
transform 1 0 6808 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2058_
timestamp 18001
transform -1 0 6348 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2059_
timestamp 18001
transform 1 0 6348 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2060_
timestamp 18001
transform 1 0 7084 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2061_
timestamp 18001
transform -1 0 7084 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2062_
timestamp 18001
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _2063_
timestamp 18001
transform -1 0 5888 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2064_
timestamp 18001
transform -1 0 5704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2065_
timestamp 18001
transform -1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2066_
timestamp 18001
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2067_
timestamp 18001
transform 1 0 4048 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2068_
timestamp 18001
transform 1 0 3956 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _2069_
timestamp 18001
transform -1 0 5244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_2  _2070_
timestamp 18001
transform 1 0 12144 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _2071_
timestamp 18001
transform 1 0 5704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2072_
timestamp 18001
transform 1 0 8740 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2073_
timestamp 18001
transform 1 0 15916 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _2074_
timestamp 18001
transform 1 0 14904 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2075_
timestamp 18001
transform -1 0 14904 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _2076_
timestamp 18001
transform -1 0 6992 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2077_
timestamp 18001
transform -1 0 5888 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2078_
timestamp 18001
transform 1 0 4600 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2079_
timestamp 18001
transform -1 0 5244 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _2080_
timestamp 18001
transform -1 0 5796 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2081_
timestamp 18001
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2082_
timestamp 18001
transform 1 0 6532 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2083_
timestamp 18001
transform -1 0 5796 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2084_
timestamp 18001
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2085_
timestamp 18001
transform 1 0 5796 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2086_
timestamp 18001
transform -1 0 5796 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2087_
timestamp 18001
transform -1 0 6256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2088_
timestamp 18001
transform -1 0 5244 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2089_
timestamp 18001
transform 1 0 4416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2090_
timestamp 18001
transform 1 0 6348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2091_
timestamp 18001
transform -1 0 4600 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2092_
timestamp 18001
transform 1 0 3864 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2093_
timestamp 18001
transform 1 0 3588 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2094_
timestamp 18001
transform -1 0 4968 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2095_
timestamp 18001
transform 1 0 5244 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _2096_
timestamp 18001
transform 1 0 13156 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__o22ai_1  _2097_
timestamp 18001
transform -1 0 8188 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2098_
timestamp 18001
transform 1 0 9108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2099_
timestamp 18001
transform -1 0 10028 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2100_
timestamp 18001
transform -1 0 7360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2101_
timestamp 18001
transform -1 0 7176 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2102_
timestamp 18001
transform 1 0 6532 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _2103_
timestamp 18001
transform 1 0 6624 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2104_
timestamp 18001
transform -1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2105_
timestamp 18001
transform 1 0 6808 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2106_
timestamp 18001
transform 1 0 5152 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2107_
timestamp 18001
transform 1 0 5612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2108_
timestamp 18001
transform -1 0 6072 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2109_
timestamp 18001
transform 1 0 5612 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2110_
timestamp 18001
transform 1 0 5888 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_1  _2111_
timestamp 18001
transform 1 0 4968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2112_
timestamp 18001
transform 1 0 12328 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2113_
timestamp 18001
transform 1 0 12972 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2114_
timestamp 18001
transform -1 0 9108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _2115_
timestamp 18001
transform 1 0 7360 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2116_
timestamp 18001
transform 1 0 4508 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2117_
timestamp 18001
transform 1 0 2944 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2118_
timestamp 18001
transform 1 0 3772 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _2119_
timestamp 18001
transform 1 0 4140 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__a221oi_2  _2120_
timestamp 18001
transform 1 0 11776 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _2121_
timestamp 18001
transform 1 0 7084 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2122_
timestamp 18001
transform 1 0 6900 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _2123_
timestamp 18001
transform 1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _2124_
timestamp 18001
transform -1 0 8096 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2125_
timestamp 18001
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2126_
timestamp 18001
transform 1 0 7820 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2127_
timestamp 18001
transform 1 0 7912 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2128_
timestamp 18001
transform -1 0 12880 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2129_
timestamp 18001
transform -1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _2130_
timestamp 18001
transform 1 0 8556 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2131_
timestamp 18001
transform 1 0 8280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2132_
timestamp 18001
transform -1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2133_
timestamp 18001
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2134_
timestamp 18001
transform 1 0 11040 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _2135_
timestamp 18001
transform -1 0 11960 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2136_
timestamp 18001
transform -1 0 11408 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2137_
timestamp 18001
transform -1 0 11316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2138_
timestamp 18001
transform -1 0 12052 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2139_
timestamp 18001
transform 1 0 10764 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2140_
timestamp 18001
transform -1 0 12144 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2141_
timestamp 18001
transform -1 0 11960 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _2142_
timestamp 18001
transform 1 0 12052 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__o2bb2a_1  _2143_
timestamp 18001
transform 1 0 10948 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _2144_
timestamp 18001
transform 1 0 10764 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2145_
timestamp 18001
transform -1 0 9568 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _2146_
timestamp 18001
transform -1 0 12328 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2147_
timestamp 18001
transform -1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2148_
timestamp 18001
transform 1 0 10304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2149_
timestamp 18001
transform 1 0 12052 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2150_
timestamp 18001
transform -1 0 11960 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2151_
timestamp 18001
transform 1 0 11316 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _2152_
timestamp 18001
transform -1 0 12328 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2153_
timestamp 18001
transform 1 0 10212 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2154_
timestamp 18001
transform 1 0 9476 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2155_
timestamp 18001
transform 1 0 10120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2156_
timestamp 18001
transform 1 0 10304 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _2157_
timestamp 18001
transform 1 0 8924 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _2158_
timestamp 18001
transform -1 0 9660 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2159_
timestamp 18001
transform 1 0 9936 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2160_
timestamp 18001
transform -1 0 9476 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2161_
timestamp 18001
transform 1 0 14260 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _2162_
timestamp 18001
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2163_
timestamp 18001
transform 1 0 13248 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2164_
timestamp 18001
transform 1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2165_
timestamp 18001
transform 1 0 11408 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _2166_
timestamp 18001
transform 1 0 10580 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _2167_
timestamp 18001
transform 1 0 12236 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2168_
timestamp 18001
transform 1 0 11500 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2169_
timestamp 18001
transform -1 0 10488 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _2170_
timestamp 18001
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _2171_
timestamp 18001
transform -1 0 9936 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2172_
timestamp 18001
transform -1 0 10304 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2173_
timestamp 18001
transform 1 0 10764 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2174_
timestamp 18001
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2175_
timestamp 18001
transform 1 0 9016 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _2176_
timestamp 18001
transform -1 0 10580 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2177_
timestamp 18001
transform -1 0 11408 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  _2178_
timestamp 18001
transform 1 0 11500 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2179_
timestamp 18001
transform -1 0 14260 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _2180_
timestamp 18001
transform 1 0 12144 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2181_
timestamp 18001
transform 1 0 11776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2182_
timestamp 18001
transform -1 0 10764 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2183_
timestamp 18001
transform 1 0 9660 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2184_
timestamp 18001
transform 1 0 8188 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2185_
timestamp 18001
transform -1 0 9752 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _2186_
timestamp 18001
transform 1 0 8740 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2187_
timestamp 18001
transform -1 0 16100 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2188_
timestamp 18001
transform 1 0 15824 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2189_
timestamp 18001
transform 1 0 15456 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2190_
timestamp 18001
transform -1 0 18860 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2191_
timestamp 18001
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2192_
timestamp 18001
transform -1 0 17020 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2193_
timestamp 18001
transform 1 0 15916 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2194_
timestamp 18001
transform 1 0 15916 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2195_
timestamp 18001
transform 1 0 15824 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2196_
timestamp 18001
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2197_
timestamp 18001
transform -1 0 13432 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2198_
timestamp 18001
transform 1 0 9752 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _2199_
timestamp 18001
transform -1 0 10120 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _2200_
timestamp 18001
transform 1 0 7912 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2201_
timestamp 18001
transform 1 0 7360 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2202_
timestamp 18001
transform 1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2203_
timestamp 18001
transform 1 0 5888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2204_
timestamp 18001
transform -1 0 5980 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _2205_
timestamp 18001
transform 1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2206_
timestamp 18001
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2207_
timestamp 18001
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2208_
timestamp 18001
transform -1 0 4784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2209_
timestamp 18001
transform 1 0 4324 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2210_
timestamp 18001
transform -1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2211_
timestamp 18001
transform 1 0 7544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2212_
timestamp 18001
transform -1 0 7636 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2213_
timestamp 18001
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2214_
timestamp 18001
transform 1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _2215_
timestamp 18001
transform -1 0 10580 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _2216_
timestamp 18001
transform -1 0 10488 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_2  _2217_
timestamp 18001
transform 1 0 17296 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2218_
timestamp 18001
transform -1 0 5888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2219_
timestamp 18001
transform 1 0 7544 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2220_
timestamp 18001
transform 1 0 7176 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2221_
timestamp 18001
transform -1 0 7636 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2222_
timestamp 18001
transform -1 0 8832 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2223_
timestamp 18001
transform 1 0 2760 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2224_
timestamp 18001
transform -1 0 5060 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2225_
timestamp 18001
transform -1 0 3496 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2226_
timestamp 18001
transform -1 0 5152 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2227_
timestamp 18001
transform -1 0 2852 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2228_
timestamp 18001
transform -1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2229_
timestamp 18001
transform -1 0 5796 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2230_
timestamp 18001
transform 1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2231_
timestamp 18001
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2232_
timestamp 18001
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2233_
timestamp 18001
transform -1 0 4600 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2234_
timestamp 18001
transform 1 0 5888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2235_
timestamp 18001
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2236_
timestamp 18001
transform -1 0 8464 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2237_
timestamp 18001
transform 1 0 5612 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2238_
timestamp 18001
transform 1 0 6348 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2239_
timestamp 18001
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2240_
timestamp 18001
transform -1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2241_
timestamp 18001
transform -1 0 12880 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2242_
timestamp 18001
transform 1 0 18124 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2243_
timestamp 18001
transform -1 0 13984 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2244_
timestamp 18001
transform 1 0 12144 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2245_
timestamp 18001
transform 1 0 12236 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2246_
timestamp 18001
transform -1 0 11408 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2247_
timestamp 18001
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2248_
timestamp 18001
transform 1 0 19136 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _2249_
timestamp 18001
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _2250_
timestamp 18001
transform 1 0 19228 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2251_
timestamp 18001
transform -1 0 11408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2252_
timestamp 18001
transform 1 0 11592 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2253_
timestamp 18001
transform 1 0 9016 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _2254_
timestamp 18001
transform 1 0 10028 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _2255_
timestamp 18001
transform 1 0 10580 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2256_
timestamp 18001
transform -1 0 12420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _2257_
timestamp 18001
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _2258_
timestamp 18001
transform -1 0 18124 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2259_
timestamp 18001
transform -1 0 13432 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2260_
timestamp 18001
transform -1 0 11776 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _2261_
timestamp 18001
transform 1 0 26772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2262_
timestamp 18001
transform -1 0 12052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _2263_
timestamp 18001
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2264_
timestamp 18001
transform 1 0 7268 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2265_
timestamp 18001
transform -1 0 9752 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2266_
timestamp 18001
transform 1 0 9844 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2267_
timestamp 18001
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _2268_
timestamp 18001
transform -1 0 12328 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2269_
timestamp 18001
transform -1 0 15548 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2270_
timestamp 18001
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2271_
timestamp 18001
transform 1 0 9936 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2272_
timestamp 18001
transform -1 0 21712 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2273_
timestamp 18001
transform -1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2274_
timestamp 18001
transform 1 0 11960 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2275_
timestamp 18001
transform 1 0 13156 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2276_
timestamp 18001
transform -1 0 15640 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2277_
timestamp 18001
transform 1 0 15088 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2278_
timestamp 18001
transform 1 0 19320 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2279_
timestamp 18001
transform -1 0 15824 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2280_
timestamp 18001
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2281_
timestamp 18001
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2282_
timestamp 18001
transform 1 0 12788 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _2283_
timestamp 18001
transform 1 0 18308 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2284_
timestamp 18001
transform -1 0 17940 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2285_
timestamp 18001
transform -1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2286_
timestamp 18001
transform 1 0 15916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2287_
timestamp 18001
transform -1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2288_
timestamp 18001
transform -1 0 17940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2289_
timestamp 18001
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2290_
timestamp 18001
transform 1 0 15180 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _2291_
timestamp 18001
transform 1 0 14904 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2292_
timestamp 18001
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2293_
timestamp 18001
transform -1 0 11592 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2294_
timestamp 18001
transform -1 0 9476 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2295_
timestamp 18001
transform 1 0 10304 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2296_
timestamp 18001
transform -1 0 8832 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2297_
timestamp 18001
transform 1 0 9016 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2298_
timestamp 18001
transform 1 0 9476 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2299_
timestamp 18001
transform 1 0 11868 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _2300_
timestamp 18001
transform 1 0 20148 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2301_
timestamp 18001
transform 1 0 20884 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2302_
timestamp 18001
transform 1 0 20056 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2303_
timestamp 18001
transform 1 0 20148 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2304_
timestamp 18001
transform 1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2305_
timestamp 18001
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2306_
timestamp 18001
transform -1 0 20424 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2307_
timestamp 18001
transform -1 0 23828 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2308_
timestamp 18001
transform 1 0 22632 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _2309_
timestamp 18001
transform -1 0 24932 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _2310_
timestamp 18001
transform 1 0 21160 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2311_
timestamp 18001
transform 1 0 22080 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2312_
timestamp 18001
transform -1 0 22632 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2313_
timestamp 18001
transform -1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2314_
timestamp 18001
transform 1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2315_
timestamp 18001
transform -1 0 20516 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2316_
timestamp 18001
transform 1 0 19872 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2317_
timestamp 18001
transform 1 0 18216 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2318_
timestamp 18001
transform 1 0 17664 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _2319_
timestamp 18001
transform -1 0 18952 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2320_
timestamp 18001
transform 1 0 19228 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2321_
timestamp 18001
transform -1 0 19044 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _2322_
timestamp 18001
transform 1 0 18860 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2323_
timestamp 18001
transform 1 0 13984 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2324_
timestamp 18001
transform 1 0 14076 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _2325_
timestamp 18001
transform -1 0 18768 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2326_
timestamp 18001
transform 1 0 8556 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2327_
timestamp 18001
transform 1 0 9016 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2328_
timestamp 18001
transform 1 0 8832 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2329_
timestamp 18001
transform 1 0 8924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2330_
timestamp 18001
transform 1 0 8740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2331_
timestamp 18001
transform 1 0 7452 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2332_
timestamp 18001
transform -1 0 6072 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2333_
timestamp 18001
transform 1 0 7176 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2334_
timestamp 18001
transform 1 0 7452 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2335_
timestamp 18001
transform -1 0 7728 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2336_
timestamp 18001
transform 1 0 7728 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2337_
timestamp 18001
transform -1 0 7268 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2338_
timestamp 18001
transform -1 0 7544 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2339_
timestamp 18001
transform 1 0 7820 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2340_
timestamp 18001
transform 1 0 7084 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2341_
timestamp 18001
transform -1 0 8188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2342_
timestamp 18001
transform -1 0 8464 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2343_
timestamp 18001
transform -1 0 8740 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2344_
timestamp 18001
transform -1 0 9200 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2345_
timestamp 18001
transform -1 0 9476 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2346_
timestamp 18001
transform -1 0 11040 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2347_
timestamp 18001
transform 1 0 11500 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2348_
timestamp 18001
transform -1 0 12604 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2349_
timestamp 18001
transform 1 0 9568 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2350_
timestamp 18001
transform 1 0 7636 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2351_
timestamp 18001
transform 1 0 7084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2352_
timestamp 18001
transform -1 0 7452 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2353_
timestamp 18001
transform 1 0 6900 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2354_
timestamp 18001
transform -1 0 8740 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2355_
timestamp 18001
transform -1 0 9752 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2356_
timestamp 18001
transform 1 0 9292 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2357_
timestamp 18001
transform 1 0 9660 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _2358_
timestamp 18001
transform 1 0 9752 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2359_
timestamp 18001
transform -1 0 6992 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2360_
timestamp 18001
transform 1 0 5612 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2361_
timestamp 18001
transform 1 0 6532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _2362_
timestamp 18001
transform 1 0 14536 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _2363_
timestamp 18001
transform 1 0 6348 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2364_
timestamp 18001
transform 1 0 6716 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2365_
timestamp 18001
transform -1 0 9476 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2366_
timestamp 18001
transform 1 0 9476 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2367_
timestamp 18001
transform 1 0 9108 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _2368_
timestamp 18001
transform -1 0 5520 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2369_
timestamp 18001
transform -1 0 5060 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2370_
timestamp 18001
transform 1 0 4324 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2371_
timestamp 18001
transform 1 0 9292 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2372_
timestamp 18001
transform -1 0 10396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2373_
timestamp 18001
transform 1 0 11776 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2374_
timestamp 18001
transform 1 0 9384 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2375_
timestamp 18001
transform 1 0 9844 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _2376_
timestamp 18001
transform -1 0 14996 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2377_
timestamp 18001
transform -1 0 11316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2378_
timestamp 18001
transform 1 0 9752 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2379_
timestamp 18001
transform -1 0 10580 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2380_
timestamp 18001
transform 1 0 10580 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2381_
timestamp 18001
transform 1 0 10672 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2382_
timestamp 18001
transform 1 0 11040 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _2383_
timestamp 18001
transform 1 0 11684 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_4  _2384_
timestamp 18001
transform -1 0 13064 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_1  _2385_
timestamp 18001
transform 1 0 9936 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2386_
timestamp 18001
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2387_
timestamp 18001
transform 1 0 11316 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2388_
timestamp 18001
transform -1 0 12052 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2389_
timestamp 18001
transform 1 0 11500 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2390_
timestamp 18001
transform -1 0 13984 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2391_
timestamp 18001
transform -1 0 13800 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2392_
timestamp 18001
transform 1 0 12052 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2393_
timestamp 18001
transform -1 0 14352 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2394_
timestamp 18001
transform -1 0 13432 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2395_
timestamp 18001
transform 1 0 14352 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2396_
timestamp 18001
transform 1 0 12328 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2397_
timestamp 18001
transform 1 0 10948 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2398_
timestamp 18001
transform -1 0 12972 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2399_
timestamp 18001
transform -1 0 8188 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _2400_
timestamp 18001
transform 1 0 7176 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _2401_
timestamp 18001
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2402_
timestamp 18001
transform -1 0 12788 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2403_
timestamp 18001
transform -1 0 13340 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2404_
timestamp 18001
transform 1 0 12236 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2405_
timestamp 18001
transform -1 0 13156 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2406_
timestamp 18001
transform 1 0 12972 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2407_
timestamp 18001
transform -1 0 15272 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_1  _2408_
timestamp 18001
transform 1 0 10672 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2409_
timestamp 18001
transform -1 0 14996 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2410_
timestamp 18001
transform -1 0 7728 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _2411_
timestamp 18001
transform 1 0 7176 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2412_
timestamp 18001
transform 1 0 16192 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2413_
timestamp 18001
transform 1 0 14996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2414_
timestamp 18001
transform -1 0 13616 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2415_
timestamp 18001
transform 1 0 13616 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2416_
timestamp 18001
transform 1 0 14720 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2417_
timestamp 18001
transform -1 0 15824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2418_
timestamp 18001
transform -1 0 15088 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2419_
timestamp 18001
transform 1 0 15824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2420_
timestamp 18001
transform 1 0 12788 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _2421_
timestamp 18001
transform 1 0 14076 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2422_
timestamp 18001
transform -1 0 13800 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2423_
timestamp 18001
transform 1 0 14076 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2424_
timestamp 18001
transform 1 0 15824 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2425_
timestamp 18001
transform 1 0 15180 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2426_
timestamp 18001
transform 1 0 4876 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_4  _2427_
timestamp 18001
transform 1 0 4876 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  _2428_
timestamp 18001
transform 1 0 21344 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _2429_
timestamp 18001
transform 1 0 14904 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2430_
timestamp 18001
transform -1 0 15824 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2431_
timestamp 18001
transform 1 0 15088 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _2432_
timestamp 18001
transform 1 0 15180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2433_
timestamp 18001
transform 1 0 17388 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2434_
timestamp 18001
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2435_
timestamp 18001
transform 1 0 17296 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2436_
timestamp 18001
transform 1 0 15916 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2437_
timestamp 18001
transform 1 0 8556 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _2438_
timestamp 18001
transform -1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2439_
timestamp 18001
transform 1 0 15916 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2440_
timestamp 18001
transform 1 0 15272 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2441_
timestamp 18001
transform 1 0 16008 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2442_
timestamp 18001
transform -1 0 14904 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2443_
timestamp 18001
transform 1 0 16652 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2444_
timestamp 18001
transform 1 0 16652 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2445_
timestamp 18001
transform 1 0 17296 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2446_
timestamp 18001
transform 1 0 16652 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2447_
timestamp 18001
transform -1 0 19136 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2448_
timestamp 18001
transform 1 0 17572 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2449_
timestamp 18001
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2450_
timestamp 18001
transform -1 0 18308 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2451_
timestamp 18001
transform -1 0 5612 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _2452_
timestamp 18001
transform -1 0 6348 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2453_
timestamp 18001
transform -1 0 19136 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2454_
timestamp 18001
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2455_
timestamp 18001
transform 1 0 18032 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _2456_
timestamp 18001
transform 1 0 17112 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2457_
timestamp 18001
transform 1 0 16284 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2458_
timestamp 18001
transform 1 0 16928 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _2459_
timestamp 18001
transform 1 0 18584 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2460_
timestamp 18001
transform 1 0 19136 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2461_
timestamp 18001
transform 1 0 8924 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2462_
timestamp 18001
transform 1 0 8648 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _2463_
timestamp 18001
transform 1 0 17756 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2464_
timestamp 18001
transform -1 0 19044 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2465_
timestamp 18001
transform 1 0 17848 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _2466_
timestamp 18001
transform 1 0 20516 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_4  _2467_
timestamp 18001
transform 1 0 19228 0 1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2468_
timestamp 18001
transform 1 0 8924 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2469_
timestamp 18001
transform 1 0 9752 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2470_
timestamp 18001
transform 1 0 2300 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2471_
timestamp 18001
transform 1 0 1748 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2472_
timestamp 18001
transform 1 0 3772 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2473_
timestamp 18001
transform 1 0 6256 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2474_
timestamp 18001
transform 1 0 2116 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2475_
timestamp 18001
transform 1 0 7360 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _2476_
timestamp 18001
transform 1 0 26312 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2477_
timestamp 18001
transform -1 0 23644 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _2478_
timestamp 18001
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2479_
timestamp 18001
transform 1 0 9016 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2480_
timestamp 18001
transform 1 0 10212 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2481_
timestamp 18001
transform 1 0 2024 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2482_
timestamp 18001
transform 1 0 2024 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2483_
timestamp 18001
transform 1 0 3220 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2484_
timestamp 18001
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2485_
timestamp 18001
transform 1 0 1932 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2486_
timestamp 18001
transform 1 0 6716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2487_
timestamp 18001
transform 1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2488_
timestamp 18001
transform 1 0 18032 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_1  _2489_
timestamp 18001
transform 1 0 22816 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _2490_
timestamp 18001
transform -1 0 21804 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2491_
timestamp 18001
transform 1 0 24288 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2492_
timestamp 18001
transform 1 0 23092 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2493_
timestamp 18001
transform 1 0 23552 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2494_
timestamp 18001
transform -1 0 23552 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2495_
timestamp 18001
transform -1 0 20700 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2496_
timestamp 18001
transform 1 0 20516 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2497_
timestamp 18001
transform -1 0 20332 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _2498_
timestamp 18001
transform 1 0 18584 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _2499_
timestamp 18001
transform 1 0 19780 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2500_
timestamp 18001
transform 1 0 20516 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2501_
timestamp 18001
transform 1 0 21988 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2502_
timestamp 18001
transform 1 0 25208 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2503_
timestamp 18001
transform 1 0 23092 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 18001
transform 1 0 24380 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2505_
timestamp 18001
transform 1 0 20148 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 18001
transform 1 0 22816 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2507_
timestamp 18001
transform 1 0 24472 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2508_
timestamp 18001
transform 1 0 13156 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2509_
timestamp 18001
transform 1 0 13064 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2510_
timestamp 18001
transform -1 0 10764 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2511_
timestamp 18001
transform 1 0 10488 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2512_
timestamp 18001
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2513_
timestamp 18001
transform -1 0 11592 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2514_
timestamp 18001
transform -1 0 11408 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2515_
timestamp 18001
transform 1 0 11592 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2516_
timestamp 18001
transform -1 0 11500 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2517_
timestamp 18001
transform 1 0 10120 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2518_
timestamp 18001
transform 1 0 9200 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2519_
timestamp 18001
transform -1 0 10120 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2520_
timestamp 18001
transform 1 0 10120 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2521_
timestamp 18001
transform 1 0 9568 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2522_
timestamp 18001
transform 1 0 9016 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2523_
timestamp 18001
transform -1 0 6072 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2524_
timestamp 18001
transform -1 0 8556 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2525_
timestamp 18001
transform 1 0 7544 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2526_
timestamp 18001
transform 1 0 5520 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2527_
timestamp 18001
transform 1 0 5520 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2528_
timestamp 18001
transform 1 0 4784 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2529_
timestamp 18001
transform 1 0 7544 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2530_
timestamp 18001
transform 1 0 6900 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2531_
timestamp 18001
transform 1 0 5060 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2532_
timestamp 18001
transform -1 0 6348 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2533_
timestamp 18001
transform 1 0 6348 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2534_
timestamp 18001
transform -1 0 4600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2535_
timestamp 18001
transform 1 0 4508 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2536_
timestamp 18001
transform 1 0 6348 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2537_
timestamp 18001
transform 1 0 6348 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2538_
timestamp 18001
transform 1 0 4784 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2539_
timestamp 18001
transform -1 0 5336 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _2540_
timestamp 18001
transform -1 0 5888 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2541_
timestamp 18001
transform -1 0 6256 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _2542_
timestamp 18001
transform -1 0 7636 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2543_
timestamp 18001
transform -1 0 5888 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _2544_
timestamp 18001
transform -1 0 7452 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _2545_
timestamp 18001
transform 1 0 6532 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2546_
timestamp 18001
transform 1 0 3956 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2547_
timestamp 18001
transform -1 0 6900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2548_
timestamp 18001
transform -1 0 6532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2549_
timestamp 18001
transform 1 0 6348 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2550_
timestamp 18001
transform -1 0 6992 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2551_
timestamp 18001
transform -1 0 6256 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2552_
timestamp 18001
transform -1 0 6808 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2553_
timestamp 18001
transform -1 0 8188 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2554_
timestamp 18001
transform -1 0 8832 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2555_
timestamp 18001
transform -1 0 7820 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2556_
timestamp 18001
transform 1 0 8004 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2557_
timestamp 18001
transform 1 0 8372 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2558_
timestamp 18001
transform 1 0 7820 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2559_
timestamp 18001
transform 1 0 24932 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2560_
timestamp 18001
transform 1 0 25484 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _2561_
timestamp 18001
transform -1 0 21804 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2562_
timestamp 18001
transform 1 0 7912 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2563_
timestamp 18001
transform 1 0 9844 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2564_
timestamp 18001
transform 1 0 4416 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2565_
timestamp 18001
transform 1 0 2208 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2566_
timestamp 18001
transform 1 0 4784 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2567_
timestamp 18001
transform 1 0 4784 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2568_
timestamp 18001
transform 1 0 1748 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2569_
timestamp 18001
transform 1 0 3772 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2570_
timestamp 18001
transform -1 0 22356 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2571_
timestamp 18001
transform 1 0 21804 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2572_
timestamp 18001
transform 1 0 23460 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _2573_
timestamp 18001
transform -1 0 23460 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2574_
timestamp 18001
transform 1 0 21252 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _2575_
timestamp 18001
transform -1 0 20516 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a221oi_1  _2576_
timestamp 18001
transform 1 0 18768 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _2577_
timestamp 18001
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2578_
timestamp 18001
transform 1 0 3772 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2579_
timestamp 18001
transform 1 0 3864 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2580_
timestamp 18001
transform 1 0 2208 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2581_
timestamp 18001
transform 1 0 3772 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2582_
timestamp 18001
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2583_
timestamp 18001
transform 1 0 3128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2584_
timestamp 18001
transform 1 0 1840 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2585_
timestamp 18001
transform 1 0 2300 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2586_
timestamp 18001
transform 1 0 9016 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2587_
timestamp 18001
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2588_
timestamp 18001
transform -1 0 12144 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2589_
timestamp 18001
transform -1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2590_
timestamp 18001
transform -1 0 12788 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _2591_
timestamp 18001
transform -1 0 27508 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _2592_
timestamp 18001
transform 1 0 10580 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2593_
timestamp 18001
transform -1 0 11040 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2594_
timestamp 18001
transform -1 0 10764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2595_
timestamp 18001
transform 1 0 9108 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _2596_
timestamp 18001
transform 1 0 9936 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _2597_
timestamp 18001
transform 1 0 17756 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2598_
timestamp 18001
transform -1 0 15548 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2599_
timestamp 18001
transform -1 0 13156 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2600_
timestamp 18001
transform -1 0 13340 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2601_
timestamp 18001
transform -1 0 12696 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _2602_
timestamp 18001
transform -1 0 10580 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2603_
timestamp 18001
transform -1 0 2208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2604_
timestamp 18001
transform 1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2605_
timestamp 18001
transform 1 0 9200 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2606_
timestamp 18001
transform 1 0 8004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2607_
timestamp 18001
transform 1 0 7728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2608_
timestamp 18001
transform -1 0 9200 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2609_
timestamp 18001
transform -1 0 9936 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2610_
timestamp 18001
transform 1 0 2208 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2611_
timestamp 18001
transform -1 0 11316 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2612_
timestamp 18001
transform 1 0 8924 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2613_
timestamp 18001
transform -1 0 10396 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2614_
timestamp 18001
transform 1 0 2300 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2615_
timestamp 18001
transform 1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2616_
timestamp 18001
transform 1 0 2392 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2617_
timestamp 18001
transform 1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2618_
timestamp 18001
transform -1 0 6256 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2619_
timestamp 18001
transform -1 0 7176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2620_
timestamp 18001
transform 1 0 6256 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2621_
timestamp 18001
transform -1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2622_
timestamp 18001
transform 1 0 1748 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2623_
timestamp 18001
transform -1 0 3220 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2624_
timestamp 18001
transform 1 0 3036 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2625_
timestamp 18001
transform 1 0 3680 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _2626_
timestamp 18001
transform 1 0 3220 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2627_
timestamp 18001
transform -1 0 5244 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2628_
timestamp 18001
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2629_
timestamp 18001
transform 1 0 5060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2630_
timestamp 18001
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2631_
timestamp 18001
transform -1 0 4232 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _2632_
timestamp 18001
transform 1 0 5336 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2633_
timestamp 18001
transform -1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2634_
timestamp 18001
transform 1 0 3772 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2635_
timestamp 18001
transform 1 0 1840 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2636_
timestamp 18001
transform 1 0 3220 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2637_
timestamp 18001
transform 1 0 2392 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2638_
timestamp 18001
transform -1 0 6256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2639_
timestamp 18001
transform 1 0 5428 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _2640_
timestamp 18001
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2641_
timestamp 18001
transform 1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _2642_
timestamp 18001
transform 1 0 4784 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2643_
timestamp 18001
transform -1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2644_
timestamp 18001
transform 1 0 4600 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2645_
timestamp 18001
transform -1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2646_
timestamp 18001
transform -1 0 4600 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2647_
timestamp 18001
transform 1 0 4048 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2648_
timestamp 18001
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2649_
timestamp 18001
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2650_
timestamp 18001
transform -1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2651_
timestamp 18001
transform -1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2652_
timestamp 18001
transform 1 0 6164 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2653_
timestamp 18001
transform 1 0 5244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2654_
timestamp 18001
transform -1 0 6256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _2655_
timestamp 18001
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2656_
timestamp 18001
transform -1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2657_
timestamp 18001
transform 1 0 4508 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _2658_
timestamp 18001
transform 1 0 5152 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2659_
timestamp 18001
transform -1 0 5244 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2660_
timestamp 18001
transform -1 0 10580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2661_
timestamp 18001
transform -1 0 9568 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2662_
timestamp 18001
transform 1 0 8188 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2663_
timestamp 18001
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2664_
timestamp 18001
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2665_
timestamp 18001
transform 1 0 8740 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2666_
timestamp 18001
transform -1 0 9108 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _2667_
timestamp 18001
transform -1 0 5888 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2668_
timestamp 18001
transform 1 0 6624 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2669_
timestamp 18001
transform 1 0 25300 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_4  _2670_
timestamp 18001
transform 1 0 21988 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2671_
timestamp 18001
transform 1 0 8556 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2672_
timestamp 18001
transform 1 0 10580 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2673_
timestamp 18001
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2674_
timestamp 18001
transform 1 0 3220 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2675_
timestamp 18001
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2676_
timestamp 18001
transform 1 0 6072 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2677_
timestamp 18001
transform 1 0 4508 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2678_
timestamp 18001
transform 1 0 7176 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2679_
timestamp 18001
transform -1 0 13248 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2680_
timestamp 18001
transform 1 0 12420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _2681_
timestamp 18001
transform -1 0 25116 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2682_
timestamp 18001
transform -1 0 25484 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _2683_
timestamp 18001
transform 1 0 18216 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2684_
timestamp 18001
transform 1 0 12420 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _2685_
timestamp 18001
transform 1 0 25484 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 18001
transform 1 0 27416 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 18001
transform -1 0 31372 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 18001
transform -1 0 23644 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 18001
transform 1 0 32108 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 18001
transform -1 0 25024 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2691_
timestamp 18001
transform -1 0 26128 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2692_
timestamp 18001
transform -1 0 26680 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 18001
transform 1 0 26312 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 18001
transform 1 0 24472 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 18001
transform -1 0 29992 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 18001
transform 1 0 22080 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2697_
timestamp 18001
transform -1 0 31740 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _2698_
timestamp 18001
transform 1 0 23736 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2699_
timestamp 18001
transform 1 0 21252 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2700_
timestamp 18001
transform 1 0 22264 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 18001
transform 1 0 23368 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 18001
transform -1 0 26220 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2703_
timestamp 18001
transform 1 0 22172 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2704_
timestamp 18001
transform 1 0 22172 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2705_
timestamp 18001
transform -1 0 15088 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2706_
timestamp 18001
transform -1 0 36156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2707_
timestamp 18001
transform -1 0 36156 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2708_
timestamp 18001
transform 1 0 33488 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2709_
timestamp 18001
transform 1 0 34224 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2710_
timestamp 18001
transform 1 0 34040 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2711_
timestamp 18001
transform 1 0 32016 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2712_
timestamp 18001
transform 1 0 11132 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2713_
timestamp 18001
transform 1 0 9568 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2714_
timestamp 18001
transform 1 0 12328 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2715_
timestamp 18001
transform 1 0 9568 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2716_
timestamp 18001
transform 1 0 9476 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2717_
timestamp 18001
transform 1 0 14168 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2718_
timestamp 18001
transform 1 0 19780 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2719_
timestamp 18001
transform -1 0 15916 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2720_
timestamp 18001
transform 1 0 11776 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2721_
timestamp 18001
transform -1 0 18952 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2722_
timestamp 18001
transform -1 0 17664 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2723_
timestamp 18001
transform 1 0 17204 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2724_
timestamp 18001
transform 1 0 14444 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2725_
timestamp 18001
transform 1 0 16652 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2726_
timestamp 18001
transform -1 0 14076 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2727_
timestamp 18001
transform 1 0 13800 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2728_
timestamp 18001
transform 1 0 11408 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2729_
timestamp 18001
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2730_
timestamp 18001
transform 1 0 8924 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2731_
timestamp 18001
transform -1 0 11224 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2732_
timestamp 18001
transform -1 0 11316 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2733_
timestamp 18001
transform -1 0 9936 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2734_
timestamp 18001
transform -1 0 10764 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2735_
timestamp 18001
transform 1 0 11500 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2736_
timestamp 18001
transform 1 0 10120 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2737_
timestamp 18001
transform -1 0 11408 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2738_
timestamp 18001
transform 1 0 12604 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2739_
timestamp 18001
transform 1 0 14076 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2740_
timestamp 18001
transform -1 0 16836 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2741_
timestamp 18001
transform -1 0 18768 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2742_
timestamp 18001
transform 1 0 18400 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2743_
timestamp 18001
transform 1 0 19228 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2744_
timestamp 18001
transform 1 0 8372 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2745_
timestamp 18001
transform 1 0 8924 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2746_
timestamp 18001
transform 1 0 1380 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2747_
timestamp 18001
transform 1 0 1564 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2748_
timestamp 18001
transform -1 0 4416 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2749_
timestamp 18001
transform 1 0 6348 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2750_
timestamp 18001
transform 1 0 1380 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2751_
timestamp 18001
transform 1 0 6624 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2752_
timestamp 18001
transform 1 0 8924 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2753_
timestamp 18001
transform 1 0 9660 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2754_
timestamp 18001
transform 1 0 1380 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2755_
timestamp 18001
transform 1 0 1380 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2756_
timestamp 18001
transform 1 0 1380 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2757_
timestamp 18001
transform 1 0 5336 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2758_
timestamp 18001
transform 1 0 1380 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2759_
timestamp 18001
transform 1 0 6348 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2760_
timestamp 18001
transform 1 0 18676 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2761_
timestamp 18001
transform 1 0 19596 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2762_
timestamp 18001
transform 1 0 20976 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2763_
timestamp 18001
transform -1 0 23920 0 1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2764_
timestamp 18001
transform 1 0 22540 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2765_
timestamp 18001
transform -1 0 23920 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2766_
timestamp 18001
transform 1 0 19872 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2767_
timestamp 18001
transform 1 0 19320 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2768_
timestamp 18001
transform 1 0 22356 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2769_
timestamp 18001
transform -1 0 14996 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2770_
timestamp 18001
transform -1 0 13432 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2771_
timestamp 18001
transform 1 0 8740 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2772_
timestamp 18001
transform 1 0 3680 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2773_
timestamp 18001
transform 1 0 3772 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2774_
timestamp 18001
transform 1 0 4692 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2775_
timestamp 18001
transform 1 0 6348 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2776_
timestamp 18001
transform 1 0 7820 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2777_
timestamp 18001
transform 1 0 7268 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2778_
timestamp 18001
transform 1 0 9016 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2779_
timestamp 18001
transform 1 0 1380 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2780_
timestamp 18001
transform 1 0 1380 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2781_
timestamp 18001
transform 1 0 2576 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2782_
timestamp 18001
transform 1 0 3680 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2783_
timestamp 18001
transform 1 0 1380 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2784_
timestamp 18001
transform 1 0 2208 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2785_
timestamp 18001
transform -1 0 3680 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2786_
timestamp 18001
transform -1 0 3864 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2787_
timestamp 18001
transform -1 0 3496 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2788_
timestamp 18001
transform -1 0 3680 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2789_
timestamp 18001
transform -1 0 3588 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2790_
timestamp 18001
transform -1 0 4508 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2791_
timestamp 18001
transform 1 0 1472 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2792_
timestamp 18001
transform -1 0 3588 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2793_
timestamp 18001
transform 1 0 9568 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2794_
timestamp 18001
transform 1 0 9016 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2795_
timestamp 18001
transform 1 0 1380 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2796_
timestamp 18001
transform 1 0 1380 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2797_
timestamp 18001
transform 1 0 1380 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2798_
timestamp 18001
transform -1 0 4048 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2799_
timestamp 18001
transform 1 0 2484 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2800_
timestamp 18001
transform 1 0 6992 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2801_
timestamp 18001
transform 1 0 21804 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2802_
timestamp 18001
transform -1 0 25484 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2803_
timestamp 18001
transform 1 0 7820 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2804_
timestamp 18001
transform 1 0 9568 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2805_
timestamp 18001
transform 1 0 1840 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2806_
timestamp 18001
transform 1 0 1840 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2807_
timestamp 18001
transform 1 0 1932 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2808_
timestamp 18001
transform 1 0 5336 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2809_
timestamp 18001
transform 1 0 3772 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2810_
timestamp 18001
transform 1 0 6440 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2811_
timestamp 18001
transform 1 0 11868 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2812_
timestamp 18001
transform 1 0 24380 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2813_
timestamp 18001
transform 1 0 11776 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _2814_
timestamp 18001
transform -1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 18001
transform -1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 18001
transform -1 0 35236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 18001
transform 1 0 16836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform 1 0 19228 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 18001
transform 1 0 7636 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 18001
transform 1 0 7728 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 18001
transform -1 0 14352 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 18001
transform -1 0 11040 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 18001
transform -1 0 4416 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 18001
transform 1 0 3772 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 18001
transform 1 0 7452 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 18001
transform 1 0 7360 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 18001
transform -1 0 23552 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 18001
transform 1 0 22080 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 18001
transform 1 0 28152 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 18001
transform 1 0 27968 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 18001
transform -1 0 20240 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 18001
transform -1 0 19136 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 18001
transform -1 0 25944 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 18001
transform -1 0 24104 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_8  clkload0
timestamp 18001
transform 1 0 7636 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload1
timestamp 18001
transform 1 0 7728 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  clkload2
timestamp 18001
transform 1 0 15088 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_6  clkload3
timestamp 18001
transform 1 0 11500 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  clkload4
timestamp 18001
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  clkload5
timestamp 18001
transform -1 0 8096 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload6
timestamp 18001
transform 1 0 8096 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  clkload7
timestamp 18001
transform 1 0 22540 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload8
timestamp 18001
transform -1 0 22908 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload9
timestamp 18001
transform 1 0 28152 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  clkload10
timestamp 18001
transform 1 0 27968 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_6  clkload11
timestamp 18001
transform 1 0 20240 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload12
timestamp 18001
transform -1 0 19136 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload13
timestamp 18001
transform 1 0 24840 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload14
timestamp 18001
transform 1 0 22264 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 18001
transform 1 0 15364 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 18001
transform -1 0 10764 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 18001
transform 1 0 32660 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 18001
transform 1 0 7544 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 18001
transform -1 0 11316 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 18001
transform -1 0 11960 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 18001
transform -1 0 17296 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 18001
transform -1 0 17020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 18001
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 18001
transform 1 0 25024 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout29
timestamp 18001
transform -1 0 5244 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 18001
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 18001
transform -1 0 10764 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout32
timestamp 18001
transform 1 0 10304 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 18001
transform -1 0 28336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 18001
transform 1 0 31372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout35
timestamp 18001
transform -1 0 33120 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 18001
transform 1 0 29532 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout37
timestamp 18001
transform 1 0 27508 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 18001
transform -1 0 26772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 18001
transform -1 0 24288 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 18001
transform -1 0 30452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 18001
transform -1 0 24288 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 18001
transform -1 0 24288 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 18001
transform 1 0 11500 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 18001
transform -1 0 12512 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 18001
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 18001
transform -1 0 14720 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 18001
transform 1 0 21804 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 18001
transform -1 0 17204 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 18001
transform -1 0 16744 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 18001
transform -1 0 16836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout51
timestamp 18001
transform 1 0 19228 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 18001
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp 18001
transform 1 0 19596 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 18001
transform 1 0 14260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 18001
transform -1 0 20424 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout56
timestamp 18001
transform 1 0 20424 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp 18001
transform -1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 18001
transform 1 0 25760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout59
timestamp 18001
transform 1 0 28520 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 18001
transform 1 0 32844 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout61
timestamp 18001
transform -1 0 17572 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 18001
transform 1 0 26128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout63
timestamp 18001
transform -1 0 15364 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout64
timestamp 18001
transform 1 0 21528 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout65
timestamp 18001
transform -1 0 26588 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout66
timestamp 18001
transform 1 0 26312 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 18001
transform 1 0 24472 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 18001
transform -1 0 25392 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 18001
transform -1 0 26496 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 18001
transform -1 0 19136 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout71
timestamp 18001
transform -1 0 21712 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 18001
transform 1 0 30452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout73
timestamp 18001
transform 1 0 32292 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout74
timestamp 18001
transform -1 0 29348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout75
timestamp 18001
transform 1 0 32844 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 18001
transform -1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout77
timestamp 18001
transform 1 0 31372 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp 18001
transform -1 0 26312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout79
timestamp 18001
transform 1 0 34684 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 18001
transform 1 0 31280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 18001
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout82
timestamp 18001
transform -1 0 32844 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 18001
transform -1 0 26404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout84
timestamp 18001
transform -1 0 35972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout85
timestamp 18001
transform -1 0 24748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout86
timestamp 18001
transform -1 0 23368 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout87
timestamp 18001
transform 1 0 29808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout88
timestamp 18001
transform -1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout89
timestamp 18001
transform -1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout90
timestamp 18001
transform -1 0 30176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp 18001
transform 1 0 33028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout92
timestamp 18001
transform -1 0 35604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 18001
transform -1 0 30452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout94
timestamp 18001
transform -1 0 30452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout95
timestamp 18001
transform -1 0 33764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout96
timestamp 18001
transform 1 0 34684 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout97
timestamp 18001
transform -1 0 28428 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  fanout98
timestamp 18001
transform 1 0 28980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 18001
transform 1 0 35236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout100
timestamp 18001
transform 1 0 35052 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout101
timestamp 18001
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout102
timestamp 18001
transform 1 0 34868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout103
timestamp 18001
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout104
timestamp 18001
transform 1 0 24380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout105
timestamp 18001
transform 1 0 22908 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp 18001
transform -1 0 19872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout107
timestamp 18001
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 18001
transform -1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout109
timestamp 18001
transform 1 0 23736 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout110
timestamp 18001
transform 1 0 23276 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp 18001
transform -1 0 21988 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout112
timestamp 18001
transform -1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout113
timestamp 18001
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout114
timestamp 18001
transform -1 0 23092 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 18001
transform 1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout116
timestamp 18001
transform -1 0 18492 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout117
timestamp 18001
transform -1 0 26220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 18001
transform 1 0 17572 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout119
timestamp 18001
transform -1 0 21620 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout120
timestamp 18001
transform -1 0 19136 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout121
timestamp 18001
transform 1 0 21988 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout122
timestamp 18001
transform 1 0 24932 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout123
timestamp 18001
transform 1 0 26588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout124
timestamp 18001
transform -1 0 26588 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout125
timestamp 18001
transform 1 0 26496 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout126
timestamp 18001
transform 1 0 29532 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout127
timestamp 18001
transform -1 0 11316 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout128
timestamp 18001
transform 1 0 19780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout129
timestamp 18001
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout130
timestamp 18001
transform 1 0 9568 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout131
timestamp 18001
transform -1 0 9936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout132
timestamp 18001
transform -1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout133
timestamp 18001
transform 1 0 35604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout134
timestamp 18001
transform -1 0 10212 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout135
timestamp 18001
transform -1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout136
timestamp 18001
transform 1 0 17020 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout137
timestamp 18001
transform -1 0 11132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout138
timestamp 18001
transform -1 0 15548 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout139
timestamp 18001
transform -1 0 22540 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout140
timestamp 18001
transform -1 0 29624 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout141
timestamp 18001
transform -1 0 25760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout142
timestamp 18001
transform -1 0 32844 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout143
timestamp 18001
transform 1 0 35696 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout144
timestamp 18001
transform -1 0 36156 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout145
timestamp 18001
transform -1 0 31740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout146
timestamp 18001
transform -1 0 28612 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout147
timestamp 18001
transform -1 0 29256 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69
timestamp 18001
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 18001
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_189
timestamp 18001
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 18001
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636986456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_209
timestamp 18001
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_217
timestamp 18001
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 18001
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 18001
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_259
timestamp 1636986456
transform 1 0 24932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_271
timestamp 18001
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 18001
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636986456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636986456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 18001
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636986456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636986456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 18001
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1636986456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1636986456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 18001
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1636986456
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_377
timestamp 18001
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_69
timestamp 18001
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 18001
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_213
timestamp 18001
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_217
timestamp 18001
transform 1 0 21068 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_265
timestamp 1636986456
transform 1 0 25484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 18001
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636986456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636986456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636986456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 18001
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_373
timestamp 18001
transform 1 0 35420 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_65
timestamp 18001
transform 1 0 7084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 18001
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_110
timestamp 18001
transform 1 0 11224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_197
timestamp 18001
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 18001
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_273
timestamp 18001
transform 1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_291
timestamp 1636986456
transform 1 0 27876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_303
timestamp 18001
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 18001
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636986456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636986456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1636986456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1636986456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 18001
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 18001
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_377
timestamp 18001
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636986456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636986456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 18001
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 18001
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 18001
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_136
timestamp 18001
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 18001
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_198
timestamp 1636986456
transform 1 0 19320 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_210
timestamp 18001
transform 1 0 20424 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_216
timestamp 18001
transform 1 0 20976 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_225
timestamp 18001
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_257
timestamp 18001
transform 1 0 24748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_270
timestamp 18001
transform 1 0 25944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_278
timestamp 18001
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636986456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_293
timestamp 18001
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_304
timestamp 1636986456
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_316
timestamp 1636986456
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_328
timestamp 18001
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_373
timestamp 18001
transform 1 0 35420 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_65
timestamp 18001
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_73
timestamp 18001
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_126
timestamp 18001
transform 1 0 12696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_170
timestamp 18001
transform 1 0 16744 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_190
timestamp 18001
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636986456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_209
timestamp 18001
transform 1 0 20332 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_217
timestamp 18001
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_243
timestamp 18001
transform 1 0 23460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 18001
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636986456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1636986456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1636986456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1636986456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 18001
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 18001
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1636986456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 18001
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1636986456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_377
timestamp 18001
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_69
timestamp 18001
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_75
timestamp 18001
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_96
timestamp 18001
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_157
timestamp 18001
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 18001
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1636986456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1636986456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_193
timestamp 18001
transform 1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1636986456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 18001
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 18001
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 18001
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_239
timestamp 1636986456
transform 1 0 23092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_251
timestamp 1636986456
transform 1 0 24196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_263
timestamp 1636986456
transform 1 0 25300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_275
timestamp 18001
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_286
timestamp 1636986456
transform 1 0 27416 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_298
timestamp 1636986456
transform 1 0 28520 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_310
timestamp 18001
transform 1 0 29624 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_319
timestamp 1636986456
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_331
timestamp 18001
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 18001
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1636986456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1636986456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_373
timestamp 18001
transform 1 0 35420 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_41
timestamp 18001
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_47
timestamp 1636986456
transform 1 0 5428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_59
timestamp 18001
transform 1 0 6532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_67
timestamp 18001
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_73
timestamp 18001
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 18001
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_95
timestamp 18001
transform 1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_115
timestamp 18001
transform 1 0 11684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_149
timestamp 18001
transform 1 0 14812 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_158
timestamp 18001
transform 1 0 15640 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_168
timestamp 18001
transform 1 0 16560 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_181
timestamp 1636986456
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_193
timestamp 18001
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_197
timestamp 18001
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_207
timestamp 18001
transform 1 0 20148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_211
timestamp 18001
transform 1 0 20516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_226
timestamp 18001
transform 1 0 21896 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_234
timestamp 18001
transform 1 0 22632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_253
timestamp 18001
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_261
timestamp 1636986456
transform 1 0 25116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_273
timestamp 18001
transform 1 0 26220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_285
timestamp 18001
transform 1 0 27324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_302
timestamp 18001
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_309
timestamp 18001
transform 1 0 29532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_336
timestamp 18001
transform 1 0 32016 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_348
timestamp 1636986456
transform 1 0 33120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_360
timestamp 18001
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1636986456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_377
timestamp 18001
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_27
timestamp 18001
transform 1 0 3588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_48
timestamp 18001
transform 1 0 5520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 18001
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_60
timestamp 18001
transform 1 0 6624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_84
timestamp 18001
transform 1 0 8832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_139
timestamp 18001
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_148
timestamp 18001
transform 1 0 14720 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_152
timestamp 18001
transform 1 0 15088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_158
timestamp 18001
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 18001
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1636986456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_186
timestamp 18001
transform 1 0 18216 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_195
timestamp 1636986456
transform 1 0 19044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_207
timestamp 18001
transform 1 0 20148 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_215
timestamp 18001
transform 1 0 20884 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_221
timestamp 18001
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1636986456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_237
timestamp 18001
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_243
timestamp 18001
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_253
timestamp 18001
transform 1 0 24380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_276
timestamp 18001
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_281
timestamp 18001
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_328
timestamp 18001
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_360
timestamp 1636986456
transform 1 0 34224 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_372
timestamp 18001
transform 1 0 35328 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_380
timestamp 18001
transform 1 0 36064 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 18001
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_58
timestamp 18001
transform 1 0 6440 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_120
timestamp 18001
transform 1 0 12144 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_134
timestamp 18001
transform 1 0 13432 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_147
timestamp 1636986456
transform 1 0 14628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_159
timestamp 1636986456
transform 1 0 15732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_171
timestamp 18001
transform 1 0 16836 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_179
timestamp 18001
transform 1 0 17572 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 18001
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_210
timestamp 1636986456
transform 1 0 20424 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_222
timestamp 1636986456
transform 1 0 21528 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_234
timestamp 1636986456
transform 1 0 22632 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_246
timestamp 18001
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1636986456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1636986456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_277
timestamp 18001
transform 1 0 26588 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_290
timestamp 1636986456
transform 1 0 27784 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_302
timestamp 18001
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_309
timestamp 18001
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_315
timestamp 1636986456
transform 1 0 30084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_327
timestamp 1636986456
transform 1 0 31188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_351
timestamp 1636986456
transform 1 0 33396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 18001
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1636986456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_377
timestamp 18001
transform 1 0 35788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 18001
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_11
timestamp 18001
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_41
timestamp 18001
transform 1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_69
timestamp 18001
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_92
timestamp 18001
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 18001
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 18001
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_149
timestamp 18001
transform 1 0 14812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_155
timestamp 18001
transform 1 0 15364 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_160
timestamp 18001
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_175
timestamp 18001
transform 1 0 17204 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_183
timestamp 18001
transform 1 0 17940 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_194
timestamp 18001
transform 1 0 18952 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_211
timestamp 18001
transform 1 0 20516 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_219
timestamp 18001
transform 1 0 21252 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_241
timestamp 1636986456
transform 1 0 23276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_253
timestamp 18001
transform 1 0 24380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_269
timestamp 18001
transform 1 0 25852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_277
timestamp 18001
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_281
timestamp 18001
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_292
timestamp 1636986456
transform 1 0 27968 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_304
timestamp 1636986456
transform 1 0 29072 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_316
timestamp 18001
transform 1 0 30176 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 18001
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_337
timestamp 18001
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_348
timestamp 1636986456
transform 1 0 33120 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_360
timestamp 1636986456
transform 1 0 34224 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_372
timestamp 18001
transform 1 0 35328 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_380
timestamp 18001
transform 1 0 36064 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 18001
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_41
timestamp 18001
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_45
timestamp 18001
transform 1 0 5244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_54
timestamp 18001
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 18001
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_94
timestamp 18001
transform 1 0 9752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_103
timestamp 18001
transform 1 0 10580 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 18001
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_155
timestamp 18001
transform 1 0 15364 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_162
timestamp 1636986456
transform 1 0 16008 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_174
timestamp 1636986456
transform 1 0 17112 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_186
timestamp 18001
transform 1 0 18216 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 18001
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1636986456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_209
timestamp 18001
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_218
timestamp 1636986456
transform 1 0 21160 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_230
timestamp 18001
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_234
timestamp 18001
transform 1 0 22632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_244
timestamp 18001
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_260
timestamp 18001
transform 1 0 25024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_272
timestamp 18001
transform 1 0 26128 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_295
timestamp 18001
transform 1 0 28244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_302
timestamp 18001
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_327
timestamp 1636986456
transform 1 0 31188 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_339
timestamp 1636986456
transform 1 0 32292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_351
timestamp 1636986456
transform 1 0 33396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 18001
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_376
timestamp 18001
transform 1 0 35696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_380
timestamp 18001
transform 1 0 36064 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_35
timestamp 18001
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_90
timestamp 18001
transform 1 0 9384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_106
timestamp 18001
transform 1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_127
timestamp 1636986456
transform 1 0 12788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_139
timestamp 1636986456
transform 1 0 13892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_151
timestamp 18001
transform 1 0 14996 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_159
timestamp 18001
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_176
timestamp 18001
transform 1 0 17296 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_184
timestamp 18001
transform 1 0 18032 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1636986456
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_205
timestamp 18001
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_213
timestamp 18001
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_221
timestamp 18001
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1636986456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_237
timestamp 18001
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_246
timestamp 1636986456
transform 1 0 23736 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_258
timestamp 18001
transform 1 0 24840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_262
timestamp 18001
transform 1 0 25208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 18001
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 18001
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1636986456
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1636986456
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_305
timestamp 18001
transform 1 0 29164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_327
timestamp 18001
transform 1 0 31188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 18001
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_337
timestamp 18001
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_343
timestamp 18001
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_360
timestamp 18001
transform 1 0 34224 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_15
timestamp 18001
transform 1 0 2484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_23
timestamp 18001
transform 1 0 3220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_51
timestamp 18001
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_116
timestamp 18001
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_120
timestamp 18001
transform 1 0 12144 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_130
timestamp 18001
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 18001
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1636986456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1636986456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_165
timestamp 18001
transform 1 0 16284 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_186
timestamp 18001
transform 1 0 18216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 18001
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_197
timestamp 18001
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_205
timestamp 18001
transform 1 0 19964 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_214
timestamp 1636986456
transform 1 0 20792 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_226
timestamp 1636986456
transform 1 0 21896 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_238
timestamp 18001
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_247
timestamp 18001
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 18001
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636986456
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1636986456
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_277
timestamp 18001
transform 1 0 26588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_287
timestamp 18001
transform 1 0 27508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_295
timestamp 18001
transform 1 0 28244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_301
timestamp 18001
transform 1 0 28796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_309
timestamp 18001
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_318
timestamp 18001
transform 1 0 30360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_348
timestamp 18001
transform 1 0 33120 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_354
timestamp 18001
transform 1 0 33672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_362
timestamp 18001
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_365
timestamp 18001
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_375
timestamp 18001
transform 1 0 35604 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 18001
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_11
timestamp 18001
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_23
timestamp 18001
transform 1 0 3220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_34
timestamp 18001
transform 1 0 4232 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_60
timestamp 18001
transform 1 0 6624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_69
timestamp 18001
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_76
timestamp 18001
transform 1 0 8096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_92
timestamp 18001
transform 1 0 9568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 18001
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_119
timestamp 18001
transform 1 0 12052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_134
timestamp 18001
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_142
timestamp 18001
transform 1 0 14168 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_154
timestamp 1636986456
transform 1 0 15272 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 18001
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_175
timestamp 1636986456
transform 1 0 17204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_187
timestamp 18001
transform 1 0 18308 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_195
timestamp 18001
transform 1 0 19044 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_201
timestamp 18001
transform 1 0 19596 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_209
timestamp 18001
transform 1 0 20332 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_219
timestamp 18001
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 18001
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_238
timestamp 1636986456
transform 1 0 23000 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_250
timestamp 1636986456
transform 1 0 24104 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_262
timestamp 18001
transform 1 0 25208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 18001
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_285
timestamp 1636986456
transform 1 0 27324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_297
timestamp 1636986456
transform 1 0 28428 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_309
timestamp 18001
transform 1 0 29532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_316
timestamp 18001
transform 1 0 30176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_322
timestamp 18001
transform 1 0 30728 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_334
timestamp 18001
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_342
timestamp 18001
transform 1 0 32568 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_348
timestamp 18001
transform 1 0 33120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_3
timestamp 18001
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_19
timestamp 18001
transform 1 0 2852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 18001
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_44
timestamp 18001
transform 1 0 5152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_66
timestamp 18001
transform 1 0 7176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_71
timestamp 18001
transform 1 0 7636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_75
timestamp 18001
transform 1 0 8004 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 18001
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_111
timestamp 18001
transform 1 0 11316 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_120
timestamp 18001
transform 1 0 12144 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_127
timestamp 1636986456
transform 1 0 12788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 18001
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_141
timestamp 18001
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_147
timestamp 18001
transform 1 0 14628 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_155
timestamp 1636986456
transform 1 0 15364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_167
timestamp 18001
transform 1 0 16468 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_175
timestamp 18001
transform 1 0 17204 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_183
timestamp 18001
transform 1 0 17940 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 18001
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 18001
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1636986456
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_209
timestamp 18001
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_213
timestamp 18001
transform 1 0 20700 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_219
timestamp 1636986456
transform 1 0 21252 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_231
timestamp 18001
transform 1 0 22356 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_243
timestamp 18001
transform 1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 18001
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp 18001
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_275
timestamp 18001
transform 1 0 26404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_306
timestamp 18001
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_328
timestamp 18001
transform 1 0 31280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_345
timestamp 18001
transform 1 0 32844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 18001
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 18001
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1636986456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_69
timestamp 18001
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_73
timestamp 18001
transform 1 0 7820 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 18001
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 18001
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1636986456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1636986456
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1636986456
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_149
timestamp 18001
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_157
timestamp 18001
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 18001
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_169
timestamp 18001
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_175
timestamp 18001
transform 1 0 17204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_205
timestamp 18001
transform 1 0 19964 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_225
timestamp 18001
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_233
timestamp 18001
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_242
timestamp 18001
transform 1 0 23368 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_254
timestamp 18001
transform 1 0 24472 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_260
timestamp 18001
transform 1 0 25024 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_268
timestamp 1636986456
transform 1 0 25760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_281
timestamp 18001
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_289
timestamp 18001
transform 1 0 27692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_293
timestamp 18001
transform 1 0 28060 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_319
timestamp 1636986456
transform 1 0 30452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_331
timestamp 18001
transform 1 0 31556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 18001
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_351
timestamp 18001
transform 1 0 33396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_359
timestamp 18001
transform 1 0 34132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_380
timestamp 18001
transform 1 0 36064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 18001
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 18001
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_101
timestamp 18001
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_108
timestamp 18001
transform 1 0 11040 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 18001
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 18001
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_141
timestamp 18001
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_151
timestamp 1636986456
transform 1 0 14996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_163
timestamp 18001
transform 1 0 16100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_169
timestamp 18001
transform 1 0 16652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_179
timestamp 18001
transform 1 0 17572 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 18001
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 18001
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_202
timestamp 1636986456
transform 1 0 19688 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_214
timestamp 1636986456
transform 1 0 20792 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_226
timestamp 18001
transform 1 0 21896 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_246
timestamp 18001
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_257
timestamp 1636986456
transform 1 0 24748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_269
timestamp 1636986456
transform 1 0 25852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_281
timestamp 18001
transform 1 0 26956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_285
timestamp 18001
transform 1 0 27324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_289
timestamp 18001
transform 1 0 27692 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 18001
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_316
timestamp 1636986456
transform 1 0 30176 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_328
timestamp 18001
transform 1 0 31280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_334
timestamp 18001
transform 1 0 31832 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_350
timestamp 1636986456
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_362
timestamp 18001
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_379
timestamp 18001
transform 1 0 35972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 18001
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_11
timestamp 18001
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_22
timestamp 1636986456
transform 1 0 3128 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_34
timestamp 18001
transform 1 0 4232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 18001
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_105
timestamp 18001
transform 1 0 10764 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_133
timestamp 1636986456
transform 1 0 13340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_145
timestamp 18001
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_158
timestamp 18001
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 18001
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_184
timestamp 1636986456
transform 1 0 18032 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_196
timestamp 1636986456
transform 1 0 19136 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_208
timestamp 18001
transform 1 0 20240 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 18001
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 18001
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1636986456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_237
timestamp 18001
transform 1 0 22908 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_242
timestamp 1636986456
transform 1 0 23368 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_254
timestamp 1636986456
transform 1 0 24472 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_266
timestamp 18001
transform 1 0 25576 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_274
timestamp 18001
transform 1 0 26312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_290
timestamp 18001
transform 1 0 27784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_297
timestamp 18001
transform 1 0 28428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_307
timestamp 18001
transform 1 0 29348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_323
timestamp 18001
transform 1 0 30820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_327
timestamp 18001
transform 1 0 31188 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_337
timestamp 18001
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_351
timestamp 18001
transform 1 0 33396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_359
timestamp 18001
transform 1 0 34132 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 18001
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 18001
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_23
timestamp 18001
transform 1 0 3220 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_40
timestamp 18001
transform 1 0 4784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_48
timestamp 18001
transform 1 0 5520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_64
timestamp 18001
transform 1 0 6992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 18001
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_108
timestamp 18001
transform 1 0 11040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_117
timestamp 18001
transform 1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_125
timestamp 18001
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_131
timestamp 18001
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 18001
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_148
timestamp 18001
transform 1 0 14720 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_157
timestamp 1636986456
transform 1 0 15548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_169
timestamp 18001
transform 1 0 16652 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_175
timestamp 18001
transform 1 0 17204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 18001
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1636986456
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_209
timestamp 18001
transform 1 0 20332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_217
timestamp 18001
transform 1 0 21068 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_224
timestamp 18001
transform 1 0 21712 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_232
timestamp 18001
transform 1 0 22448 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_242
timestamp 18001
transform 1 0 23368 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 18001
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_269
timestamp 18001
transform 1 0 25852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_277
timestamp 18001
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_298
timestamp 18001
transform 1 0 28520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_306
timestamp 18001
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_317
timestamp 18001
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_328
timestamp 1636986456
transform 1 0 31280 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_346
timestamp 18001
transform 1 0 32936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_354
timestamp 18001
transform 1 0 33672 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_373
timestamp 18001
transform 1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_32
timestamp 18001
transform 1 0 4048 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 18001
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 18001
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 18001
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1636986456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1636986456
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_137
timestamp 18001
transform 1 0 13708 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_162
timestamp 18001
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1636986456
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1636986456
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_193
timestamp 18001
transform 1 0 18860 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_199
timestamp 18001
transform 1 0 19412 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1636986456
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 18001
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 18001
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_231
timestamp 18001
transform 1 0 22356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_235
timestamp 18001
transform 1 0 22724 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_241
timestamp 18001
transform 1 0 23276 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_251
timestamp 1636986456
transform 1 0 24196 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_263
timestamp 1636986456
transform 1 0 25300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_275
timestamp 18001
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 18001
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1636986456
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1636986456
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1636986456
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1636986456
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 18001
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 18001
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1636986456
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1636986456
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1636986456
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_373
timestamp 18001
transform 1 0 35420 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 18001
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_11
timestamp 18001
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_23
timestamp 18001
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 18001
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_34
timestamp 18001
transform 1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_45
timestamp 18001
transform 1 0 5244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_50
timestamp 18001
transform 1 0 5704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_60
timestamp 18001
transform 1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_71
timestamp 18001
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 18001
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 18001
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_93
timestamp 18001
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_106
timestamp 1636986456
transform 1 0 10856 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_118
timestamp 18001
transform 1 0 11960 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_130
timestamp 18001
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 18001
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 18001
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_151
timestamp 18001
transform 1 0 14996 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_159
timestamp 18001
transform 1 0 15732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_174
timestamp 18001
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_184
timestamp 1636986456
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_212
timestamp 1636986456
transform 1 0 20608 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_224
timestamp 1636986456
transform 1 0 21712 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_236
timestamp 1636986456
transform 1 0 22816 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_248
timestamp 18001
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1636986456
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_265
timestamp 18001
transform 1 0 25484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_271
timestamp 18001
transform 1 0 26036 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_278
timestamp 1636986456
transform 1 0 26680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_290
timestamp 1636986456
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_302
timestamp 18001
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_316
timestamp 18001
transform 1 0 30176 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_324
timestamp 1636986456
transform 1 0 30912 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_336
timestamp 18001
transform 1 0 32016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_340
timestamp 18001
transform 1 0 32384 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_349
timestamp 1636986456
transform 1 0 33212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_361
timestamp 18001
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1636986456
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_377
timestamp 18001
transform 1 0 35788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_45
timestamp 18001
transform 1 0 5244 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 18001
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_72
timestamp 18001
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_86
timestamp 18001
transform 1 0 9016 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_126
timestamp 1636986456
transform 1 0 12696 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_138
timestamp 18001
transform 1 0 13800 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_145
timestamp 1636986456
transform 1 0 14444 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_157
timestamp 18001
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 18001
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_176
timestamp 1636986456
transform 1 0 17296 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_188
timestamp 1636986456
transform 1 0 18400 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_200
timestamp 1636986456
transform 1 0 19504 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_212
timestamp 18001
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 18001
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 18001
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_241
timestamp 18001
transform 1 0 23276 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_255
timestamp 18001
transform 1 0 24564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_267
timestamp 18001
transform 1 0 25668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_271
timestamp 18001
transform 1 0 26036 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 18001
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_281
timestamp 18001
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_289
timestamp 18001
transform 1 0 27692 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_295
timestamp 18001
transform 1 0 28244 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_304
timestamp 1636986456
transform 1 0 29072 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_316
timestamp 18001
transform 1 0 30176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_324
timestamp 18001
transform 1 0 30912 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_333
timestamp 18001
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_337
timestamp 18001
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_346
timestamp 18001
transform 1 0 32936 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_352
timestamp 18001
transform 1 0 33488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_359
timestamp 18001
transform 1 0 34132 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_378
timestamp 18001
transform 1 0 35880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 18001
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_7
timestamp 18001
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_51
timestamp 18001
transform 1 0 5796 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_61
timestamp 18001
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_71
timestamp 18001
transform 1 0 7636 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 18001
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_114
timestamp 1636986456
transform 1 0 11592 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_126
timestamp 18001
transform 1 0 12696 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 18001
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1636986456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1636986456
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1636986456
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_177
timestamp 18001
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_185
timestamp 18001
transform 1 0 18124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 18001
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_218
timestamp 1636986456
transform 1 0 21160 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_230
timestamp 18001
transform 1 0 22264 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_247
timestamp 18001
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 18001
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_253
timestamp 18001
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_259
timestamp 18001
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_274
timestamp 18001
transform 1 0 26312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_299
timestamp 18001
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 18001
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_309
timestamp 18001
transform 1 0 29532 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_318
timestamp 1636986456
transform 1 0 30360 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_330
timestamp 1636986456
transform 1 0 31464 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_342
timestamp 1636986456
transform 1 0 32568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_354
timestamp 18001
transform 1 0 33672 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_361
timestamp 18001
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1636986456
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_377
timestamp 18001
transform 1 0 35788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_3
timestamp 18001
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 18001
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_63
timestamp 18001
transform 1 0 6900 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_72
timestamp 18001
transform 1 0 7728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 18001
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1636986456
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1636986456
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1636986456
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_159
timestamp 18001
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 18001
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1636986456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_188
timestamp 18001
transform 1 0 18400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_199
timestamp 18001
transform 1 0 19412 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_207
timestamp 18001
transform 1 0 20148 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_212
timestamp 1636986456
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1636986456
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_237
timestamp 18001
transform 1 0 22908 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_245
timestamp 18001
transform 1 0 23644 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1636986456
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 18001
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 18001
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_281
timestamp 18001
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_292
timestamp 1636986456
transform 1 0 27968 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_304
timestamp 1636986456
transform 1 0 29072 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_316
timestamp 1636986456
transform 1 0 30176 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_328
timestamp 18001
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_345
timestamp 1636986456
transform 1 0 32844 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_357
timestamp 1636986456
transform 1 0 33948 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_369
timestamp 1636986456
transform 1 0 35052 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 18001
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_7
timestamp 18001
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 18001
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_88
timestamp 18001
transform 1 0 9200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_120
timestamp 18001
transform 1 0 12144 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_129
timestamp 18001
transform 1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 18001
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_141
timestamp 18001
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_147
timestamp 18001
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_156
timestamp 18001
transform 1 0 15456 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_168
timestamp 1636986456
transform 1 0 16560 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_180
timestamp 18001
transform 1 0 17664 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_188
timestamp 18001
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_201
timestamp 18001
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_223
timestamp 1636986456
transform 1 0 21620 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_235
timestamp 18001
transform 1 0 22724 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 18001
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 18001
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1636986456
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1636986456
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1636986456
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1636986456
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 18001
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 18001
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_309
timestamp 18001
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_317
timestamp 18001
transform 1 0 30268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_335
timestamp 18001
transform 1 0 31924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_354
timestamp 18001
transform 1 0 33672 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 18001
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_371
timestamp 18001
transform 1 0 35236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_379
timestamp 18001
transform 1 0 35972 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_32
timestamp 18001
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_36
timestamp 18001
transform 1 0 4416 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 18001
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 18001
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_78
timestamp 18001
transform 1 0 8280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_90
timestamp 18001
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_122
timestamp 18001
transform 1 0 12328 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_134
timestamp 18001
transform 1 0 13432 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_154
timestamp 1636986456
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 18001
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 18001
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 18001
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1636986456
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1636986456
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1636986456
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 18001
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 18001
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_243
timestamp 18001
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_247
timestamp 18001
transform 1 0 23828 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_263
timestamp 18001
transform 1 0 25300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_272
timestamp 18001
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_281
timestamp 18001
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_289
timestamp 18001
transform 1 0 27692 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_310
timestamp 1636986456
transform 1 0 29624 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_322
timestamp 18001
transform 1 0 30728 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_333
timestamp 18001
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1636986456
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1636986456
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_361
timestamp 18001
transform 1 0 34316 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_371
timestamp 18001
transform 1 0 35236 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_379
timestamp 18001
transform 1 0 35972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_3
timestamp 18001
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_18
timestamp 18001
transform 1 0 2760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_43
timestamp 18001
transform 1 0 5060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_71
timestamp 18001
transform 1 0 7636 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 18001
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_98
timestamp 18001
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_119
timestamp 18001
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_128
timestamp 1636986456
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1636986456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1636986456
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1636986456
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1636986456
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 18001
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 18001
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1636986456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1636986456
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1636986456
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_244
timestamp 18001
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_261
timestamp 18001
transform 1 0 25116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_271
timestamp 18001
transform 1 0 26036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_288
timestamp 18001
transform 1 0 27600 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_305
timestamp 18001
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1636986456
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1636986456
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_333
timestamp 18001
transform 1 0 31740 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_359
timestamp 18001
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 18001
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_365
timestamp 18001
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_38
timestamp 18001
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 18001
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_66
timestamp 18001
transform 1 0 7176 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_87
timestamp 18001
transform 1 0 9108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_103
timestamp 18001
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 18001
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 18001
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_127
timestamp 1636986456
transform 1 0 12788 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_139
timestamp 1636986456
transform 1 0 13892 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_151
timestamp 18001
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_156
timestamp 18001
transform 1 0 15456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 18001
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 18001
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_177
timestamp 18001
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_183
timestamp 1636986456
transform 1 0 17940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_195
timestamp 18001
transform 1 0 19044 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_211
timestamp 1636986456
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 18001
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_246
timestamp 1636986456
transform 1 0 23736 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_258
timestamp 18001
transform 1 0 24840 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_266
timestamp 1636986456
transform 1 0 25576 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 18001
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_281
timestamp 18001
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_303
timestamp 1636986456
transform 1 0 28980 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_315
timestamp 18001
transform 1 0 30084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_323
timestamp 18001
transform 1 0 30820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_327
timestamp 18001
transform 1 0 31188 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_342
timestamp 1636986456
transform 1 0 32568 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_354
timestamp 1636986456
transform 1 0 33672 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_366
timestamp 1636986456
transform 1 0 34776 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_378
timestamp 18001
transform 1 0 35880 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636986456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_15
timestamp 18001
transform 1 0 2484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_23
timestamp 18001
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 18001
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_45
timestamp 18001
transform 1 0 5244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 18001
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_96
timestamp 18001
transform 1 0 9936 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_103
timestamp 18001
transform 1 0 10580 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_128
timestamp 1636986456
transform 1 0 12880 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_150
timestamp 18001
transform 1 0 14904 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_163
timestamp 1636986456
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 18001
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_197
timestamp 18001
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_205
timestamp 18001
transform 1 0 19964 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_230
timestamp 18001
transform 1 0 22264 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_240
timestamp 18001
transform 1 0 23184 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_248
timestamp 18001
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1636986456
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1636986456
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1636986456
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_289
timestamp 18001
transform 1 0 27692 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_305
timestamp 18001
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_322
timestamp 1636986456
transform 1 0 30728 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_334
timestamp 1636986456
transform 1 0 31832 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_346
timestamp 1636986456
transform 1 0 32936 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_358
timestamp 18001
transform 1 0 34040 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1636986456
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_377
timestamp 18001
transform 1 0 35788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_3
timestamp 18001
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_9
timestamp 18001
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1636986456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1636986456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 18001
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 18001
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_57
timestamp 18001
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_67
timestamp 18001
transform 1 0 7268 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_84
timestamp 18001
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_135
timestamp 18001
transform 1 0 13524 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_141
timestamp 1636986456
transform 1 0 14076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_153
timestamp 1636986456
transform 1 0 15180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 18001
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1636986456
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1636986456
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1636986456
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_205
timestamp 18001
transform 1 0 19964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 18001
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 18001
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_237
timestamp 18001
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_243
timestamp 18001
transform 1 0 23460 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_259
timestamp 18001
transform 1 0 24932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_269
timestamp 18001
transform 1 0 25852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_274
timestamp 18001
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_281
timestamp 18001
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_291
timestamp 1636986456
transform 1 0 27876 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_303
timestamp 1636986456
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_315
timestamp 1636986456
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_327
timestamp 18001
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 18001
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_351
timestamp 18001
transform 1 0 33396 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_359
timestamp 18001
transform 1 0 34132 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_377
timestamp 18001
transform 1 0 35788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_23
timestamp 18001
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 18001
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_29
timestamp 18001
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_42
timestamp 1636986456
transform 1 0 4968 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_54
timestamp 18001
transform 1 0 6072 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_60
timestamp 18001
transform 1 0 6624 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_70
timestamp 18001
transform 1 0 7544 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_79
timestamp 18001
transform 1 0 8372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_113
timestamp 18001
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 18001
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_141
timestamp 18001
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_149
timestamp 18001
transform 1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_165
timestamp 18001
transform 1 0 16284 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_178
timestamp 18001
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_188
timestamp 18001
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1636986456
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_209
timestamp 18001
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_217
timestamp 18001
transform 1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_227
timestamp 18001
transform 1 0 21988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 18001
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_260
timestamp 18001
transform 1 0 25024 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_264
timestamp 18001
transform 1 0 25392 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_283
timestamp 18001
transform 1 0 27140 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_295
timestamp 1636986456
transform 1 0 28244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 18001
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_317
timestamp 18001
transform 1 0 30268 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_328
timestamp 1636986456
transform 1 0 31280 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_340
timestamp 1636986456
transform 1 0 32384 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_352
timestamp 1636986456
transform 1 0 33488 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_371
timestamp 18001
transform 1 0 35236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_379
timestamp 18001
transform 1 0 35972 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_3
timestamp 18001
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_9
timestamp 18001
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_34
timestamp 18001
transform 1 0 4232 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_42
timestamp 18001
transform 1 0 4968 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_52
timestamp 18001
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_85
timestamp 18001
transform 1 0 8924 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_108
timestamp 18001
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_121
timestamp 18001
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_132
timestamp 18001
transform 1 0 13248 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_148
timestamp 18001
transform 1 0 14720 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_175
timestamp 1636986456
transform 1 0 17204 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_187
timestamp 18001
transform 1 0 18308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_192
timestamp 18001
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_211
timestamp 1636986456
transform 1 0 20516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 18001
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_225
timestamp 18001
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_244
timestamp 18001
transform 1 0 23552 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_248
timestamp 18001
transform 1 0 23920 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_255
timestamp 18001
transform 1 0 24564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_259
timestamp 18001
transform 1 0 24932 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_266
timestamp 1636986456
transform 1 0 25576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 18001
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_281
timestamp 18001
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_289
timestamp 18001
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_299
timestamp 1636986456
transform 1 0 28612 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_311
timestamp 1636986456
transform 1 0 29716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_323
timestamp 1636986456
transform 1 0 30820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 18001
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_337
timestamp 18001
transform 1 0 32108 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_343
timestamp 18001
transform 1 0 32660 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1636986456
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1636986456
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_373
timestamp 18001
transform 1 0 35420 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_23
timestamp 18001
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_36
timestamp 18001
transform 1 0 4416 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_42
timestamp 18001
transform 1 0 4968 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 18001
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_92
timestamp 18001
transform 1 0 9568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_113
timestamp 18001
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_137
timestamp 18001
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_141
timestamp 18001
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_169
timestamp 18001
transform 1 0 16652 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_176
timestamp 18001
transform 1 0 17296 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_184
timestamp 18001
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_191
timestamp 18001
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 18001
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_225
timestamp 1636986456
transform 1 0 21804 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_237
timestamp 1636986456
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_249
timestamp 18001
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1636986456
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_265
timestamp 18001
transform 1 0 25484 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_272
timestamp 1636986456
transform 1 0 26128 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_284
timestamp 18001
transform 1 0 27232 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_297
timestamp 18001
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_305
timestamp 18001
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_315
timestamp 1636986456
transform 1 0 30084 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_327
timestamp 1636986456
transform 1 0 31188 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_339
timestamp 1636986456
transform 1 0 32292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_351
timestamp 18001
transform 1 0 33396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_355
timestamp 18001
transform 1 0 33764 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_362
timestamp 18001
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1636986456
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_377
timestamp 18001
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636986456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1636986456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_27
timestamp 18001
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_50
timestamp 18001
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_57
timestamp 18001
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_77
timestamp 18001
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_107
timestamp 18001
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 18001
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_122
timestamp 18001
transform 1 0 12328 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 18001
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1636986456
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_193
timestamp 18001
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_201
timestamp 18001
transform 1 0 19596 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_210
timestamp 18001
transform 1 0 20424 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_214
timestamp 18001
transform 1 0 20792 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 18001
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_231
timestamp 18001
transform 1 0 22356 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_235
timestamp 18001
transform 1 0 22724 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_239
timestamp 18001
transform 1 0 23092 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_252
timestamp 18001
transform 1 0 24288 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_258
timestamp 18001
transform 1 0 24840 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_264
timestamp 18001
transform 1 0 25392 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_298
timestamp 1636986456
transform 1 0 28520 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_310
timestamp 18001
transform 1 0 29624 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_316
timestamp 18001
transform 1 0 30176 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_323
timestamp 18001
transform 1 0 30820 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_333
timestamp 18001
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1636986456
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1636986456
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_361
timestamp 18001
transform 1 0 34316 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_369
timestamp 1636986456
transform 1 0 35052 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_3
timestamp 18001
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 18001
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 18001
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_37
timestamp 18001
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_45
timestamp 1636986456
transform 1 0 5244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_57
timestamp 18001
transform 1 0 6348 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 18001
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_144
timestamp 18001
transform 1 0 14352 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_150
timestamp 18001
transform 1 0 14904 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_158
timestamp 18001
transform 1 0 15640 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_167
timestamp 18001
transform 1 0 16468 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1636986456
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 18001
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 18001
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_203
timestamp 1636986456
transform 1 0 19780 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_215
timestamp 18001
transform 1 0 20884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_224
timestamp 18001
transform 1 0 21712 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_228
timestamp 18001
transform 1 0 22080 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_266
timestamp 18001
transform 1 0 25576 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_283
timestamp 18001
transform 1 0 27140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_291
timestamp 18001
transform 1 0 27876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_300
timestamp 18001
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1636986456
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_321
timestamp 18001
transform 1 0 30636 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_327
timestamp 18001
transform 1 0 31188 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_334
timestamp 18001
transform 1 0 31832 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_342
timestamp 18001
transform 1 0 32568 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_350
timestamp 1636986456
transform 1 0 33304 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_362
timestamp 18001
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1636986456
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_377
timestamp 18001
transform 1 0 35788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_31
timestamp 18001
transform 1 0 3956 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1636986456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 18001
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 18001
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_120
timestamp 18001
transform 1 0 12144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_128
timestamp 18001
transform 1 0 12880 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_143
timestamp 1636986456
transform 1 0 14260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_155
timestamp 1636986456
transform 1 0 15364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 18001
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_169
timestamp 18001
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_179
timestamp 18001
transform 1 0 17572 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_185
timestamp 18001
transform 1 0 18124 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_194
timestamp 18001
transform 1 0 18952 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_211
timestamp 1636986456
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 18001
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636986456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_237
timestamp 18001
transform 1 0 22908 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_250
timestamp 1636986456
transform 1 0 24104 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_262
timestamp 1636986456
transform 1 0 25208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_274
timestamp 18001
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1636986456
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_293
timestamp 18001
transform 1 0 28060 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_313
timestamp 1636986456
transform 1 0 29900 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_325
timestamp 18001
transform 1 0 31004 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 18001
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1636986456
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1636986456
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 1636986456
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_373
timestamp 18001
transform 1 0 35420 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 18001
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_11
timestamp 18001
transform 1 0 2116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_22
timestamp 18001
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_37
timestamp 18001
transform 1 0 4508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_48
timestamp 18001
transform 1 0 5520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_65
timestamp 18001
transform 1 0 7084 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_80
timestamp 18001
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_85
timestamp 18001
transform 1 0 8924 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_106
timestamp 18001
transform 1 0 10856 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_127
timestamp 18001
transform 1 0 12788 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 18001
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_141
timestamp 18001
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_164
timestamp 18001
transform 1 0 16192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_170
timestamp 18001
transform 1 0 16744 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_178
timestamp 1636986456
transform 1 0 17480 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_190
timestamp 18001
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_197
timestamp 18001
transform 1 0 19228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_207
timestamp 18001
transform 1 0 20148 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_215
timestamp 18001
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_225
timestamp 18001
transform 1 0 21804 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_233
timestamp 18001
transform 1 0 22540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_244
timestamp 18001
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1636986456
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_265
timestamp 18001
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_276
timestamp 18001
transform 1 0 26496 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_296
timestamp 1636986456
transform 1 0 28336 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_309
timestamp 18001
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_313
timestamp 18001
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1636986456
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1636986456
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1636986456
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 18001
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 18001
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_365
timestamp 18001
transform 1 0 34684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_369
timestamp 18001
transform 1 0 35052 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_3
timestamp 18001
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_64
timestamp 18001
transform 1 0 6992 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_129
timestamp 18001
transform 1 0 12972 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_148
timestamp 18001
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_158
timestamp 18001
transform 1 0 15640 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_164
timestamp 18001
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1636986456
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_181
timestamp 18001
transform 1 0 17756 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_190
timestamp 1636986456
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_202
timestamp 18001
transform 1 0 19688 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_216
timestamp 18001
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_225
timestamp 18001
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_234
timestamp 18001
transform 1 0 22632 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_255
timestamp 18001
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_263
timestamp 18001
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_269
timestamp 18001
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 18001
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_281
timestamp 18001
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_300
timestamp 1636986456
transform 1 0 28704 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_312
timestamp 1636986456
transform 1 0 29808 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_324
timestamp 1636986456
transform 1 0 30912 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_345
timestamp 18001
transform 1 0 32844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_349
timestamp 18001
transform 1 0 33212 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_355
timestamp 18001
transform 1 0 33764 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_369
timestamp 18001
transform 1 0 35052 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 18001
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_38
timestamp 18001
transform 1 0 4600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_57
timestamp 18001
transform 1 0 6348 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_73
timestamp 18001
transform 1 0 7820 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1636986456
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_97
timestamp 18001
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 18001
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_141
timestamp 18001
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_164
timestamp 18001
transform 1 0 16192 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_170
timestamp 18001
transform 1 0 16744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_182
timestamp 18001
transform 1 0 17848 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_192
timestamp 18001
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1636986456
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1636986456
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_221
timestamp 18001
transform 1 0 21436 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_233
timestamp 18001
transform 1 0 22540 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_240
timestamp 1636986456
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1636986456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_265
timestamp 18001
transform 1 0 25484 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_271
timestamp 1636986456
transform 1 0 26036 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_283
timestamp 18001
transform 1 0 27140 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_298
timestamp 18001
transform 1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 18001
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1636986456
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1636986456
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1636986456
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1636986456
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 18001
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 18001
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1636986456
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_377
timestamp 18001
transform 1 0 35788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_3
timestamp 18001
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_65
timestamp 18001
transform 1 0 7084 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_87
timestamp 1636986456
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_99
timestamp 1636986456
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 18001
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_118
timestamp 18001
transform 1 0 11960 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_126
timestamp 18001
transform 1 0 12696 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1636986456
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_149
timestamp 18001
transform 1 0 14812 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_160
timestamp 18001
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_169
timestamp 18001
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_177
timestamp 18001
transform 1 0 17388 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_197
timestamp 18001
transform 1 0 19228 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_212
timestamp 18001
transform 1 0 20608 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 18001
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_225
timestamp 18001
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_229
timestamp 18001
transform 1 0 22172 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_235
timestamp 1636986456
transform 1 0 22724 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_247
timestamp 1636986456
transform 1 0 23828 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_259
timestamp 18001
transform 1 0 24932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_266
timestamp 18001
transform 1 0 25576 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_274
timestamp 18001
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1636986456
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_293
timestamp 18001
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_297
timestamp 18001
transform 1 0 28428 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_310
timestamp 18001
transform 1 0 29624 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_318
timestamp 18001
transform 1 0 30360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_328
timestamp 18001
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_337
timestamp 18001
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_345
timestamp 18001
transform 1 0 32844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_353
timestamp 18001
transform 1 0 33580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_361
timestamp 18001
transform 1 0 34316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_368
timestamp 1636986456
transform 1 0 34960 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_380
timestamp 18001
transform 1 0 36064 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_23
timestamp 18001
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 18001
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_29
timestamp 18001
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_37
timestamp 18001
transform 1 0 4508 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_54
timestamp 18001
transform 1 0 6072 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_79
timestamp 18001
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 18001
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_85
timestamp 18001
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_105
timestamp 18001
transform 1 0 10764 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_115
timestamp 18001
transform 1 0 11684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_119
timestamp 18001
transform 1 0 12052 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_126
timestamp 18001
transform 1 0 12696 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 18001
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 18001
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_156
timestamp 1636986456
transform 1 0 15456 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_168
timestamp 18001
transform 1 0 16560 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_180
timestamp 1636986456
transform 1 0 17664 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 18001
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_205
timestamp 18001
transform 1 0 19964 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_223
timestamp 1636986456
transform 1 0 21620 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_235
timestamp 1636986456
transform 1 0 22724 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_247
timestamp 18001
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 18001
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_264
timestamp 18001
transform 1 0 25392 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_270
timestamp 18001
transform 1 0 25944 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_292
timestamp 1636986456
transform 1 0 27968 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_304
timestamp 18001
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1636986456
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_334
timestamp 1636986456
transform 1 0 31832 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_346
timestamp 1636986456
transform 1 0 32936 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_358
timestamp 18001
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1636986456
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_377
timestamp 18001
transform 1 0 35788 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_3
timestamp 18001
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_11
timestamp 18001
transform 1 0 2116 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_21
timestamp 18001
transform 1 0 3036 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_27
timestamp 18001
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_62
timestamp 18001
transform 1 0 6808 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_66
timestamp 1636986456
transform 1 0 7176 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_78
timestamp 18001
transform 1 0 8280 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_83
timestamp 18001
transform 1 0 8740 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_95
timestamp 1636986456
transform 1 0 9844 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_107
timestamp 18001
transform 1 0 10948 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_131
timestamp 1636986456
transform 1 0 13156 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_143
timestamp 1636986456
transform 1 0 14260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_155
timestamp 18001
transform 1 0 15364 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_163
timestamp 18001
transform 1 0 16100 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_178
timestamp 18001
transform 1 0 17480 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_184
timestamp 18001
transform 1 0 18032 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_202
timestamp 1636986456
transform 1 0 19688 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_214
timestamp 18001
transform 1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_222
timestamp 18001
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_225
timestamp 18001
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_233
timestamp 18001
transform 1 0 22540 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1636986456
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_261
timestamp 18001
transform 1 0 25116 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_275
timestamp 18001
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 18001
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_281
timestamp 18001
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_290
timestamp 18001
transform 1 0 27784 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_308
timestamp 1636986456
transform 1 0 29440 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_320
timestamp 1636986456
transform 1 0 30544 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_332
timestamp 18001
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1636986456
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_349
timestamp 18001
transform 1 0 33212 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_355
timestamp 18001
transform 1 0 33764 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_361
timestamp 18001
transform 1 0 34316 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_369
timestamp 18001
transform 1 0 35052 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_23
timestamp 18001
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 18001
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_53
timestamp 18001
transform 1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_57
timestamp 18001
transform 1 0 6348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_64
timestamp 18001
transform 1 0 6992 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_69
timestamp 18001
transform 1 0 7452 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_73
timestamp 18001
transform 1 0 7820 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_81
timestamp 18001
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_85
timestamp 18001
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_98
timestamp 1636986456
transform 1 0 10120 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_110
timestamp 18001
transform 1 0 11224 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_118
timestamp 1636986456
transform 1 0 11960 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_130
timestamp 18001
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 18001
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_141
timestamp 18001
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_156
timestamp 18001
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_171
timestamp 18001
transform 1 0 16836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_186
timestamp 18001
transform 1 0 18216 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_197
timestamp 18001
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_216
timestamp 18001
transform 1 0 20976 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_231
timestamp 18001
transform 1 0 22356 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_244
timestamp 18001
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_253
timestamp 18001
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_257
timestamp 18001
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_264
timestamp 1636986456
transform 1 0 25392 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_276
timestamp 1636986456
transform 1 0 26496 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_288
timestamp 1636986456
transform 1 0 27600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_300
timestamp 18001
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1636986456
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1636986456
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_333
timestamp 18001
transform 1 0 31740 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_345
timestamp 18001
transform 1 0 32844 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_349
timestamp 18001
transform 1 0 33212 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_359
timestamp 18001
transform 1 0 34132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 18001
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_365
timestamp 18001
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_373
timestamp 18001
transform 1 0 35420 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_380
timestamp 18001
transform 1 0 36064 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_3
timestamp 18001
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_57
timestamp 18001
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_75
timestamp 18001
transform 1 0 8004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_99
timestamp 18001
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_110
timestamp 18001
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_120
timestamp 18001
transform 1 0 12144 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_130
timestamp 18001
transform 1 0 13064 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_154
timestamp 18001
transform 1 0 15272 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 18001
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_169
timestamp 18001
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_191
timestamp 18001
transform 1 0 18676 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_201
timestamp 18001
transform 1 0 19596 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_205
timestamp 18001
transform 1 0 19964 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 18001
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_232
timestamp 18001
transform 1 0 22448 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_259
timestamp 18001
transform 1 0 24932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_272
timestamp 18001
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_281
timestamp 18001
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_290
timestamp 1636986456
transform 1 0 27784 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_316
timestamp 1636986456
transform 1 0 30176 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_328
timestamp 18001
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_345
timestamp 18001
transform 1 0 32844 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_351
timestamp 18001
transform 1 0 33396 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_23
timestamp 18001
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 18001
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_38
timestamp 18001
transform 1 0 4600 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_57
timestamp 18001
transform 1 0 6348 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_65
timestamp 18001
transform 1 0 7084 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_74
timestamp 18001
transform 1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_82
timestamp 18001
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1636986456
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_97
timestamp 18001
transform 1 0 10028 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_105
timestamp 18001
transform 1 0 10764 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_111
timestamp 18001
transform 1 0 11316 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_115
timestamp 18001
transform 1 0 11684 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_123
timestamp 18001
transform 1 0 12420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_138
timestamp 18001
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_146
timestamp 18001
transform 1 0 14536 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_154
timestamp 18001
transform 1 0 15272 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_181
timestamp 18001
transform 1 0 17756 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_187
timestamp 18001
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 18001
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 18001
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_215
timestamp 18001
transform 1 0 20884 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_223
timestamp 18001
transform 1 0 21620 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_231
timestamp 18001
transform 1 0 22356 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_239
timestamp 18001
transform 1 0 23092 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 18001
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 18001
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_253
timestamp 18001
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_261
timestamp 18001
transform 1 0 25116 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_279
timestamp 18001
transform 1 0 26772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_288
timestamp 18001
transform 1 0 27600 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_297
timestamp 18001
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_305
timestamp 18001
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_316
timestamp 1636986456
transform 1 0 30176 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_328
timestamp 18001
transform 1 0 31280 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_341
timestamp 1636986456
transform 1 0 32476 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_353
timestamp 18001
transform 1 0 33580 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_361
timestamp 18001
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1636986456
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_377
timestamp 18001
transform 1 0 35788 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_3
timestamp 18001
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_11
timestamp 18001
transform 1 0 2116 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_32
timestamp 18001
transform 1 0 4048 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_45
timestamp 18001
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_53
timestamp 18001
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_57
timestamp 18001
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_76
timestamp 18001
transform 1 0 8096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_84
timestamp 18001
transform 1 0 8832 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_90
timestamp 1636986456
transform 1 0 9384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_102
timestamp 18001
transform 1 0 10488 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_113
timestamp 18001
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_119
timestamp 18001
transform 1 0 12052 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_132
timestamp 18001
transform 1 0 13248 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_140
timestamp 18001
transform 1 0 13984 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_151
timestamp 1636986456
transform 1 0 14996 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_163
timestamp 18001
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 18001
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_179
timestamp 18001
transform 1 0 17572 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_183
timestamp 18001
transform 1 0 17940 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 18001
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_225
timestamp 18001
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_257
timestamp 1636986456
transform 1 0 24748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_277
timestamp 18001
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_281
timestamp 18001
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_285
timestamp 18001
transform 1 0 27324 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_291
timestamp 1636986456
transform 1 0 27876 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_303
timestamp 1636986456
transform 1 0 28980 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_315
timestamp 1636986456
transform 1 0 30084 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_327
timestamp 18001
transform 1 0 31188 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 18001
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1636986456
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1636986456
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_361
timestamp 18001
transform 1 0 34316 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_371
timestamp 18001
transform 1 0 35236 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_379
timestamp 18001
transform 1 0 35972 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_3
timestamp 18001
transform 1 0 1380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_11
timestamp 18001
transform 1 0 2116 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_18
timestamp 18001
transform 1 0 2760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_26
timestamp 18001
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_29
timestamp 18001
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_33
timestamp 18001
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_58
timestamp 18001
transform 1 0 6440 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_66
timestamp 18001
transform 1 0 7176 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_76
timestamp 18001
transform 1 0 8096 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_92
timestamp 18001
transform 1 0 9568 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_98
timestamp 18001
transform 1 0 10120 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_102
timestamp 18001
transform 1 0 10488 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_106
timestamp 18001
transform 1 0 10856 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 18001
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_141
timestamp 18001
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_158
timestamp 1636986456
transform 1 0 15640 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_170
timestamp 18001
transform 1 0 16744 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_194
timestamp 18001
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_215
timestamp 18001
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 18001
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_253
timestamp 18001
transform 1 0 24380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_262
timestamp 18001
transform 1 0 25208 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_284
timestamp 1636986456
transform 1 0 27232 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_296
timestamp 1636986456
transform 1 0 28336 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_316
timestamp 18001
transform 1 0 30176 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_330
timestamp 18001
transform 1 0 31464 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_337
timestamp 1636986456
transform 1 0 32108 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_349
timestamp 1636986456
transform 1 0 33212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_361
timestamp 18001
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1636986456
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_377
timestamp 18001
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_26
timestamp 18001
transform 1 0 3496 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_32
timestamp 18001
transform 1 0 4048 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_57
timestamp 18001
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_72
timestamp 18001
transform 1 0 7728 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_91
timestamp 18001
transform 1 0 9476 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_101
timestamp 18001
transform 1 0 10396 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 18001
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_165
timestamp 18001
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_169
timestamp 18001
transform 1 0 16652 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_177
timestamp 18001
transform 1 0 17388 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_185
timestamp 18001
transform 1 0 18124 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_205
timestamp 18001
transform 1 0 19964 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_219
timestamp 18001
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 18001
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_225
timestamp 18001
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_241
timestamp 18001
transform 1 0 23276 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_278
timestamp 18001
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_290
timestamp 18001
transform 1 0 27784 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_296
timestamp 18001
transform 1 0 28336 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_305
timestamp 18001
transform 1 0 29164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_309
timestamp 18001
transform 1 0 29532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_325
timestamp 18001
transform 1 0 31004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_329
timestamp 18001
transform 1 0 31372 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_337
timestamp 18001
transform 1 0 32108 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_347
timestamp 1636986456
transform 1 0 33028 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_359
timestamp 1636986456
transform 1 0 34132 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_371
timestamp 18001
transform 1 0 35236 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_379
timestamp 18001
transform 1 0 35972 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_3
timestamp 18001
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_35
timestamp 18001
transform 1 0 4324 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_39
timestamp 18001
transform 1 0 4692 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_63
timestamp 18001
transform 1 0 6900 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_85
timestamp 18001
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_109
timestamp 18001
transform 1 0 11132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_158
timestamp 18001
transform 1 0 15640 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_169
timestamp 1636986456
transform 1 0 16652 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_181
timestamp 18001
transform 1 0 17756 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_189
timestamp 18001
transform 1 0 18492 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 18001
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_197
timestamp 18001
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_205
timestamp 18001
transform 1 0 19964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_218
timestamp 18001
transform 1 0 21160 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_257
timestamp 18001
transform 1 0 24748 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_281
timestamp 18001
transform 1 0 26956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1636986456
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_321
timestamp 18001
transform 1 0 30636 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_329
timestamp 18001
transform 1 0 31372 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_339
timestamp 1636986456
transform 1 0 32292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_351
timestamp 18001
transform 1 0 33396 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 18001
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_373
timestamp 18001
transform 1 0 35420 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_3
timestamp 18001
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1636986456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 18001
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 18001
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 18001
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_75
timestamp 1636986456
transform 1 0 8004 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_100
timestamp 1636986456
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_113
timestamp 18001
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_163
timestamp 18001
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 18001
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_183
timestamp 18001
transform 1 0 17940 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1636986456
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_205
timestamp 18001
transform 1 0 19964 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_222
timestamp 18001
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_231
timestamp 18001
transform 1 0 22356 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_245
timestamp 18001
transform 1 0 23644 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_277
timestamp 18001
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_289
timestamp 18001
transform 1 0 27692 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_303
timestamp 18001
transform 1 0 28980 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_310
timestamp 18001
transform 1 0 29624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_316
timestamp 18001
transform 1 0 30176 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_333
timestamp 18001
transform 1 0 31740 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1636986456
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1636986456
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_361
timestamp 18001
transform 1 0 34316 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_379
timestamp 18001
transform 1 0 35972 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_3
timestamp 18001
transform 1 0 1380 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 18001
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_38
timestamp 18001
transform 1 0 4600 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_52
timestamp 1636986456
transform 1 0 5888 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_64
timestamp 18001
transform 1 0 6992 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_79
timestamp 18001
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 18001
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_94
timestamp 18001
transform 1 0 9752 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_98
timestamp 18001
transform 1 0 10120 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_105
timestamp 18001
transform 1 0 10764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_113
timestamp 18001
transform 1 0 11500 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_147
timestamp 18001
transform 1 0 14628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_153
timestamp 18001
transform 1 0 15180 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_169
timestamp 18001
transform 1 0 16652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_175
timestamp 18001
transform 1 0 17204 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_183
timestamp 18001
transform 1 0 17940 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_194
timestamp 18001
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_204
timestamp 18001
transform 1 0 19872 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_221
timestamp 18001
transform 1 0 21436 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_250
timestamp 18001
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_253
timestamp 18001
transform 1 0 24380 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_284
timestamp 18001
transform 1 0 27232 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_296
timestamp 1636986456
transform 1 0 28336 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1636986456
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_321
timestamp 18001
transform 1 0 30636 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_340
timestamp 1636986456
transform 1 0 32384 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_352
timestamp 1636986456
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1636986456
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_377
timestamp 18001
transform 1 0 35788 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_3
timestamp 18001
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 18001
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_57
timestamp 18001
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_65
timestamp 18001
transform 1 0 7084 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_77
timestamp 18001
transform 1 0 8188 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_81
timestamp 18001
transform 1 0 8556 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_89
timestamp 18001
transform 1 0 9292 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_93
timestamp 18001
transform 1 0 9660 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 18001
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_119
timestamp 18001
transform 1 0 12052 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_127
timestamp 18001
transform 1 0 12788 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_137
timestamp 18001
transform 1 0 13708 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_143
timestamp 18001
transform 1 0 14260 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_151
timestamp 1636986456
transform 1 0 14996 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_163
timestamp 18001
transform 1 0 16100 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 18001
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_169
timestamp 18001
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_177
timestamp 18001
transform 1 0 17388 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_203
timestamp 1636986456
transform 1 0 19780 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_215
timestamp 18001
transform 1 0 20884 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 18001
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_225
timestamp 18001
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 18001
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_292
timestamp 18001
transform 1 0 27968 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_315
timestamp 18001
transform 1 0 30084 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_324
timestamp 1636986456
transform 1 0 30912 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_337
timestamp 18001
transform 1 0 32108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_345
timestamp 18001
transform 1 0 32844 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_355
timestamp 18001
transform 1 0 33764 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_363
timestamp 1636986456
transform 1 0 34500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_375
timestamp 18001
transform 1 0 35604 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_3
timestamp 18001
transform 1 0 1380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 18001
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_64
timestamp 18001
transform 1 0 6992 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_80
timestamp 18001
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_85
timestamp 18001
transform 1 0 8924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_95
timestamp 18001
transform 1 0 9844 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_118
timestamp 1636986456
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_130
timestamp 18001
transform 1 0 13064 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_150
timestamp 18001
transform 1 0 14904 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_158
timestamp 18001
transform 1 0 15640 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_175
timestamp 18001
transform 1 0 17204 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_179
timestamp 18001
transform 1 0 17572 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_185
timestamp 18001
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_189
timestamp 18001
transform 1 0 18492 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_205
timestamp 1636986456
transform 1 0 19964 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_217
timestamp 18001
transform 1 0 21068 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_256
timestamp 18001
transform 1 0 24656 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_278
timestamp 18001
transform 1 0 26680 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_297
timestamp 18001
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_314
timestamp 18001
transform 1 0 29992 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_329
timestamp 1636986456
transform 1 0 31372 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_341
timestamp 1636986456
transform 1 0 32476 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_353
timestamp 18001
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_361
timestamp 18001
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1636986456
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_377
timestamp 18001
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_3
timestamp 18001
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_7
timestamp 18001
transform 1 0 1748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_54
timestamp 18001
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_62
timestamp 18001
transform 1 0 6808 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_84
timestamp 18001
transform 1 0 8832 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_91
timestamp 18001
transform 1 0 9476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_100
timestamp 18001
transform 1 0 10304 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_108
timestamp 18001
transform 1 0 11040 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_125
timestamp 18001
transform 1 0 12604 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_157
timestamp 18001
transform 1 0 15548 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_165
timestamp 18001
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_169
timestamp 18001
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_177
timestamp 1636986456
transform 1 0 17388 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_189
timestamp 18001
transform 1 0 18492 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_196
timestamp 18001
transform 1 0 19136 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_202
timestamp 18001
transform 1 0 19688 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_221
timestamp 18001
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1636986456
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_295
timestamp 18001
transform 1 0 28244 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_313
timestamp 18001
transform 1 0 29900 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_330
timestamp 18001
transform 1 0 31464 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_337
timestamp 18001
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_353
timestamp 1636986456
transform 1 0 33580 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_365
timestamp 1636986456
transform 1 0 34684 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_377
timestamp 18001
transform 1 0 35788 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_3
timestamp 18001
transform 1 0 1380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_11
timestamp 18001
transform 1 0 2116 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_19
timestamp 18001
transform 1 0 2852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_64
timestamp 18001
transform 1 0 6992 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_77
timestamp 18001
transform 1 0 8188 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 18001
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_85
timestamp 18001
transform 1 0 8924 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_98
timestamp 18001
transform 1 0 10120 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_134
timestamp 18001
transform 1 0 13432 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 18001
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_141
timestamp 18001
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_149
timestamp 18001
transform 1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_160
timestamp 1636986456
transform 1 0 15824 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_172
timestamp 18001
transform 1 0 16928 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_178
timestamp 18001
transform 1 0 17480 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_183
timestamp 1636986456
transform 1 0 17940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 18001
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_197
timestamp 18001
transform 1 0 19228 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1636986456
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_228
timestamp 18001
transform 1 0 22080 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_278
timestamp 18001
transform 1 0 26680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_290
timestamp 18001
transform 1 0 27784 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_299
timestamp 18001
transform 1 0 28612 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_306
timestamp 18001
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_320
timestamp 18001
transform 1 0 30544 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_331
timestamp 18001
transform 1 0 31556 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_335
timestamp 18001
transform 1 0 31924 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_339
timestamp 18001
transform 1 0 32292 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1636986456
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 18001
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 18001
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1636986456
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_377
timestamp 18001
transform 1 0 35788 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_3
timestamp 18001
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1636986456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_39
timestamp 18001
transform 1 0 4692 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_54
timestamp 18001
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_76
timestamp 18001
transform 1 0 8096 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_82
timestamp 18001
transform 1 0 8648 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_109
timestamp 18001
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_113
timestamp 18001
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_124
timestamp 1636986456
transform 1 0 12512 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_136
timestamp 1636986456
transform 1 0 13616 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_148
timestamp 18001
transform 1 0 14720 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_154
timestamp 18001
transform 1 0 15272 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_169
timestamp 18001
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_177
timestamp 18001
transform 1 0 17388 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_189
timestamp 18001
transform 1 0 18492 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_193
timestamp 18001
transform 1 0 18860 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_210
timestamp 18001
transform 1 0 20424 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_218
timestamp 18001
transform 1 0 21160 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_233
timestamp 18001
transform 1 0 22540 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_256
timestamp 18001
transform 1 0 24656 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_301
timestamp 18001
transform 1 0 28796 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_337
timestamp 18001
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_352
timestamp 1636986456
transform 1 0 33488 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_364
timestamp 1636986456
transform 1 0 34592 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_376
timestamp 18001
transform 1 0 35696 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_380
timestamp 18001
transform 1 0 36064 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1636986456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1636986456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 18001
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_29
timestamp 18001
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_52
timestamp 18001
transform 1 0 5888 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_71
timestamp 18001
transform 1 0 7636 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_80
timestamp 18001
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_85
timestamp 18001
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_92
timestamp 18001
transform 1 0 9568 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_101
timestamp 18001
transform 1 0 10396 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_107
timestamp 18001
transform 1 0 10948 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_111
timestamp 18001
transform 1 0 11316 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_115
timestamp 18001
transform 1 0 11684 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1636986456
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 18001
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 18001
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_164
timestamp 1636986456
transform 1 0 16192 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_176
timestamp 1636986456
transform 1 0 17296 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_188
timestamp 18001
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_210
timestamp 1636986456
transform 1 0 20424 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_222
timestamp 18001
transform 1 0 21528 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_286
timestamp 18001
transform 1 0 27416 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 18001
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_349
timestamp 1636986456
transform 1 0 33212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_361
timestamp 18001
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1636986456
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_377
timestamp 18001
transform 1 0 35788 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1636986456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1636986456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1636986456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_39
timestamp 18001
transform 1 0 4692 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_64
timestamp 18001
transform 1 0 6992 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_103
timestamp 18001
transform 1 0 10580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_128
timestamp 18001
transform 1 0 12880 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_159
timestamp 18001
transform 1 0 15732 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 18001
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_173
timestamp 18001
transform 1 0 17020 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_187
timestamp 18001
transform 1 0 18308 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_196
timestamp 18001
transform 1 0 19136 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_253
timestamp 18001
transform 1 0 24380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_333
timestamp 18001
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_357
timestamp 1636986456
transform 1 0 33948 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_369
timestamp 1636986456
transform 1 0 35052 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1636986456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_29
timestamp 18001
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_37
timestamp 18001
transform 1 0 4508 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_74
timestamp 18001
transform 1 0 7912 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 18001
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_85
timestamp 18001
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_89
timestamp 18001
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_101
timestamp 18001
transform 1 0 10396 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_118
timestamp 18001
transform 1 0 11960 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_179
timestamp 18001
transform 1 0 17572 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 18001
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_218
timestamp 18001
transform 1 0 21160 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_222
timestamp 18001
transform 1 0 21528 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_294
timestamp 18001
transform 1 0 28152 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_304
timestamp 18001
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_319
timestamp 1636986456
transform 1 0 30452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_331
timestamp 18001
transform 1 0 31556 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_339
timestamp 18001
transform 1 0 32292 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1636986456
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 18001
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 18001
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1636986456
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_377
timestamp 18001
transform 1 0 35788 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1636986456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1636986456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1636986456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1636986456
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_51
timestamp 18001
transform 1 0 5796 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_57
timestamp 18001
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_75
timestamp 18001
transform 1 0 8004 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_83
timestamp 18001
transform 1 0 8740 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_89
timestamp 18001
transform 1 0 9292 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_98
timestamp 1636986456
transform 1 0 10120 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_110
timestamp 18001
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_113
timestamp 18001
transform 1 0 11500 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_131
timestamp 1636986456
transform 1 0 13156 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_143
timestamp 18001
transform 1 0 14260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_151
timestamp 18001
transform 1 0 14996 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_160
timestamp 18001
transform 1 0 15824 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_200
timestamp 18001
transform 1 0 19504 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_225
timestamp 18001
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_256
timestamp 18001
transform 1 0 24656 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_277
timestamp 18001
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_281
timestamp 18001
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_285
timestamp 18001
transform 1 0 27324 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_314
timestamp 1636986456
transform 1 0 29992 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_326
timestamp 18001
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_334
timestamp 18001
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1636986456
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1636986456
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1636986456
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_373
timestamp 18001
transform 1 0 35420 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1636986456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1636986456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 18001
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1636986456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_41
timestamp 18001
transform 1 0 4876 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_49
timestamp 18001
transform 1 0 5612 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_62
timestamp 18001
transform 1 0 6808 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_94
timestamp 18001
transform 1 0 9752 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_98
timestamp 18001
transform 1 0 10120 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_124
timestamp 18001
transform 1 0 12512 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_138
timestamp 18001
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_141
timestamp 18001
transform 1 0 14076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_160
timestamp 18001
transform 1 0 15824 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_168
timestamp 18001
transform 1 0 16560 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_183
timestamp 18001
transform 1 0 17940 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_215
timestamp 18001
transform 1 0 20884 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_250
timestamp 18001
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_253
timestamp 18001
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_270
timestamp 1636986456
transform 1 0 25944 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_288
timestamp 1636986456
transform 1 0 27600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_300
timestamp 18001
transform 1 0 28704 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1636986456
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1636986456
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1636986456
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1636986456
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 18001
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 18001
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1636986456
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_377
timestamp 18001
transform 1 0 35788 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1636986456
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1636986456
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1636986456
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1636986456
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 18001
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 18001
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_78
timestamp 18001
transform 1 0 8280 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_82
timestamp 18001
transform 1 0 8648 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_93
timestamp 18001
transform 1 0 9660 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_103
timestamp 18001
transform 1 0 10580 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 18001
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_147
timestamp 18001
transform 1 0 14628 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_178
timestamp 18001
transform 1 0 17480 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_186
timestamp 18001
transform 1 0 18216 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 18001
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_225
timestamp 18001
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_263
timestamp 1636986456
transform 1 0 25300 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_275
timestamp 18001
transform 1 0 26404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 18001
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1636986456
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1636986456
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1636986456
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1636986456
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 18001
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 18001
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1636986456
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1636986456
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1636986456
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_373
timestamp 18001
transform 1 0 35420 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1636986456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1636986456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 18001
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1636986456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1636986456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1636986456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_65
timestamp 18001
transform 1 0 7084 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_69
timestamp 1636986456
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_81
timestamp 18001
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_85
timestamp 18001
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_96
timestamp 18001
transform 1 0 9936 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_121
timestamp 18001
transform 1 0 12236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_203
timestamp 18001
transform 1 0 19780 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 18001
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 18001
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_271
timestamp 1636986456
transform 1 0 26036 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_283
timestamp 1636986456
transform 1 0 27140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_295
timestamp 1636986456
transform 1 0 28244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 18001
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1636986456
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1636986456
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1636986456
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1636986456
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 18001
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 18001
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1636986456
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_377
timestamp 18001
transform 1 0 35788 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1636986456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1636986456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1636986456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 18001
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 18001
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1636986456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1636986456
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_81
timestamp 18001
transform 1 0 8556 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1636986456
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_163
timestamp 18001
transform 1 0 16100 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_182
timestamp 18001
transform 1 0 17848 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_196
timestamp 18001
transform 1 0 19136 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_221
timestamp 18001
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_248
timestamp 1636986456
transform 1 0 23920 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_260
timestamp 1636986456
transform 1 0 25024 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_272
timestamp 18001
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1636986456
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1636986456
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1636986456
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1636986456
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 18001
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 18001
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1636986456
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1636986456
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1636986456
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_373
timestamp 18001
transform 1 0 35420 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1636986456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1636986456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 18001
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1636986456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1636986456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 18001
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 1636986456
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 1636986456
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 18001
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1636986456
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1636986456
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_109
timestamp 18001
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 1636986456
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1636986456
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 18001
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1636986456
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1636986456
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_165
timestamp 18001
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_169
timestamp 18001
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_182
timestamp 1636986456
transform 1 0 17848 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_194
timestamp 18001
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_197
timestamp 18001
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_205
timestamp 18001
transform 1 0 19964 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_216
timestamp 18001
transform 1 0 20976 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_248
timestamp 18001
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1636986456
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1636986456
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_277
timestamp 18001
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_281
timestamp 1636986456
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_293
timestamp 18001
transform 1 0 28060 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_301
timestamp 18001
transform 1 0 28796 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 18001
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_309
timestamp 18001
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_317
timestamp 1636986456
transform 1 0 30268 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_329
timestamp 18001
transform 1 0 31372 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_335
timestamp 18001
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_337
timestamp 1636986456
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_349
timestamp 1636986456
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_361
timestamp 18001
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1636986456
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_377
timestamp 18001
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 18001
transform -1 0 19780 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 18001
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 18001
transform -1 0 28152 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 18001
transform -1 0 16468 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 18001
transform -1 0 16192 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 18001
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 18001
transform -1 0 15088 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 18001
transform -1 0 19136 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 18001
transform 1 0 17388 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 18001
transform -1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 18001
transform -1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 18001
transform -1 0 3956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 18001
transform -1 0 12236 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 18001
transform -1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 18001
transform -1 0 8648 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 18001
transform -1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 18001
transform -1 0 8372 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 18001
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 18001
transform -1 0 11500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 18001
transform -1 0 7636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 18001
transform -1 0 11684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 18001
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 18001
transform -1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 18001
transform -1 0 5336 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 18001
transform -1 0 12144 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 18001
transform -1 0 6072 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 18001
transform 1 0 8740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 18001
transform -1 0 24380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 18001
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 18001
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 18001
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 18001
transform -1 0 8740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 18001
transform -1 0 5336 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 18001
transform 1 0 14720 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 18001
transform -1 0 4784 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 18001
transform -1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 18001
transform 1 0 12420 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 18001
transform 1 0 7912 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 18001
transform -1 0 25208 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 18001
transform -1 0 26220 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 18001
transform -1 0 7820 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 18001
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 18001
transform -1 0 11316 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 18001
transform -1 0 24196 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 18001
transform -1 0 3956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 18001
transform -1 0 10948 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 18001
transform -1 0 8832 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 18001
transform -1 0 11316 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 18001
transform -1 0 5152 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 18001
transform -1 0 12236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 18001
transform -1 0 5152 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 18001
transform 1 0 28336 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 18001
transform -1 0 20884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 18001
transform -1 0 26220 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 18001
transform -1 0 5980 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 18001
transform -1 0 6256 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 18001
transform -1 0 36156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 18001
transform -1 0 36156 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 18001
transform -1 0 36156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 18001
transform 1 0 29716 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 18001
transform 1 0 29072 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 18001
transform 1 0 35236 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 18001
transform -1 0 36156 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 18001
transform -1 0 36156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 18001
transform 1 0 35880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 18001
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 18001
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 18001
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 18001
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 18001
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 18001
transform -1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 18001
transform -1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 18001
transform -1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 18001
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 36432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 36432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 36432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 36432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 36432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 36432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 36432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 36432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 36432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 36432 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 36432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 36432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 36432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 36432 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 36432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 36432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 36432 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 36432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 36432 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 36432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 36432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 36432 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 36432 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 36432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 36432 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 36432 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 36432 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 36432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 36432 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 36432 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 36432 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 36432 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 36432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 36432 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 36432 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 36432 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 36432 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 36432 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 36432 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 36432 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 36432 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 36432 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 36432 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 36432 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 36432 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 36432 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 36432 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 36432 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 36432 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 36432 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 36432 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 36432 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 36432 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 36432 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 36432 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 36432 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 36432 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 36432 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 36432 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 36432 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 36432 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 36432 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 36432 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 36432 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_143
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_144
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_145
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_146
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_147
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_148
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_149
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_150
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_151
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_152
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_153
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_154
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_155
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_156
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_157
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_158
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_159
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_160
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_161
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_162
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_163
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_164
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_165
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_166
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_167
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_168
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_169
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_170
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_171
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_172
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_173
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_174
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_175
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_176
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_177
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_178
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_179
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_180
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_181
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_182
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_183
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_184
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_185
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_186
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_187
timestamp 18001
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_188
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_189
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_190
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_191
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_192
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_193
timestamp 18001
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_194
timestamp 18001
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_195
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_196
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_197
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_198
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_199
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_200
timestamp 18001
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_201
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_202
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_203
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_204
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_205
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_206
timestamp 18001
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_207
timestamp 18001
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_208
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_209
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_210
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_211
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_212
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_213
timestamp 18001
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_214
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_215
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_216
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_217
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_218
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_219
timestamp 18001
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_220
timestamp 18001
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_221
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_222
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_223
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_224
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_225
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_226
timestamp 18001
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_227
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_228
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_229
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_230
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_231
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_232
timestamp 18001
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_233
timestamp 18001
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_234
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_235
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_236
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_237
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_238
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_239
timestamp 18001
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_240
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_241
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_242
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_243
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_244
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_245
timestamp 18001
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_246
timestamp 18001
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_247
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_248
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_249
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_250
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_251
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_252
timestamp 18001
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_253
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_254
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_255
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_256
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_257
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_258
timestamp 18001
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_259
timestamp 18001
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_260
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_261
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_262
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_263
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_264
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_265
timestamp 18001
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_266
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_267
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_268
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_269
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_270
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_271
timestamp 18001
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_272
timestamp 18001
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_273
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_274
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_275
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_276
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_277
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_278
timestamp 18001
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_279
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_280
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_281
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_282
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_283
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_284
timestamp 18001
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_285
timestamp 18001
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_286
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_287
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_288
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_289
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_290
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_291
timestamp 18001
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_292
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_293
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_294
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_295
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_296
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_297
timestamp 18001
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_298
timestamp 18001
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_299
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_300
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_301
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_302
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_303
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_304
timestamp 18001
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_305
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_306
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_307
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_308
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_309
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_310
timestamp 18001
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_311
timestamp 18001
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_312
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_313
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_314
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_315
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_316
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_317
timestamp 18001
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_318
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_319
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_320
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_321
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_322
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_323
timestamp 18001
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_324
timestamp 18001
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_325
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_326
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_327
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_328
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_329
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_330
timestamp 18001
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_331
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_332
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_333
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_334
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_335
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_336
timestamp 18001
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_337
timestamp 18001
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_338
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_339
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_340
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_341
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_342
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_343
timestamp 18001
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_344
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_345
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_346
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_347
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_348
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_349
timestamp 18001
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_350
timestamp 18001
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_351
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_352
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_353
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_354
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_355
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_356
timestamp 18001
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_357
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_358
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_359
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_360
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_361
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_362
timestamp 18001
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_363
timestamp 18001
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_364
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_365
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_366
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_367
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_368
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_369
timestamp 18001
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_370
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_371
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_372
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_373
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_374
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_375
timestamp 18001
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_376
timestamp 18001
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_377
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_378
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_379
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_380
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_381
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_382
timestamp 18001
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_383
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_384
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_385
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_386
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_387
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_388
timestamp 18001
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_389
timestamp 18001
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_390
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_391
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_392
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_393
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_394
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_395
timestamp 18001
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_396
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_397
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_398
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_399
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_400
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_401
timestamp 18001
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_402
timestamp 18001
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_403
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_404
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_405
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_406
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_407
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_408
timestamp 18001
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_409
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_410
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_411
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_412
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_413
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_414
timestamp 18001
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_415
timestamp 18001
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_416
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_417
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_418
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_419
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_420
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_421
timestamp 18001
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_422
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_423
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_424
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_425
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_426
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_427
timestamp 18001
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_428
timestamp 18001
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_429
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_430
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_431
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_432
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_433
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_434
timestamp 18001
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_435
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_436
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_437
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_438
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_439
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_440
timestamp 18001
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_441
timestamp 18001
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_442
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_443
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_444
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_445
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_446
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_447
timestamp 18001
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_448
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_449
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_450
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_451
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_452
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_453
timestamp 18001
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_454
timestamp 18001
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_455
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_456
timestamp 18001
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_457
timestamp 18001
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_458
timestamp 18001
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_459
timestamp 18001
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_460
timestamp 18001
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_461
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_462
timestamp 18001
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_463
timestamp 18001
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_464
timestamp 18001
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_465
timestamp 18001
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_466
timestamp 18001
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_467
timestamp 18001
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_468
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_469
timestamp 18001
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_470
timestamp 18001
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_471
timestamp 18001
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_472
timestamp 18001
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_473
timestamp 18001
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_474
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_475
timestamp 18001
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_476
timestamp 18001
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_477
timestamp 18001
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_478
timestamp 18001
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_479
timestamp 18001
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_480
timestamp 18001
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_481
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_482
timestamp 18001
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_483
timestamp 18001
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_484
timestamp 18001
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_485
timestamp 18001
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_486
timestamp 18001
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_487
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_488
timestamp 18001
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_489
timestamp 18001
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_490
timestamp 18001
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_491
timestamp 18001
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_492
timestamp 18001
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_493
timestamp 18001
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_494
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_495
timestamp 18001
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_496
timestamp 18001
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_497
timestamp 18001
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_498
timestamp 18001
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_499
timestamp 18001
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_500
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_501
timestamp 18001
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_502
timestamp 18001
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_503
timestamp 18001
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_504
timestamp 18001
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_505
timestamp 18001
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_506
timestamp 18001
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_507
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_508
timestamp 18001
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_509
timestamp 18001
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_510
timestamp 18001
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_511
timestamp 18001
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_512
timestamp 18001
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_513
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_514
timestamp 18001
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_515
timestamp 18001
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_516
timestamp 18001
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_517
timestamp 18001
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_518
timestamp 18001
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_519
timestamp 18001
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_520
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_521
timestamp 18001
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_522
timestamp 18001
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_523
timestamp 18001
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_524
timestamp 18001
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_525
timestamp 18001
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_526
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_527
timestamp 18001
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_528
timestamp 18001
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_529
timestamp 18001
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_530
timestamp 18001
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_531
timestamp 18001
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_532
timestamp 18001
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_533
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_534
timestamp 18001
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_535
timestamp 18001
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_536
timestamp 18001
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_537
timestamp 18001
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_538
timestamp 18001
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_539
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_540
timestamp 18001
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_541
timestamp 18001
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_542
timestamp 18001
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_543
timestamp 18001
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_544
timestamp 18001
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_545
timestamp 18001
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_546
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_547
timestamp 18001
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_548
timestamp 18001
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_549
timestamp 18001
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_550
timestamp 18001
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_551
timestamp 18001
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_552
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_553
timestamp 18001
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_554
timestamp 18001
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_555
timestamp 18001
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_556
timestamp 18001
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_557
timestamp 18001
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_558
timestamp 18001
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_559
timestamp 18001
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_560
timestamp 18001
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_561
timestamp 18001
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_562
timestamp 18001
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_563
timestamp 18001
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_564
timestamp 18001
transform 1 0 34592 0 1 36992
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 cs
port 3 nsew signal input
flabel metal3 s 36782 21088 37582 21208 0 FreeSans 480 0 0 0 dataBusIn[0]
port 4 nsew signal input
flabel metal3 s 36782 21768 37582 21888 0 FreeSans 480 0 0 0 dataBusIn[1]
port 5 nsew signal input
flabel metal3 s 36782 22448 37582 22568 0 FreeSans 480 0 0 0 dataBusIn[2]
port 6 nsew signal input
flabel metal2 s 29642 38926 29698 39726 0 FreeSans 224 90 0 0 dataBusIn[3]
port 7 nsew signal input
flabel metal2 s 28998 38926 29054 39726 0 FreeSans 224 90 0 0 dataBusIn[4]
port 8 nsew signal input
flabel metal3 s 36782 16328 37582 16448 0 FreeSans 480 0 0 0 dataBusIn[5]
port 9 nsew signal input
flabel metal3 s 36782 24488 37582 24608 0 FreeSans 480 0 0 0 dataBusIn[6]
port 10 nsew signal input
flabel metal3 s 36782 23808 37582 23928 0 FreeSans 480 0 0 0 dataBusIn[7]
port 11 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 dataBusOut[0]
port 12 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 dataBusOut[1]
port 13 nsew signal output
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 dataBusOut[2]
port 14 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 dataBusOut[3]
port 15 nsew signal output
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 dataBusOut[4]
port 16 nsew signal output
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 dataBusOut[5]
port 17 nsew signal output
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 dataBusOut[6]
port 18 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 dataBusOut[7]
port 19 nsew signal output
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 dataBusSelect
port 20 nsew signal output
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 gpio[0]
port 21 nsew signal bidirectional
flabel metal2 s 23202 38926 23258 39726 0 FreeSans 224 90 0 0 gpio[10]
port 22 nsew signal bidirectional
flabel metal2 s 25134 38926 25190 39726 0 FreeSans 224 90 0 0 gpio[11]
port 23 nsew signal bidirectional
flabel metal2 s 22558 38926 22614 39726 0 FreeSans 224 90 0 0 gpio[12]
port 24 nsew signal bidirectional
flabel metal2 s 23846 38926 23902 39726 0 FreeSans 224 90 0 0 gpio[13]
port 25 nsew signal bidirectional
flabel metal2 s 25778 38926 25834 39726 0 FreeSans 224 90 0 0 gpio[14]
port 26 nsew signal bidirectional
flabel metal2 s 24490 38926 24546 39726 0 FreeSans 224 90 0 0 gpio[15]
port 27 nsew signal bidirectional
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 gpio[16]
port 28 nsew signal bidirectional
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpio[17]
port 29 nsew signal bidirectional
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 gpio[18]
port 30 nsew signal bidirectional
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 gpio[19]
port 31 nsew signal bidirectional
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 gpio[1]
port 32 nsew signal bidirectional
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 gpio[20]
port 33 nsew signal bidirectional
flabel metal3 s 36782 15648 37582 15768 0 FreeSans 480 0 0 0 gpio[21]
port 34 nsew signal bidirectional
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 gpio[22]
port 35 nsew signal bidirectional
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpio[23]
port 36 nsew signal bidirectional
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 gpio[24]
port 37 nsew signal bidirectional
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 gpio[25]
port 38 nsew signal bidirectional
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 gpio[2]
port 39 nsew signal bidirectional
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 gpio[3]
port 40 nsew signal bidirectional
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 gpio[4]
port 41 nsew signal bidirectional
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 gpio[5]
port 42 nsew signal bidirectional
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 gpio[6]
port 43 nsew signal bidirectional
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 gpio[7]
port 44 nsew signal bidirectional
flabel metal2 s 27066 38926 27122 39726 0 FreeSans 224 90 0 0 gpio[8]
port 45 nsew signal bidirectional
flabel metal2 s 26422 38926 26478 39726 0 FreeSans 224 90 0 0 gpio[9]
port 46 nsew signal bidirectional
flabel metal3 s 36782 3408 37582 3528 0 FreeSans 480 0 0 0 nrst
port 47 nsew signal input
rlabel metal1 18768 36992 18768 36992 0 VGND
rlabel metal1 18768 37536 18768 37536 0 VPWR
rlabel metal1 25852 32878 25852 32878 0 _0000_
rlabel metal2 28290 33694 28290 33694 0 _0001_
rlabel metal2 22402 33388 22402 33388 0 _0002_
rlabel metal2 31418 33252 31418 33252 0 _0003_
rlabel metal1 27646 32980 27646 32980 0 _0004_
rlabel metal2 30406 32640 30406 32640 0 _0005_
rlabel metal2 22770 32980 22770 32980 0 _0006_
rlabel metal1 32246 33082 32246 33082 0 _0007_
rlabel metal1 24702 31416 24702 31416 0 _0008_
rlabel metal1 25898 30158 25898 30158 0 _0009_
rlabel metal2 26358 30226 26358 30226 0 _0010_
rlabel metal2 26634 34408 26634 34408 0 _0011_
rlabel metal1 25576 31654 25576 31654 0 _0012_
rlabel metal1 24886 29070 24886 29070 0 _0013_
rlabel metal1 21390 27098 21390 27098 0 _0014_
rlabel metal2 22586 4284 22586 4284 0 _0015_
rlabel metal1 23368 27642 23368 27642 0 _0016_
rlabel metal1 25300 3570 25300 3570 0 _0017_
rlabel metal1 22540 27030 22540 27030 0 _0018_
rlabel metal1 22402 4046 22402 4046 0 _0019_
rlabel metal1 35650 14042 35650 14042 0 _0020_
rlabel metal2 34592 13396 34592 13396 0 _0021_
rlabel metal1 33718 14042 33718 14042 0 _0022_
rlabel metal1 34500 10710 34500 10710 0 _0023_
rlabel metal1 34178 25806 34178 25806 0 _0024_
rlabel metal2 32338 16796 32338 16796 0 _0025_
rlabel metal1 14444 20366 14444 20366 0 _0026_
rlabel metal1 14536 19754 14536 19754 0 _0027_
rlabel metal1 19964 33490 19964 33490 0 _0028_
rlabel metal1 15640 3094 15640 3094 0 _0029_
rlabel metal2 12834 4250 12834 4250 0 _0030_
rlabel metal1 18216 27098 18216 27098 0 _0031_
rlabel metal1 16238 2890 16238 2890 0 _0032_
rlabel metal1 18078 4726 18078 4726 0 _0033_
rlabel metal1 13202 3400 13202 3400 0 _0034_
rlabel metal1 11408 4794 11408 4794 0 _0035_
rlabel metal1 9338 2822 9338 2822 0 _0036_
rlabel metal2 10902 3740 10902 3740 0 _0037_
rlabel metal1 10994 3128 10994 3128 0 _0038_
rlabel metal1 9476 5270 9476 5270 0 _0039_
rlabel metal1 9844 3910 9844 3910 0 _0040_
rlabel metal1 11868 2482 11868 2482 0 _0041_
rlabel metal1 10488 35802 10488 35802 0 _0042_
rlabel metal1 11316 35802 11316 35802 0 _0043_
rlabel metal2 13294 36516 13294 36516 0 _0044_
rlabel metal2 14398 33150 14398 33150 0 _0045_
rlabel metal1 16192 35802 16192 35802 0 _0046_
rlabel metal1 17894 35734 17894 35734 0 _0047_
rlabel metal1 18768 35734 18768 35734 0 _0048_
rlabel metal1 19090 33898 19090 33898 0 _0049_
rlabel metal1 8832 20502 8832 20502 0 _0050_
rlabel metal2 9798 21284 9798 21284 0 _0051_
rlabel metal1 2024 22202 2024 22202 0 _0052_
rlabel metal1 1840 22746 1840 22746 0 _0053_
rlabel metal2 4094 22814 4094 22814 0 _0054_
rlabel metal1 6440 21862 6440 21862 0 _0055_
rlabel metal2 2162 21284 2162 21284 0 _0056_
rlabel metal1 7169 20026 7169 20026 0 _0057_
rlabel metal1 9154 18394 9154 18394 0 _0058_
rlabel metal2 10258 19618 10258 19618 0 _0059_
rlabel metal1 1886 19482 1886 19482 0 _0060_
rlabel metal1 1886 18394 1886 18394 0 _0061_
rlabel metal1 2231 16014 2231 16014 0 _0062_
rlabel metal1 6026 17306 6026 17306 0 _0063_
rlabel metal1 1840 16762 1840 16762 0 _0064_
rlabel metal2 6762 19108 6762 19108 0 _0065_
rlabel metal1 18814 26894 18814 26894 0 _0066_
rlabel metal2 19918 35054 19918 35054 0 _0067_
rlabel metal1 21436 34986 21436 34986 0 _0068_
rlabel metal2 25254 36822 25254 36822 0 _0069_
rlabel metal1 23000 34170 23000 34170 0 _0070_
rlabel metal2 24426 36516 24426 36516 0 _0071_
rlabel metal2 20194 36652 20194 36652 0 _0072_
rlabel metal2 19642 36516 19642 36516 0 _0073_
rlabel metal1 22678 35768 22678 35768 0 _0074_
rlabel metal1 13800 30090 13800 30090 0 _0075_
rlabel metal1 11362 31926 11362 31926 0 _0076_
rlabel metal2 9062 32096 9062 32096 0 _0077_
rlabel metal1 4416 29818 4416 29818 0 _0078_
rlabel metal2 4416 31994 4416 31994 0 _0079_
rlabel metal1 5198 33626 5198 33626 0 _0080_
rlabel metal2 6762 35428 6762 35428 0 _0081_
rlabel metal1 8004 33082 8004 33082 0 _0082_
rlabel metal2 7590 17374 7590 17374 0 _0083_
rlabel via2 9706 22219 9706 22219 0 _0084_
rlabel metal1 2224 26554 2224 26554 0 _0085_
rlabel metal2 1702 24412 1702 24412 0 _0086_
rlabel metal1 4784 25466 4784 25466 0 _0087_
rlabel metal1 4416 24378 4416 24378 0 _0088_
rlabel metal2 1702 25432 1702 25432 0 _0089_
rlabel metal1 3772 26554 3772 26554 0 _0090_
rlabel metal1 3726 29818 3726 29818 0 _0091_
rlabel metal1 3726 29070 3726 29070 0 _0092_
rlabel metal2 3174 27778 3174 27778 0 _0093_
rlabel metal1 3588 28458 3588 28458 0 _0094_
rlabel metal2 3266 30192 3266 30192 0 _0095_
rlabel metal1 3680 31994 3680 31994 0 _0096_
rlabel metal2 1794 30872 1794 30872 0 _0097_
rlabel metal1 2438 31994 2438 31994 0 _0098_
rlabel metal1 9936 13498 9936 13498 0 _0099_
rlabel metal1 9154 9690 9154 9690 0 _0100_
rlabel metal1 2116 12410 2116 12410 0 _0101_
rlabel metal2 3818 10404 3818 10404 0 _0102_
rlabel metal1 2070 13498 2070 13498 0 _0103_
rlabel metal1 3910 7310 3910 7310 0 _0104_
rlabel metal1 3726 8398 3726 8398 0 _0105_
rlabel metal1 7268 6358 7268 6358 0 _0106_
rlabel metal2 8142 15470 8142 15470 0 _0107_
rlabel metal2 10626 15844 10626 15844 0 _0108_
rlabel metal1 3818 15572 3818 15572 0 _0109_
rlabel metal2 2438 14178 2438 14178 0 _0110_
rlabel metal2 2254 14756 2254 14756 0 _0111_
rlabel metal1 5888 15538 5888 15538 0 _0112_
rlabel metal2 4094 15470 4094 15470 0 _0113_
rlabel metal2 7222 15844 7222 15844 0 _0114_
rlabel metal1 12236 19890 12236 19890 0 _0115_
rlabel metal1 25070 33082 25070 33082 0 _0116_
rlabel metal2 12466 5984 12466 5984 0 _0117_
rlabel metal1 5520 7718 5520 7718 0 _0118_
rlabel viali 5566 10030 5566 10030 0 _0119_
rlabel metal1 5336 9486 5336 9486 0 _0120_
rlabel metal1 3450 16762 3450 16762 0 _0121_
rlabel metal2 4876 18020 4876 18020 0 _0122_
rlabel metal1 4416 17306 4416 17306 0 _0123_
rlabel metal2 5566 19805 5566 19805 0 _0124_
rlabel metal1 6440 27438 6440 27438 0 _0125_
rlabel metal1 5290 26962 5290 26962 0 _0126_
rlabel metal1 8050 25466 8050 25466 0 _0127_
rlabel metal1 15686 22610 15686 22610 0 _0128_
rlabel metal1 14812 22746 14812 22746 0 _0129_
rlabel metal1 14030 24378 14030 24378 0 _0130_
rlabel metal1 6302 25194 6302 25194 0 _0131_
rlabel metal1 5290 27030 5290 27030 0 _0132_
rlabel via2 4278 22933 4278 22933 0 _0133_
rlabel metal1 4462 13328 4462 13328 0 _0134_
rlabel metal1 7130 12818 7130 12818 0 _0135_
rlabel metal1 8556 5542 8556 5542 0 _0136_
rlabel metal1 6394 12614 6394 12614 0 _0137_
rlabel metal1 5060 22746 5060 22746 0 _0138_
rlabel via2 5842 22627 5842 22627 0 _0139_
rlabel metal2 6072 18190 6072 18190 0 _0140_
rlabel metal1 5198 13498 5198 13498 0 _0141_
rlabel metal1 5014 13294 5014 13294 0 _0142_
rlabel metal1 5704 13430 5704 13430 0 _0143_
rlabel metal1 5980 12750 5980 12750 0 _0144_
rlabel metal1 4922 12716 4922 12716 0 _0145_
rlabel metal1 4140 12818 4140 12818 0 _0146_
rlabel metal3 4646 18088 4646 18088 0 _0147_
rlabel metal1 4370 18768 4370 18768 0 _0148_
rlabel metal1 5198 18938 5198 18938 0 _0149_
rlabel metal2 7222 19686 7222 19686 0 _0150_
rlabel metal2 7774 29206 7774 29206 0 _0151_
rlabel metal2 6946 28424 6946 28424 0 _0152_
rlabel metal2 9982 24378 9982 24378 0 _0153_
rlabel metal1 7314 24208 7314 24208 0 _0154_
rlabel metal1 7130 20502 7130 20502 0 _0155_
rlabel metal1 7084 28118 7084 28118 0 _0156_
rlabel metal1 2392 22610 2392 22610 0 _0157_
rlabel metal1 7360 14450 7360 14450 0 _0158_
rlabel metal1 9430 6358 9430 6358 0 _0159_
rlabel metal1 6578 14314 6578 14314 0 _0160_
rlabel via1 5658 23087 5658 23087 0 _0161_
rlabel metal1 6164 23290 6164 23290 0 _0162_
rlabel metal1 5750 29614 5750 29614 0 _0163_
rlabel metal2 2070 13889 2070 13889 0 _0164_
rlabel metal2 5934 13056 5934 13056 0 _0165_
rlabel via1 5014 11118 5014 11118 0 _0166_
rlabel metal2 13018 24922 13018 24922 0 _0167_
rlabel metal2 12282 23936 12282 23936 0 _0168_
rlabel metal2 7498 21301 7498 21301 0 _0169_
rlabel metal1 7728 26962 7728 26962 0 _0170_
rlabel metal1 4462 20400 4462 20400 0 _0171_
rlabel metal2 4554 20604 4554 20604 0 _0172_
rlabel metal1 4646 20026 4646 20026 0 _0173_
rlabel metal1 7498 29614 7498 29614 0 _0174_
rlabel metal1 7544 30226 7544 30226 0 _0175_
rlabel metal2 7314 27676 7314 27676 0 _0176_
rlabel metal2 2714 24225 2714 24225 0 _0177_
rlabel metal1 7452 12818 7452 12818 0 _0178_
rlabel metal1 7820 13226 7820 13226 0 _0179_
rlabel metal1 8786 6630 8786 6630 0 _0180_
rlabel metal1 8418 12852 8418 12852 0 _0181_
rlabel viali 7866 12750 7866 12750 0 _0182_
rlabel metal1 8878 21420 8878 21420 0 _0183_
rlabel metal1 8142 21386 8142 21386 0 _0184_
rlabel metal3 8717 13668 8717 13668 0 _0185_
rlabel metal1 7866 12614 7866 12614 0 _0186_
rlabel metal1 6964 11730 6964 11730 0 _0187_
rlabel metal1 11914 24922 11914 24922 0 _0188_
rlabel metal1 11316 24378 11316 24378 0 _0189_
rlabel metal2 11362 24990 11362 24990 0 _0190_
rlabel metal2 11362 24412 11362 24412 0 _0191_
rlabel metal2 11362 26758 11362 26758 0 _0192_
rlabel metal1 11868 17306 11868 17306 0 _0193_
rlabel metal1 11638 21080 11638 21080 0 _0194_
rlabel metal2 11546 21182 11546 21182 0 _0195_
rlabel metal1 12006 21114 12006 21114 0 _0196_
rlabel metal2 12374 28288 12374 28288 0 _0197_
rlabel metal1 10994 26894 10994 26894 0 _0198_
rlabel metal2 10258 24123 10258 24123 0 _0199_
rlabel metal1 9706 12274 9706 12274 0 _0200_
rlabel metal2 12926 17340 12926 17340 0 _0201_
rlabel metal1 11684 4794 11684 4794 0 _0202_
rlabel metal1 10120 14314 10120 14314 0 _0203_
rlabel metal1 12052 22678 12052 22678 0 _0204_
rlabel via1 11365 23086 11365 23086 0 _0205_
rlabel metal1 12282 22576 12282 22576 0 _0206_
rlabel metal1 10350 29614 10350 29614 0 _0207_
rlabel via2 9982 14467 9982 14467 0 _0208_
rlabel viali 9983 11730 9983 11730 0 _0209_
rlabel metal1 8648 10642 8648 10642 0 _0210_
rlabel metal1 10442 17170 10442 17170 0 _0211_
rlabel metal1 9567 17170 9567 17170 0 _0212_
rlabel metal1 9430 18802 9430 18802 0 _0213_
rlabel via2 9982 17323 9982 17323 0 _0214_
rlabel metal1 10074 28084 10074 28084 0 _0215_
rlabel metal1 13984 27574 13984 27574 0 _0216_
rlabel metal1 13938 27438 13938 27438 0 _0217_
rlabel metal1 13018 27506 13018 27506 0 _0218_
rlabel metal1 10166 28084 10166 28084 0 _0219_
rlabel metal1 11914 25908 11914 25908 0 _0220_
rlabel viali 11822 25806 11822 25806 0 _0221_
rlabel viali 11730 25806 11730 25806 0 _0222_
rlabel metal1 10212 18326 10212 18326 0 _0223_
rlabel metal1 10304 27642 10304 27642 0 _0224_
rlabel metal2 9476 20978 9476 20978 0 _0225_
rlabel metal2 10166 16218 10166 16218 0 _0226_
rlabel metal1 9982 18054 9982 18054 0 _0227_
rlabel metal1 11132 14790 11132 14790 0 _0228_
rlabel metal1 13984 3502 13984 3502 0 _0229_
rlabel metal2 9430 14722 9430 14722 0 _0230_
rlabel metal1 10166 14926 10166 14926 0 _0231_
rlabel metal1 11454 22406 11454 22406 0 _0232_
rlabel metal1 12466 22032 12466 22032 0 _0233_
rlabel metal1 13478 21658 13478 21658 0 _0234_
rlabel metal3 10833 15164 10833 15164 0 _0235_
rlabel metal2 13294 30294 13294 30294 0 _0236_
rlabel metal1 10258 14994 10258 14994 0 _0237_
rlabel metal2 9706 13940 9706 13940 0 _0238_
rlabel metal1 10028 12818 10028 12818 0 _0239_
rlabel metal1 10350 12886 10350 12886 0 _0240_
rlabel metal1 9338 13294 9338 13294 0 _0241_
rlabel via2 15318 17323 15318 17323 0 _0242_
rlabel metal1 16284 15674 16284 15674 0 _0243_
rlabel metal2 15410 17340 15410 17340 0 _0244_
rlabel metal1 16974 8874 16974 8874 0 _0245_
rlabel metal1 17618 9146 17618 9146 0 _0246_
rlabel metal1 16238 17034 16238 17034 0 _0247_
rlabel via1 16154 20502 16154 20502 0 _0248_
rlabel metal2 16330 18700 16330 18700 0 _0249_
rlabel metal1 15134 17136 15134 17136 0 _0250_
rlabel metal1 13386 16116 13386 16116 0 _0251_
rlabel metal1 10488 12818 10488 12818 0 _0252_
rlabel metal1 9476 12614 9476 12614 0 _0253_
rlabel metal1 7958 11696 7958 11696 0 _0254_
rlabel metal1 7084 11118 7084 11118 0 _0255_
rlabel metal1 7452 11730 7452 11730 0 _0256_
rlabel metal2 7406 11390 7406 11390 0 _0257_
rlabel metal2 4830 10914 4830 10914 0 _0258_
rlabel metal2 5290 11424 5290 11424 0 _0259_
rlabel metal1 4554 10982 4554 10982 0 _0260_
rlabel metal1 1978 10098 1978 10098 0 _0261_
rlabel metal1 4094 12172 4094 12172 0 _0262_
rlabel metal2 4692 11084 4692 11084 0 _0263_
rlabel metal1 4830 8806 4830 8806 0 _0264_
rlabel metal1 6624 8466 6624 8466 0 _0265_
rlabel metal2 7314 6868 7314 6868 0 _0266_
rlabel metal1 7636 8058 7636 8058 0 _0267_
rlabel metal2 13294 7174 13294 7174 0 _0268_
rlabel via1 10074 8602 10074 8602 0 _0269_
rlabel metal1 4692 7854 4692 7854 0 _0270_
rlabel metal2 5520 9690 5520 9690 0 _0271_
rlabel via1 6943 9554 6943 9554 0 _0272_
rlabel metal2 5612 12274 5612 12274 0 _0273_
rlabel metal1 7452 8466 7452 8466 0 _0274_
rlabel metal2 7222 7820 7222 7820 0 _0275_
rlabel metal1 1978 11084 1978 11084 0 _0276_
rlabel metal1 1886 9996 1886 9996 0 _0277_
rlabel metal2 3450 9860 3450 9860 0 _0278_
rlabel metal1 4692 10438 4692 10438 0 _0279_
rlabel metal1 2162 9996 2162 9996 0 _0280_
rlabel metal1 3818 8976 3818 8976 0 _0281_
rlabel metal2 2438 12070 2438 12070 0 _0282_
rlabel metal1 5290 8432 5290 8432 0 _0283_
rlabel metal1 6854 7888 6854 7888 0 _0284_
rlabel metal1 6348 6766 6348 6766 0 _0285_
rlabel metal1 6348 6426 6348 6426 0 _0286_
rlabel metal1 4370 7888 4370 7888 0 _0287_
rlabel metal2 4186 6630 4186 6630 0 _0288_
rlabel metal2 5658 5984 5658 5984 0 _0289_
rlabel metal2 6854 6800 6854 6800 0 _0290_
rlabel metal1 4830 6834 4830 6834 0 _0291_
rlabel metal1 5566 7276 5566 7276 0 _0292_
rlabel metal1 5750 6834 5750 6834 0 _0293_
rlabel metal2 8602 7106 8602 7106 0 _0294_
rlabel metal2 13386 18088 13386 18088 0 _0295_
rlabel metal1 12650 9010 12650 9010 0 _0296_
rlabel metal3 15479 18836 15479 18836 0 _0297_
rlabel metal2 12466 6494 12466 6494 0 _0298_
rlabel metal1 12696 8602 12696 8602 0 _0299_
rlabel metal2 12006 8636 12006 8636 0 _0300_
rlabel metal1 12098 8432 12098 8432 0 _0301_
rlabel metal1 19504 9622 19504 9622 0 _0302_
rlabel metal1 19090 13158 19090 13158 0 _0303_
rlabel metal1 13478 5576 13478 5576 0 _0304_
rlabel metal2 11086 6018 11086 6018 0 _0305_
rlabel metal1 11362 6970 11362 6970 0 _0306_
rlabel metal1 10120 5610 10120 5610 0 _0307_
rlabel metal1 10856 5882 10856 5882 0 _0308_
rlabel metal2 13202 6596 13202 6596 0 _0309_
rlabel metal2 13386 7344 13386 7344 0 _0310_
rlabel metal2 14076 18394 14076 18394 0 _0311_
rlabel metal2 11730 9350 11730 9350 0 _0312_
rlabel metal2 18538 10846 18538 10846 0 _0313_
rlabel metal1 11086 9520 11086 9520 0 _0314_
rlabel metal1 8924 7922 8924 7922 0 _0315_
rlabel metal1 9898 7718 9898 7718 0 _0316_
rlabel metal1 10534 7412 10534 7412 0 _0317_
rlabel metal1 11730 7344 11730 7344 0 _0318_
rlabel via1 12374 6171 12374 6171 0 _0319_
rlabel metal1 14628 3638 14628 3638 0 _0320_
rlabel metal2 13570 6664 13570 6664 0 _0321_
rlabel metal1 13064 20910 13064 20910 0 _0322_
rlabel metal2 15686 20570 15686 20570 0 _0323_
rlabel metal1 16468 3026 16468 3026 0 _0324_
rlabel metal2 16422 3604 16422 3604 0 _0325_
rlabel metal1 17940 26962 17940 26962 0 _0326_
rlabel metal2 15962 3876 15962 3876 0 _0327_
rlabel metal2 17158 3468 17158 3468 0 _0328_
rlabel metal1 15840 6358 15840 6358 0 _0329_
rlabel metal2 15502 5882 15502 5882 0 _0330_
rlabel metal2 14766 4624 14766 4624 0 _0331_
rlabel metal1 21022 28730 21022 28730 0 _0332_
rlabel metal1 20562 29172 20562 29172 0 _0333_
rlabel metal2 20562 24157 20562 24157 0 _0334_
rlabel metal1 13570 32402 13570 32402 0 _0335_
rlabel metal1 20332 20434 20332 20434 0 _0336_
rlabel metal1 20194 14858 20194 14858 0 _0337_
rlabel metal2 20378 21012 20378 21012 0 _0338_
rlabel metal1 23138 22746 23138 22746 0 _0339_
rlabel metal1 22494 22610 22494 22610 0 _0340_
rlabel metal2 23414 24038 23414 24038 0 _0341_
rlabel metal1 21712 22066 21712 22066 0 _0342_
rlabel metal2 22586 22814 22586 22814 0 _0343_
rlabel metal1 20378 22508 20378 22508 0 _0344_
rlabel metal2 22862 20604 22862 20604 0 _0345_
rlabel metal1 21712 21862 21712 21862 0 _0346_
rlabel metal1 20332 22406 20332 22406 0 _0347_
rlabel metal1 19826 22746 19826 22746 0 _0348_
rlabel metal1 18676 29274 18676 29274 0 _0349_
rlabel metal1 18814 30260 18814 30260 0 _0350_
rlabel metal1 19182 29614 19182 29614 0 _0351_
rlabel metal1 18308 30226 18308 30226 0 _0352_
rlabel metal1 18998 25874 18998 25874 0 _0353_
rlabel metal1 15042 30226 15042 30226 0 _0354_
rlabel metal2 14122 30498 14122 30498 0 _0355_
rlabel metal1 15318 33490 15318 33490 0 _0356_
rlabel metal1 17020 35054 17020 35054 0 _0357_
rlabel metal1 6946 33524 6946 33524 0 _0358_
rlabel metal2 9614 35836 9614 35836 0 _0359_
rlabel metal2 8970 35972 8970 35972 0 _0360_
rlabel metal1 8878 35258 8878 35258 0 _0361_
rlabel metal2 8602 35258 8602 35258 0 _0362_
rlabel metal2 7866 35700 7866 35700 0 _0363_
rlabel metal2 6026 35700 6026 35700 0 _0364_
rlabel metal2 7130 35530 7130 35530 0 _0365_
rlabel metal2 7314 34816 7314 34816 0 _0366_
rlabel metal1 7774 34612 7774 34612 0 _0367_
rlabel metal2 7222 34170 7222 34170 0 _0368_
rlabel metal1 7452 32538 7452 32538 0 _0369_
rlabel metal1 7866 32436 7866 32436 0 _0370_
rlabel metal1 7130 31382 7130 31382 0 _0371_
rlabel metal1 7406 31246 7406 31246 0 _0372_
rlabel metal1 8418 30736 8418 30736 0 _0373_
rlabel metal1 8096 31314 8096 31314 0 _0374_
rlabel metal1 8234 31790 8234 31790 0 _0375_
rlabel metal1 9430 31280 9430 31280 0 _0376_
rlabel metal2 9798 32045 9798 32045 0 _0377_
rlabel metal2 10074 32436 10074 32436 0 _0378_
rlabel metal1 11960 32198 11960 32198 0 _0379_
rlabel metal1 10074 32912 10074 32912 0 _0380_
rlabel metal2 10350 32606 10350 32606 0 _0381_
rlabel metal1 7590 31858 7590 31858 0 _0382_
rlabel metal1 6578 34102 6578 34102 0 _0383_
rlabel metal1 7268 33830 7268 33830 0 _0384_
rlabel metal2 7038 34748 7038 34748 0 _0385_
rlabel metal2 9338 35700 9338 35700 0 _0386_
rlabel metal1 11316 34986 11316 34986 0 _0387_
rlabel metal1 9706 36074 9706 36074 0 _0388_
rlabel metal2 10166 35836 10166 35836 0 _0389_
rlabel metal2 6946 30396 6946 30396 0 _0390_
rlabel metal2 5842 31518 5842 31518 0 _0391_
rlabel metal1 6624 32810 6624 32810 0 _0392_
rlabel metal1 10028 34034 10028 34034 0 _0393_
rlabel metal1 13846 28458 13846 28458 0 _0394_
rlabel metal1 7866 27948 7866 27948 0 _0395_
rlabel metal2 8878 30124 8878 30124 0 _0396_
rlabel metal1 9476 28186 9476 28186 0 _0397_
rlabel metal1 9752 28730 9752 28730 0 _0398_
rlabel metal1 13846 32844 13846 32844 0 _0399_
rlabel metal1 5106 30634 5106 30634 0 _0400_
rlabel metal1 4708 32810 4708 32810 0 _0401_
rlabel metal2 9706 33252 9706 33252 0 _0402_
rlabel metal2 10258 33524 10258 33524 0 _0403_
rlabel metal2 9522 34102 9522 34102 0 _0404_
rlabel metal2 14950 33762 14950 33762 0 _0405_
rlabel metal2 9890 34374 9890 34374 0 _0406_
rlabel metal1 9890 34714 9890 34714 0 _0407_
rlabel metal2 14030 32708 14030 32708 0 _0408_
rlabel metal2 8096 32878 8096 32878 0 _0409_
rlabel metal2 10902 35462 10902 35462 0 _0410_
rlabel metal1 11730 35190 11730 35190 0 _0411_
rlabel metal2 11638 35258 11638 35258 0 _0412_
rlabel metal1 11638 27982 11638 27982 0 _0413_
rlabel metal1 12190 27370 12190 27370 0 _0414_
rlabel metal1 12466 34000 12466 34000 0 _0415_
rlabel metal1 10856 33490 10856 33490 0 _0416_
rlabel metal1 11500 33626 11500 33626 0 _0417_
rlabel metal1 11684 34170 11684 34170 0 _0418_
rlabel metal2 12006 35428 12006 35428 0 _0419_
rlabel metal2 12926 35394 12926 35394 0 _0420_
rlabel metal1 13708 35462 13708 35462 0 _0421_
rlabel metal1 13754 35054 13754 35054 0 _0422_
rlabel metal2 14306 35054 14306 35054 0 _0423_
rlabel metal1 13892 35258 13892 35258 0 _0424_
rlabel metal1 13708 35802 13708 35802 0 _0425_
rlabel metal1 12788 35802 12788 35802 0 _0426_
rlabel metal1 14582 33456 14582 33456 0 _0427_
rlabel metal1 12696 34170 12696 34170 0 _0428_
rlabel metal2 8142 29818 8142 29818 0 _0429_
rlabel metal2 9384 33626 9384 33626 0 _0430_
rlabel metal2 13846 34323 13846 34323 0 _0431_
rlabel metal1 12696 34714 12696 34714 0 _0432_
rlabel metal1 13110 33966 13110 33966 0 _0433_
rlabel metal2 13110 34204 13110 34204 0 _0434_
rlabel metal2 13846 33660 13846 33660 0 _0435_
rlabel metal1 15548 34102 15548 34102 0 _0436_
rlabel metal1 14214 34034 14214 34034 0 _0437_
rlabel metal1 14950 33524 14950 33524 0 _0438_
rlabel metal2 7222 28662 7222 28662 0 _0439_
rlabel metal1 13110 33422 13110 33422 0 _0440_
rlabel metal2 16330 33728 16330 33728 0 _0441_
rlabel metal2 13386 33371 13386 33371 0 _0442_
rlabel metal1 13616 33490 13616 33490 0 _0443_
rlabel metal1 16054 36788 16054 36788 0 _0444_
rlabel metal1 15594 36686 15594 36686 0 _0445_
rlabel metal1 15272 36754 15272 36754 0 _0446_
rlabel metal2 14306 36380 14306 36380 0 _0447_
rlabel metal1 13478 35088 13478 35088 0 _0448_
rlabel metal2 14122 34578 14122 34578 0 _0449_
rlabel metal2 14214 35700 14214 35700 0 _0450_
rlabel metal1 15272 35666 15272 35666 0 _0451_
rlabel metal1 15962 34170 15962 34170 0 _0452_
rlabel metal2 15318 34816 15318 34816 0 _0453_
rlabel metal1 4968 27642 4968 27642 0 _0454_
rlabel metal2 21390 35479 21390 35479 0 _0455_
rlabel metal2 22586 35955 22586 35955 0 _0456_
rlabel metal1 15318 35122 15318 35122 0 _0457_
rlabel metal1 15364 35258 15364 35258 0 _0458_
rlabel metal1 16698 36822 16698 36822 0 _0459_
rlabel metal2 17526 35666 17526 35666 0 _0460_
rlabel viali 16867 36754 16867 36754 0 _0461_
rlabel metal2 17434 34986 17434 34986 0 _0462_
rlabel metal1 16882 35632 16882 35632 0 _0463_
rlabel metal1 8463 28050 8463 28050 0 _0464_
rlabel via2 9706 27965 9706 27965 0 _0465_
rlabel metal1 17802 34544 17802 34544 0 _0466_
rlabel metal1 15916 34510 15916 34510 0 _0467_
rlabel metal1 14858 35020 14858 35020 0 _0468_
rlabel metal1 17020 34578 17020 34578 0 _0469_
rlabel metal2 16698 35190 16698 35190 0 _0470_
rlabel metal2 17802 36244 17802 36244 0 _0471_
rlabel metal1 17342 36822 17342 36822 0 _0472_
rlabel metal2 17710 35802 17710 35802 0 _0473_
rlabel metal1 18216 35802 18216 35802 0 _0474_
rlabel via2 18078 34595 18078 34595 0 _0475_
rlabel metal2 19274 35360 19274 35360 0 _0476_
rlabel metal1 5951 28526 5951 28526 0 _0477_
rlabel metal2 6302 28713 6302 28713 0 _0478_
rlabel metal1 19458 36108 19458 36108 0 _0479_
rlabel metal1 18630 36346 18630 36346 0 _0480_
rlabel metal2 17158 35258 17158 35258 0 _0481_
rlabel metal1 16974 34034 16974 34034 0 _0482_
rlabel metal1 18078 33932 18078 33932 0 _0483_
rlabel metal2 19182 34068 19182 34068 0 _0484_
rlabel metal2 18998 34170 18998 34170 0 _0485_
rlabel metal1 8970 29648 8970 29648 0 _0486_
rlabel metal1 18170 33490 18170 33490 0 _0487_
rlabel metal1 18216 33626 18216 33626 0 _0488_
rlabel metal1 17940 33966 17940 33966 0 _0489_
rlabel metal1 20010 14416 20010 14416 0 _0490_
rlabel metal1 10488 20978 10488 20978 0 _0491_
rlabel metal1 24380 15538 24380 15538 0 _0492_
rlabel metal2 12098 16252 12098 16252 0 _0493_
rlabel metal2 2622 18734 2622 18734 0 _0494_
rlabel metal2 18170 26758 18170 26758 0 _0495_
rlabel metal1 22067 21930 22067 21930 0 _0496_
rlabel metal1 20654 21862 20654 21862 0 _0497_
rlabel metal1 23874 25806 23874 25806 0 _0498_
rlabel metal1 23276 25398 23276 25398 0 _0499_
rlabel metal1 23506 25976 23506 25976 0 _0500_
rlabel viali 20666 25874 20666 25874 0 _0501_
rlabel metal1 20286 26010 20286 26010 0 _0502_
rlabel metal2 20562 31484 20562 31484 0 _0503_
rlabel metal2 20194 31042 20194 31042 0 _0504_
rlabel metal1 19412 31246 19412 31246 0 _0505_
rlabel metal2 21114 33524 21114 33524 0 _0506_
rlabel metal2 13202 30362 13202 30362 0 _0507_
rlabel metal1 10626 29818 10626 29818 0 _0508_
rlabel metal2 10902 30464 10902 30464 0 _0509_
rlabel metal1 11546 30362 11546 30362 0 _0510_
rlabel metal1 11086 30838 11086 30838 0 _0511_
rlabel metal1 11546 31450 11546 31450 0 _0512_
rlabel metal2 11454 31994 11454 31994 0 _0513_
rlabel metal1 9844 30770 9844 30770 0 _0514_
rlabel metal1 9752 30838 9752 30838 0 _0515_
rlabel metal1 10166 32844 10166 32844 0 _0516_
rlabel metal1 9844 31994 9844 31994 0 _0517_
rlabel metal1 9430 31450 9430 31450 0 _0518_
rlabel metal2 5842 30634 5842 30634 0 _0519_
rlabel metal1 8050 31178 8050 31178 0 _0520_
rlabel metal1 6026 30634 6026 30634 0 _0521_
rlabel metal1 6072 30362 6072 30362 0 _0522_
rlabel metal1 5428 29614 5428 29614 0 _0523_
rlabel metal1 7498 32198 7498 32198 0 _0524_
rlabel metal1 6808 31926 6808 31926 0 _0525_
rlabel metal2 5106 32028 5106 32028 0 _0526_
rlabel metal1 5014 31348 5014 31348 0 _0527_
rlabel metal1 4554 30770 4554 30770 0 _0528_
rlabel metal1 4600 30906 4600 30906 0 _0529_
rlabel metal1 5152 31450 5152 31450 0 _0530_
rlabel metal1 6808 31450 6808 31450 0 _0531_
rlabel metal1 5244 32946 5244 32946 0 _0532_
rlabel metal2 5290 33218 5290 33218 0 _0533_
rlabel metal2 5566 33252 5566 33252 0 _0534_
rlabel metal1 7268 32878 7268 32878 0 _0535_
rlabel metal2 7314 33218 7314 33218 0 _0536_
rlabel metal1 6900 34578 6900 34578 0 _0537_
rlabel metal1 6532 34714 6532 34714 0 _0538_
rlabel metal1 6118 32402 6118 32402 0 _0539_
rlabel metal2 6670 33694 6670 33694 0 _0540_
rlabel metal1 6578 33456 6578 33456 0 _0541_
rlabel metal2 6762 32640 6762 32640 0 _0542_
rlabel metal1 6302 33626 6302 33626 0 _0543_
rlabel metal2 6118 34884 6118 34884 0 _0544_
rlabel metal1 8326 35020 8326 35020 0 _0545_
rlabel metal1 8326 32912 8326 32912 0 _0546_
rlabel metal2 8142 33796 8142 33796 0 _0547_
rlabel metal1 8372 33898 8372 33898 0 _0548_
rlabel metal2 8418 33490 8418 33490 0 _0549_
rlabel metal2 21390 17476 21390 17476 0 _0550_
rlabel metal1 21114 17646 21114 17646 0 _0551_
rlabel via2 5474 24259 5474 24259 0 _0552_
rlabel metal1 21482 25228 21482 25228 0 _0553_
rlabel metal2 21758 25466 21758 25466 0 _0554_
rlabel metal1 23322 24718 23322 24718 0 _0555_
rlabel metal2 22770 25092 22770 25092 0 _0556_
rlabel metal1 20608 25194 20608 25194 0 _0557_
rlabel metal1 19734 25466 19734 25466 0 _0558_
rlabel metal2 19366 30430 19366 30430 0 _0559_
rlabel metal1 2346 31280 2346 31280 0 _0560_
rlabel metal1 10810 13328 10810 13328 0 _0561_
rlabel metal1 10350 13294 10350 13294 0 _0562_
rlabel metal1 6440 9962 6440 9962 0 _0563_
rlabel metal1 6164 12682 6164 12682 0 _0564_
rlabel metal2 12098 10370 12098 10370 0 _0565_
rlabel metal2 26726 8823 26726 8823 0 _0566_
rlabel metal2 10948 11118 10948 11118 0 _0567_
rlabel metal1 10488 12410 10488 12410 0 _0568_
rlabel metal2 10074 12002 10074 12002 0 _0569_
rlabel metal1 9936 12206 9936 12206 0 _0570_
rlabel metal1 10350 12342 10350 12342 0 _0571_
rlabel metal1 16652 12206 16652 12206 0 _0572_
rlabel metal1 13754 12206 13754 12206 0 _0573_
rlabel metal2 12926 11798 12926 11798 0 _0574_
rlabel metal1 12282 11662 12282 11662 0 _0575_
rlabel metal2 10350 13090 10350 13090 0 _0576_
rlabel metal1 2208 10098 2208 10098 0 _0577_
rlabel metal1 9108 9418 9108 9418 0 _0578_
rlabel metal1 8694 11696 8694 11696 0 _0579_
rlabel metal2 8970 11084 8970 11084 0 _0580_
rlabel metal2 8878 11118 8878 11118 0 _0581_
rlabel metal2 9522 10540 9522 10540 0 _0582_
rlabel metal1 9706 9554 9706 9554 0 _0583_
rlabel metal1 3404 9894 3404 9894 0 _0584_
rlabel metal1 9430 9588 9430 9588 0 _0585_
rlabel metal2 2346 10030 2346 10030 0 _0586_
rlabel metal2 2714 10370 2714 10370 0 _0587_
rlabel metal1 2208 10234 2208 10234 0 _0588_
rlabel metal1 2254 11118 2254 11118 0 _0589_
rlabel metal1 6486 11594 6486 11594 0 _0590_
rlabel metal1 6348 12274 6348 12274 0 _0591_
rlabel metal1 6532 11866 6532 11866 0 _0592_
rlabel metal1 3082 11764 3082 11764 0 _0593_
rlabel metal1 3082 11866 3082 11866 0 _0594_
rlabel metal2 2898 11730 2898 11730 0 _0595_
rlabel metal2 3726 10846 3726 10846 0 _0596_
rlabel metal2 4140 10030 4140 10030 0 _0597_
rlabel metal1 4094 10064 4094 10064 0 _0598_
rlabel metal2 4922 11322 4922 11322 0 _0599_
rlabel metal1 5290 10676 5290 10676 0 _0600_
rlabel metal2 4002 10234 4002 10234 0 _0601_
rlabel metal1 3910 12274 3910 12274 0 _0602_
rlabel metal1 5371 12818 5371 12818 0 _0603_
rlabel metal2 4278 12342 4278 12342 0 _0604_
rlabel metal1 3726 12410 3726 12410 0 _0605_
rlabel metal1 3266 12172 3266 12172 0 _0606_
rlabel metal2 3266 13090 3266 13090 0 _0607_
rlabel metal1 6026 9486 6026 9486 0 _0608_
rlabel metal1 5888 9350 5888 9350 0 _0609_
rlabel metal2 5198 9146 5198 9146 0 _0610_
rlabel metal2 4830 9146 4830 9146 0 _0611_
rlabel metal2 4830 8330 4830 8330 0 _0612_
rlabel metal1 4140 6834 4140 6834 0 _0613_
rlabel metal1 4462 6834 4462 6834 0 _0614_
rlabel metal2 4370 6596 4370 6596 0 _0615_
rlabel metal1 4600 6970 4600 6970 0 _0616_
rlabel metal1 6394 8330 6394 8330 0 _0617_
rlabel metal2 6394 8704 6394 8704 0 _0618_
rlabel metal2 6670 9146 6670 9146 0 _0619_
rlabel metal2 6762 9146 6762 9146 0 _0620_
rlabel metal1 5980 8942 5980 8942 0 _0621_
rlabel metal1 5152 8534 5152 8534 0 _0622_
rlabel metal1 5980 7242 5980 7242 0 _0623_
rlabel metal2 5382 6596 5382 6596 0 _0624_
rlabel metal2 5290 6052 5290 6052 0 _0625_
rlabel metal1 5198 6426 5198 6426 0 _0626_
rlabel metal1 5244 7514 5244 7514 0 _0627_
rlabel metal1 9752 7990 9752 7990 0 _0628_
rlabel metal1 9062 7514 9062 7514 0 _0629_
rlabel metal1 9154 8976 9154 8976 0 _0630_
rlabel metal2 8970 9418 8970 9418 0 _0631_
rlabel metal1 9292 8466 9292 8466 0 _0632_
rlabel metal2 8878 7854 8878 7854 0 _0633_
rlabel viali 7126 6766 7126 6766 0 _0634_
rlabel metal1 6348 6834 6348 6834 0 _0635_
rlabel metal1 22724 13906 22724 13906 0 _0636_
rlabel metal2 12558 15164 12558 15164 0 _0637_
rlabel metal1 12788 19142 12788 19142 0 _0638_
rlabel viali 25162 32950 25162 32950 0 _0639_
rlabel metal1 13110 6290 13110 6290 0 _0640_
rlabel metal1 23552 11050 23552 11050 0 _0641_
rlabel metal1 28428 10166 28428 10166 0 _0642_
rlabel metal1 19182 15130 19182 15130 0 _0643_
rlabel metal2 19366 32572 19366 32572 0 _0644_
rlabel metal1 12926 5032 12926 5032 0 _0645_
rlabel metal1 13708 6426 13708 6426 0 _0646_
rlabel metal2 9154 22984 9154 22984 0 _0647_
rlabel metal2 13018 20145 13018 20145 0 _0648_
rlabel metal1 15364 4454 15364 4454 0 _0649_
rlabel metal2 26634 32844 26634 32844 0 _0650_
rlabel metal1 26634 29614 26634 29614 0 _0651_
rlabel metal1 25760 32538 25760 32538 0 _0652_
rlabel metal1 22448 2482 22448 2482 0 _0653_
rlabel metal1 31234 16048 31234 16048 0 _0654_
rlabel metal1 28106 7786 28106 7786 0 _0655_
rlabel metal2 22034 24990 22034 24990 0 _0656_
rlabel metal1 27646 12614 27646 12614 0 _0657_
rlabel metal2 27922 7616 27922 7616 0 _0658_
rlabel metal2 20010 6205 20010 6205 0 _0659_
rlabel metal1 31832 10506 31832 10506 0 _0660_
rlabel metal1 21390 5712 21390 5712 0 _0661_
rlabel metal1 27508 5542 27508 5542 0 _0662_
rlabel metal2 21390 18734 21390 18734 0 _0663_
rlabel metal1 22954 11084 22954 11084 0 _0664_
rlabel metal1 18124 13294 18124 13294 0 _0665_
rlabel via2 34454 10251 34454 10251 0 _0666_
rlabel metal1 24886 25908 24886 25908 0 _0667_
rlabel metal1 32798 9146 32798 9146 0 _0668_
rlabel metal2 27462 3842 27462 3842 0 _0669_
rlabel metal1 15318 15028 15318 15028 0 _0670_
rlabel metal2 24702 15810 24702 15810 0 _0671_
rlabel metal3 34339 20740 34339 20740 0 _0672_
rlabel metal1 14858 7922 14858 7922 0 _0673_
rlabel metal2 20838 9503 20838 9503 0 _0674_
rlabel metal1 26266 20944 26266 20944 0 _0675_
rlabel metal2 23046 19839 23046 19839 0 _0676_
rlabel metal2 19274 32606 19274 32606 0 _0677_
rlabel metal1 19504 21318 19504 21318 0 _0678_
rlabel metal1 20378 32198 20378 32198 0 _0679_
rlabel metal1 19274 19380 19274 19380 0 _0680_
rlabel via2 20286 26469 20286 26469 0 _0681_
rlabel metal2 29302 16830 29302 16830 0 _0682_
rlabel metal2 32890 7922 32890 7922 0 _0683_
rlabel metal2 19044 15028 19044 15028 0 _0684_
rlabel metal1 31050 13158 31050 13158 0 _0685_
rlabel metal2 30682 7480 30682 7480 0 _0686_
rlabel metal1 24104 18258 24104 18258 0 _0687_
rlabel metal1 33442 9520 33442 9520 0 _0688_
rlabel metal1 33534 9622 33534 9622 0 _0689_
rlabel via1 34845 12206 34845 12206 0 _0690_
rlabel metal1 29923 8330 29923 8330 0 _0691_
rlabel metal1 24748 6426 24748 6426 0 _0692_
rlabel metal2 29854 8262 29854 8262 0 _0693_
rlabel metal1 34178 16218 34178 16218 0 _0694_
rlabel metal2 32338 7361 32338 7361 0 _0695_
rlabel metal2 10626 11577 10626 11577 0 _0696_
rlabel metal2 17802 9010 17802 9010 0 _0697_
rlabel metal2 21574 8500 21574 8500 0 _0698_
rlabel metal1 23000 17510 23000 17510 0 _0699_
rlabel metal2 32982 11849 32982 11849 0 _0700_
rlabel metal2 25714 7650 25714 7650 0 _0701_
rlabel via2 32154 15147 32154 15147 0 _0702_
rlabel metal2 20562 7616 20562 7616 0 _0703_
rlabel metal2 21390 28577 21390 28577 0 _0704_
rlabel metal2 21574 6018 21574 6018 0 _0705_
rlabel metal1 28658 8942 28658 8942 0 _0706_
rlabel via2 31234 10251 31234 10251 0 _0707_
rlabel metal2 24978 7616 24978 7616 0 _0708_
rlabel metal2 23046 7548 23046 7548 0 _0709_
rlabel metal1 23138 7412 23138 7412 0 _0710_
rlabel metal1 22632 2414 22632 2414 0 _0711_
rlabel metal1 16928 18938 16928 18938 0 _0712_
rlabel metal1 19090 24378 19090 24378 0 _0713_
rlabel metal3 19872 18972 19872 18972 0 _0714_
rlabel metal1 21114 3706 21114 3706 0 _0715_
rlabel metal2 14306 21495 14306 21495 0 _0716_
rlabel metal1 32798 12818 32798 12818 0 _0717_
rlabel metal1 32890 9962 32890 9962 0 _0718_
rlabel metal2 28750 10812 28750 10812 0 _0719_
rlabel metal4 19228 25908 19228 25908 0 _0720_
rlabel metal1 31372 11254 31372 11254 0 _0721_
rlabel metal2 29026 10812 29026 10812 0 _0722_
rlabel via1 29946 6851 29946 6851 0 _0723_
rlabel metal1 20562 15470 20562 15470 0 _0724_
rlabel metal1 27278 6426 27278 6426 0 _0725_
rlabel metal1 27094 3638 27094 3638 0 _0726_
rlabel metal1 27738 6324 27738 6324 0 _0727_
rlabel metal1 26956 3502 26956 3502 0 _0728_
rlabel metal1 27002 3366 27002 3366 0 _0729_
rlabel metal2 27370 6460 27370 6460 0 _0730_
rlabel metal1 27048 3434 27048 3434 0 _0731_
rlabel metal1 20654 15062 20654 15062 0 _0732_
rlabel metal2 21114 3553 21114 3553 0 _0733_
rlabel metal1 20148 15470 20148 15470 0 _0734_
rlabel metal1 13524 19142 13524 19142 0 _0735_
rlabel metal1 19274 15538 19274 15538 0 _0736_
rlabel metal1 20976 15674 20976 15674 0 _0737_
rlabel metal1 20194 8908 20194 8908 0 _0738_
rlabel metal2 32982 18207 32982 18207 0 _0739_
rlabel metal1 21344 23290 21344 23290 0 _0740_
rlabel metal3 21827 22508 21827 22508 0 _0741_
rlabel metal1 21942 12920 21942 12920 0 _0742_
rlabel metal2 21666 7259 21666 7259 0 _0743_
rlabel metal1 25714 24378 25714 24378 0 _0744_
rlabel metal1 21114 9996 21114 9996 0 _0745_
rlabel metal2 20102 7038 20102 7038 0 _0746_
rlabel metal2 22678 9690 22678 9690 0 _0747_
rlabel metal2 21068 13396 21068 13396 0 _0748_
rlabel metal1 21206 12614 21206 12614 0 _0749_
rlabel metal1 18814 17850 18814 17850 0 _0750_
rlabel metal1 31694 17136 31694 17136 0 _0751_
rlabel metal2 23230 12529 23230 12529 0 _0752_
rlabel metal2 21206 11050 21206 11050 0 _0753_
rlabel metal1 21988 12818 21988 12818 0 _0754_
rlabel metal2 21390 20162 21390 20162 0 _0755_
rlabel metal1 28980 15334 28980 15334 0 _0756_
rlabel metal1 17296 9418 17296 9418 0 _0757_
rlabel metal1 23414 20774 23414 20774 0 _0758_
rlabel metal1 21850 13940 21850 13940 0 _0759_
rlabel metal1 21850 20298 21850 20298 0 _0760_
rlabel metal1 21390 20298 21390 20298 0 _0761_
rlabel metal1 21712 20502 21712 20502 0 _0762_
rlabel metal1 22264 20570 22264 20570 0 _0763_
rlabel metal1 22448 20774 22448 20774 0 _0764_
rlabel metal2 27646 17119 27646 17119 0 _0765_
rlabel via2 26266 21981 26266 21981 0 _0766_
rlabel metal1 26082 16762 26082 16762 0 _0767_
rlabel metal2 25254 15504 25254 15504 0 _0768_
rlabel metal2 32292 16524 32292 16524 0 _0769_
rlabel metal1 25070 16592 25070 16592 0 _0770_
rlabel metal1 21758 8330 21758 8330 0 _0771_
rlabel metal1 25162 16116 25162 16116 0 _0772_
rlabel via2 22218 15997 22218 15997 0 _0773_
rlabel metal1 17986 10506 17986 10506 0 _0774_
rlabel metal1 17342 11254 17342 11254 0 _0775_
rlabel metal1 32522 25704 32522 25704 0 _0776_
rlabel metal1 26082 14416 26082 14416 0 _0777_
rlabel metal2 27508 14484 27508 14484 0 _0778_
rlabel metal2 28014 20825 28014 20825 0 _0779_
rlabel metal1 25484 18734 25484 18734 0 _0780_
rlabel metal1 26358 18802 26358 18802 0 _0781_
rlabel metal1 28106 19720 28106 19720 0 _0782_
rlabel metal2 25438 23103 25438 23103 0 _0783_
rlabel metal2 25438 16286 25438 16286 0 _0784_
rlabel metal1 24886 14586 24886 14586 0 _0785_
rlabel metal1 20056 19346 20056 19346 0 _0786_
rlabel metal2 17434 16320 17434 16320 0 _0787_
rlabel metal1 21804 12818 21804 12818 0 _0788_
rlabel metal1 25806 8058 25806 8058 0 _0789_
rlabel metal1 26128 16150 26128 16150 0 _0790_
rlabel metal2 25898 18445 25898 18445 0 _0791_
rlabel metal2 19182 14586 19182 14586 0 _0792_
rlabel metal1 18216 10166 18216 10166 0 _0793_
rlabel metal2 17526 11169 17526 11169 0 _0794_
rlabel metal2 25898 9248 25898 9248 0 _0795_
rlabel metal1 27646 18938 27646 18938 0 _0796_
rlabel metal1 27048 9418 27048 9418 0 _0797_
rlabel metal2 22310 14518 22310 14518 0 _0798_
rlabel metal2 25990 15776 25990 15776 0 _0799_
rlabel metal1 25760 14042 25760 14042 0 _0800_
rlabel metal1 26220 14586 26220 14586 0 _0801_
rlabel metal1 22540 16116 22540 16116 0 _0802_
rlabel metal2 18354 29954 18354 29954 0 _0803_
rlabel metal1 32062 29716 32062 29716 0 _0804_
rlabel metal1 17802 31960 17802 31960 0 _0805_
rlabel metal1 18998 30736 18998 30736 0 _0806_
rlabel metal1 21022 31178 21022 31178 0 _0807_
rlabel metal1 16836 19754 16836 19754 0 _0808_
rlabel metal1 15364 16082 15364 16082 0 _0809_
rlabel metal2 22678 28934 22678 28934 0 _0810_
rlabel metal1 17940 32538 17940 32538 0 _0811_
rlabel via3 15755 19244 15755 19244 0 _0812_
rlabel metal1 22448 30022 22448 30022 0 _0813_
rlabel metal1 16468 32470 16468 32470 0 _0814_
rlabel metal1 22494 30770 22494 30770 0 _0815_
rlabel metal1 15962 32266 15962 32266 0 _0816_
rlabel via3 22885 6868 22885 6868 0 _0817_
rlabel metal1 22586 29070 22586 29070 0 _0818_
rlabel metal1 23414 28662 23414 28662 0 _0819_
rlabel metal1 20792 26962 20792 26962 0 _0820_
rlabel metal1 24886 24922 24886 24922 0 _0821_
rlabel metal2 32062 26554 32062 26554 0 _0822_
rlabel metal1 26266 28186 26266 28186 0 _0823_
rlabel via2 18446 4267 18446 4267 0 _0824_
rlabel metal3 22632 28764 22632 28764 0 _0825_
rlabel metal1 31786 28424 31786 28424 0 _0826_
rlabel metal1 29394 23630 29394 23630 0 _0827_
rlabel metal1 29532 31994 29532 31994 0 _0828_
rlabel metal1 27922 30906 27922 30906 0 _0829_
rlabel via1 27904 26350 27904 26350 0 _0830_
rlabel metal1 29118 30770 29118 30770 0 _0831_
rlabel metal1 31326 32334 31326 32334 0 _0832_
rlabel metal1 27554 30226 27554 30226 0 _0833_
rlabel metal2 26910 29818 26910 29818 0 _0834_
rlabel metal2 27554 27200 27554 27200 0 _0835_
rlabel metal1 32246 26520 32246 26520 0 _0836_
rlabel metal1 32292 32810 32292 32810 0 _0837_
rlabel metal1 31824 31382 31824 31382 0 _0838_
rlabel metal1 32246 31722 32246 31722 0 _0839_
rlabel metal1 32292 31994 32292 31994 0 _0840_
rlabel metal1 32016 32538 32016 32538 0 _0841_
rlabel metal1 33258 32300 33258 32300 0 _0842_
rlabel via1 32622 31654 32622 31654 0 _0843_
rlabel metal2 30406 32079 30406 32079 0 _0844_
rlabel metal2 32798 32164 32798 32164 0 _0845_
rlabel metal1 33028 32402 33028 32402 0 _0846_
rlabel metal2 33442 32708 33442 32708 0 _0847_
rlabel metal2 28934 29750 28934 29750 0 _0848_
rlabel metal1 27830 32538 27830 32538 0 _0849_
rlabel via1 32325 14994 32325 14994 0 _0850_
rlabel metal2 27922 30940 27922 30940 0 _0851_
rlabel via1 27462 31773 27462 31773 0 _0852_
rlabel metal2 30176 19380 30176 19380 0 _0853_
rlabel metal1 25622 31382 25622 31382 0 _0854_
rlabel metal1 27600 30838 27600 30838 0 _0855_
rlabel metal1 26910 30804 26910 30804 0 _0856_
rlabel metal1 22908 32402 22908 32402 0 _0857_
rlabel metal1 21620 32538 21620 32538 0 _0858_
rlabel metal1 29992 30702 29992 30702 0 _0859_
rlabel metal1 29992 31994 29992 31994 0 _0860_
rlabel metal2 29578 30396 29578 30396 0 _0861_
rlabel metal2 29670 29036 29670 29036 0 _0862_
rlabel metal2 32062 11373 32062 11373 0 _0863_
rlabel metal1 26680 31790 26680 31790 0 _0864_
rlabel metal1 27922 31790 27922 31790 0 _0865_
rlabel metal2 25714 19278 25714 19278 0 _0866_
rlabel metal1 29532 32198 29532 32198 0 _0867_
rlabel metal1 30590 32300 30590 32300 0 _0868_
rlabel metal2 28842 32334 28842 32334 0 _0869_
rlabel metal1 26450 31450 26450 31450 0 _0870_
rlabel metal1 28566 32334 28566 32334 0 _0871_
rlabel metal1 28290 31994 28290 31994 0 _0872_
rlabel metal1 26082 31790 26082 31790 0 _0873_
rlabel metal2 33350 29563 33350 29563 0 _0874_
rlabel metal2 33166 29036 33166 29036 0 _0875_
rlabel metal1 27094 26316 27094 26316 0 _0876_
rlabel metal1 27554 26316 27554 26316 0 _0877_
rlabel via1 29670 18734 29670 18734 0 _0878_
rlabel metal1 29716 26010 29716 26010 0 _0879_
rlabel viali 33810 25877 33810 25877 0 _0880_
rlabel metal1 28796 17238 28796 17238 0 _0881_
rlabel metal1 35374 24718 35374 24718 0 _0882_
rlabel metal1 32246 22576 32246 22576 0 _0883_
rlabel viali 34638 26962 34638 26962 0 _0884_
rlabel metal1 35236 24786 35236 24786 0 _0885_
rlabel metal1 35742 24582 35742 24582 0 _0886_
rlabel metal1 31878 20910 31878 20910 0 _0887_
rlabel metal1 28382 24378 28382 24378 0 _0888_
rlabel metal2 33718 18496 33718 18496 0 _0889_
rlabel metal1 28152 24752 28152 24752 0 _0890_
rlabel metal1 31970 24582 31970 24582 0 _0891_
rlabel metal1 25714 26384 25714 26384 0 _0892_
rlabel metal1 26082 20434 26082 20434 0 _0893_
rlabel metal2 26634 24582 26634 24582 0 _0894_
rlabel metal2 27462 27591 27462 27591 0 _0895_
rlabel metal1 26266 27404 26266 27404 0 _0896_
rlabel metal2 32982 19380 32982 19380 0 _0897_
rlabel metal2 25990 25772 25990 25772 0 _0898_
rlabel metal2 28750 24633 28750 24633 0 _0899_
rlabel metal1 34730 23732 34730 23732 0 _0900_
rlabel metal1 27554 23834 27554 23834 0 _0901_
rlabel metal1 32798 23664 32798 23664 0 _0902_
rlabel metal1 28290 22610 28290 22610 0 _0903_
rlabel via1 27646 18734 27646 18734 0 _0904_
rlabel metal1 28842 23290 28842 23290 0 _0905_
rlabel metal1 33994 23494 33994 23494 0 _0906_
rlabel metal1 32798 28016 32798 28016 0 _0907_
rlabel metal1 34638 16116 34638 16116 0 _0908_
rlabel viali 32705 18258 32705 18258 0 _0909_
rlabel metal2 33074 20740 33074 20740 0 _0910_
rlabel metal1 32062 28050 32062 28050 0 _0911_
rlabel metal2 31878 27642 31878 27642 0 _0912_
rlabel viali 27462 28523 27462 28523 0 _0913_
rlabel metal2 29578 28934 29578 28934 0 _0914_
rlabel metal1 32476 28594 32476 28594 0 _0915_
rlabel metal2 31694 28016 31694 28016 0 _0916_
rlabel metal1 28658 27982 28658 27982 0 _0917_
rlabel metal2 27278 28050 27278 28050 0 _0918_
rlabel metal1 28290 28186 28290 28186 0 _0919_
rlabel metal1 31694 27404 31694 27404 0 _0920_
rlabel metal2 33534 26486 33534 26486 0 _0921_
rlabel metal1 31970 14994 31970 14994 0 _0922_
rlabel metal1 30866 15674 30866 15674 0 _0923_
rlabel metal1 32384 15606 32384 15606 0 _0924_
rlabel metal1 35512 18258 35512 18258 0 _0925_
rlabel metal1 27002 20502 27002 20502 0 _0926_
rlabel metal1 28060 20502 28060 20502 0 _0927_
rlabel metal1 28014 20434 28014 20434 0 _0928_
rlabel metal2 29578 20128 29578 20128 0 _0929_
rlabel metal1 27646 20400 27646 20400 0 _0930_
rlabel metal1 27784 14042 27784 14042 0 _0931_
rlabel metal2 27462 14688 27462 14688 0 _0932_
rlabel metal1 30406 17612 30406 17612 0 _0933_
rlabel metal2 34086 14586 34086 14586 0 _0934_
rlabel metal1 30084 16966 30084 16966 0 _0935_
rlabel metal1 32062 14586 32062 14586 0 _0936_
rlabel metal2 33074 30668 33074 30668 0 _0937_
rlabel via2 32522 13379 32522 13379 0 _0938_
rlabel metal1 33718 14450 33718 14450 0 _0939_
rlabel metal1 34224 14314 34224 14314 0 _0940_
rlabel metal1 34638 14246 34638 14246 0 _0941_
rlabel metal1 34270 17612 34270 17612 0 _0942_
rlabel metal1 27324 18258 27324 18258 0 _0943_
rlabel metal1 27876 18394 27876 18394 0 _0944_
rlabel metal1 28566 18598 28566 18598 0 _0945_
rlabel metal1 29302 13498 29302 13498 0 _0946_
rlabel metal1 33764 13702 33764 13702 0 _0947_
rlabel metal1 34868 15674 34868 15674 0 _0948_
rlabel metal1 35420 19890 35420 19890 0 _0949_
rlabel metal2 33350 14110 33350 14110 0 _0950_
rlabel metal1 35420 13906 35420 13906 0 _0951_
rlabel metal2 32798 15402 32798 15402 0 _0952_
rlabel metal1 33212 13498 33212 13498 0 _0953_
rlabel metal1 31050 24038 31050 24038 0 _0954_
rlabel metal2 32522 15606 32522 15606 0 _0955_
rlabel metal2 33350 18428 33350 18428 0 _0956_
rlabel metal1 34086 18360 34086 18360 0 _0957_
rlabel metal2 32798 17187 32798 17187 0 _0958_
rlabel metal1 33534 18122 33534 18122 0 _0959_
rlabel metal1 35190 18734 35190 18734 0 _0960_
rlabel metal2 31878 23222 31878 23222 0 _0961_
rlabel metal1 33442 22644 33442 22644 0 _0962_
rlabel metal1 33534 22440 33534 22440 0 _0963_
rlabel metal2 32798 23052 32798 23052 0 _0964_
rlabel metal1 33810 20026 33810 20026 0 _0965_
rlabel metal3 31073 23732 31073 23732 0 _0966_
rlabel metal1 32062 13906 32062 13906 0 _0967_
rlabel metal1 30038 17714 30038 17714 0 _0968_
rlabel metal2 32890 19040 32890 19040 0 _0969_
rlabel metal1 33074 14042 33074 14042 0 _0970_
rlabel metal2 35374 18462 35374 18462 0 _0971_
rlabel metal2 30038 20502 30038 20502 0 _0972_
rlabel metal1 30636 20434 30636 20434 0 _0973_
rlabel metal2 31326 20604 31326 20604 0 _0974_
rlabel metal1 30406 27914 30406 27914 0 _0975_
rlabel metal1 30084 27506 30084 27506 0 _0976_
rlabel metal2 32798 20230 32798 20230 0 _0977_
rlabel metal2 28842 20774 28842 20774 0 _0978_
rlabel metal1 28704 21590 28704 21590 0 _0979_
rlabel metal1 31326 20230 31326 20230 0 _0980_
rlabel metal2 33994 20060 33994 20060 0 _0981_
rlabel metal1 33948 19754 33948 19754 0 _0982_
rlabel metal1 34132 13906 34132 13906 0 _0983_
rlabel metal2 30314 19635 30314 19635 0 _0984_
rlabel metal1 32016 17306 32016 17306 0 _0985_
rlabel metal1 33212 11322 33212 11322 0 _0986_
rlabel metal2 34638 23052 34638 23052 0 _0987_
rlabel metal1 34822 15538 34822 15538 0 _0988_
rlabel metal1 35006 21998 35006 21998 0 _0989_
rlabel metal1 34914 21862 34914 21862 0 _0990_
rlabel metal1 33810 15402 33810 15402 0 _0991_
rlabel metal2 32430 25976 32430 25976 0 _0992_
rlabel metal2 34546 19040 34546 19040 0 _0993_
rlabel metal2 34638 20570 34638 20570 0 _0994_
rlabel metal2 28566 19448 28566 19448 0 _0995_
rlabel metal1 30728 20026 30728 20026 0 _0996_
rlabel metal1 34454 20570 34454 20570 0 _0997_
rlabel metal1 33258 25398 33258 25398 0 _0998_
rlabel metal2 33350 25670 33350 25670 0 _0999_
rlabel metal2 31786 25466 31786 25466 0 _1000_
rlabel metal2 32154 26214 32154 26214 0 _1001_
rlabel metal2 28014 27914 28014 27914 0 _1002_
rlabel metal2 27738 25500 27738 25500 0 _1003_
rlabel metal1 29946 26282 29946 26282 0 _1004_
rlabel via2 32269 25092 32269 25092 0 _1005_
rlabel metal1 32798 20298 32798 20298 0 _1006_
rlabel metal2 34730 16354 34730 16354 0 _1007_
rlabel metal2 30314 17374 30314 17374 0 _1008_
rlabel metal1 32154 17204 32154 17204 0 _1009_
rlabel metal2 16882 11526 16882 11526 0 _1010_
rlabel metal2 15778 13022 15778 13022 0 _1011_
rlabel metal2 15226 11288 15226 11288 0 _1012_
rlabel metal1 15226 10608 15226 10608 0 _1013_
rlabel metal1 15732 12818 15732 12818 0 _1014_
rlabel metal2 18078 9146 18078 9146 0 _1015_
rlabel metal2 14904 12580 14904 12580 0 _1016_
rlabel metal2 14490 8908 14490 8908 0 _1017_
rlabel metal1 19054 31314 19054 31314 0 _1018_
rlabel metal2 16790 29036 16790 29036 0 _1019_
rlabel metal2 17342 30464 17342 30464 0 _1020_
rlabel metal1 16698 30770 16698 30770 0 _1021_
rlabel metal1 16330 28492 16330 28492 0 _1022_
rlabel metal2 15778 28934 15778 28934 0 _1023_
rlabel metal4 13892 25568 13892 25568 0 _1024_
rlabel metal1 14490 18666 14490 18666 0 _1025_
rlabel metal2 17710 18156 17710 18156 0 _1026_
rlabel metal1 19734 14314 19734 14314 0 _1027_
rlabel metal2 14766 13872 14766 13872 0 _1028_
rlabel metal2 17158 13702 17158 13702 0 _1029_
rlabel metal1 15364 13362 15364 13362 0 _1030_
rlabel metal2 20654 17408 20654 17408 0 _1031_
rlabel metal1 14398 15878 14398 15878 0 _1032_
rlabel metal1 14076 13158 14076 13158 0 _1033_
rlabel via1 13294 14365 13294 14365 0 _1034_
rlabel metal1 11178 16762 11178 16762 0 _1035_
rlabel metal1 17296 13906 17296 13906 0 _1036_
rlabel metal1 14950 17646 14950 17646 0 _1037_
rlabel metal1 15364 10030 15364 10030 0 _1038_
rlabel metal1 22402 10132 22402 10132 0 _1039_
rlabel metal2 21114 17884 21114 17884 0 _1040_
rlabel metal1 18308 17578 18308 17578 0 _1041_
rlabel metal1 15226 10064 15226 10064 0 _1042_
rlabel metal1 12604 13906 12604 13906 0 _1043_
rlabel metal1 17296 13702 17296 13702 0 _1044_
rlabel metal1 15134 10234 15134 10234 0 _1045_
rlabel metal1 13892 10778 13892 10778 0 _1046_
rlabel metal1 11500 11322 11500 11322 0 _1047_
rlabel metal1 10672 11866 10672 11866 0 _1048_
rlabel metal1 18814 32266 18814 32266 0 _1049_
rlabel metal1 17986 30906 17986 30906 0 _1050_
rlabel metal2 20010 32572 20010 32572 0 _1051_
rlabel metal1 17802 32436 17802 32436 0 _1052_
rlabel metal2 17710 32164 17710 32164 0 _1053_
rlabel metal1 15962 17680 15962 17680 0 _1054_
rlabel metal1 14076 17850 14076 17850 0 _1055_
rlabel metal1 16054 18122 16054 18122 0 _1056_
rlabel metal1 16652 31790 16652 31790 0 _1057_
rlabel metal1 14398 19278 14398 19278 0 _1058_
rlabel metal1 18216 7174 18216 7174 0 _1059_
rlabel metal2 12926 10472 12926 10472 0 _1060_
rlabel metal1 12650 13498 12650 13498 0 _1061_
rlabel metal1 17434 11050 17434 11050 0 _1062_
rlabel metal1 14490 12750 14490 12750 0 _1063_
rlabel metal1 13248 13294 13248 13294 0 _1064_
rlabel metal1 14490 12886 14490 12886 0 _1065_
rlabel metal2 14306 13090 14306 13090 0 _1066_
rlabel metal1 12696 13158 12696 13158 0 _1067_
rlabel metal3 15479 21556 15479 21556 0 _1068_
rlabel metal2 15502 32062 15502 32062 0 _1069_
rlabel metal2 12650 16065 12650 16065 0 _1070_
rlabel metal1 9200 13906 9200 13906 0 _1071_
rlabel metal1 4554 11866 4554 11866 0 _1072_
rlabel metal2 18170 9248 18170 9248 0 _1073_
rlabel metal2 17618 9129 17618 9129 0 _1074_
rlabel via2 17158 16235 17158 16235 0 _1075_
rlabel metal1 16146 27574 16146 27574 0 _1076_
rlabel metal2 13386 26588 13386 26588 0 _1077_
rlabel metal1 25944 9418 25944 9418 0 _1078_
rlabel metal2 20562 8704 20562 8704 0 _1079_
rlabel metal1 20470 8908 20470 8908 0 _1080_
rlabel metal2 20838 10336 20838 10336 0 _1081_
rlabel metal2 20746 11084 20746 11084 0 _1082_
rlabel metal1 19274 10574 19274 10574 0 _1083_
rlabel metal1 19412 19346 19412 19346 0 _1084_
rlabel metal1 18676 19482 18676 19482 0 _1085_
rlabel metal1 20010 10506 20010 10506 0 _1086_
rlabel metal2 20286 9724 20286 9724 0 _1087_
rlabel metal3 19435 15164 19435 15164 0 _1088_
rlabel metal1 15502 19380 15502 19380 0 _1089_
rlabel metal1 15686 19346 15686 19346 0 _1090_
rlabel metal1 5934 19924 5934 19924 0 _1091_
rlabel metal1 8786 18598 8786 18598 0 _1092_
rlabel metal1 17986 24752 17986 24752 0 _1093_
rlabel metal1 17526 24378 17526 24378 0 _1094_
rlabel metal1 16192 24242 16192 24242 0 _1095_
rlabel metal2 14490 24820 14490 24820 0 _1096_
rlabel metal1 17434 24752 17434 24752 0 _1097_
rlabel metal1 15824 25262 15824 25262 0 _1098_
rlabel metal1 18308 25466 18308 25466 0 _1099_
rlabel metal1 18446 25806 18446 25806 0 _1100_
rlabel metal1 21252 25942 21252 25942 0 _1101_
rlabel metal3 16836 18156 16836 18156 0 _1102_
rlabel metal1 21160 18122 21160 18122 0 _1103_
rlabel metal2 20010 25874 20010 25874 0 _1104_
rlabel metal1 17158 25942 17158 25942 0 _1105_
rlabel metal2 15226 25262 15226 25262 0 _1106_
rlabel metal2 17250 27982 17250 27982 0 _1107_
rlabel metal1 14214 6834 14214 6834 0 _1108_
rlabel metal2 16698 7956 16698 7956 0 _1109_
rlabel metal1 16606 8262 16606 8262 0 _1110_
rlabel metal1 16836 11526 16836 11526 0 _1111_
rlabel metal2 19182 6222 19182 6222 0 _1112_
rlabel metal2 18170 8024 18170 8024 0 _1113_
rlabel metal1 15594 19686 15594 19686 0 _1114_
rlabel metal2 16054 26622 16054 26622 0 _1115_
rlabel metal1 16652 25806 16652 25806 0 _1116_
rlabel metal1 14306 26316 14306 26316 0 _1117_
rlabel metal2 16054 25704 16054 25704 0 _1118_
rlabel metal1 14950 25840 14950 25840 0 _1119_
rlabel metal2 9614 25500 9614 25500 0 _1120_
rlabel metal1 14996 25330 14996 25330 0 _1121_
rlabel metal1 9154 24820 9154 24820 0 _1122_
rlabel metal1 14490 19346 14490 19346 0 _1123_
rlabel metal1 16836 5882 16836 5882 0 _1124_
rlabel metal1 15824 14042 15824 14042 0 _1125_
rlabel metal1 13110 15878 13110 15878 0 _1126_
rlabel metal2 11178 25092 11178 25092 0 _1127_
rlabel metal1 7360 26554 7360 26554 0 _1128_
rlabel metal1 8786 23664 8786 23664 0 _1129_
rlabel metal2 9430 25313 9430 25313 0 _1130_
rlabel metal2 13662 25092 13662 25092 0 _1131_
rlabel metal1 9565 24174 9565 24174 0 _1132_
rlabel metal2 9062 24684 9062 24684 0 _1133_
rlabel metal1 12926 23834 12926 23834 0 _1134_
rlabel metal2 12374 24106 12374 24106 0 _1135_
rlabel metal2 6118 26690 6118 26690 0 _1136_
rlabel metal2 9522 28458 9522 28458 0 _1137_
rlabel metal1 13984 19414 13984 19414 0 _1138_
rlabel metal1 14674 28662 14674 28662 0 _1139_
rlabel metal1 17020 20026 17020 20026 0 _1140_
rlabel metal1 15226 28458 15226 28458 0 _1141_
rlabel metal1 13570 27540 13570 27540 0 _1142_
rlabel metal1 5978 27438 5978 27438 0 _1143_
rlabel metal2 9246 28594 9246 28594 0 _1144_
rlabel metal1 12834 16592 12834 16592 0 _1145_
rlabel metal2 12834 16966 12834 16966 0 _1146_
rlabel metal2 12650 17476 12650 17476 0 _1147_
rlabel metal2 12466 17748 12466 17748 0 _1148_
rlabel metal1 20700 7718 20700 7718 0 _1149_
rlabel metal1 20056 8602 20056 8602 0 _1150_
rlabel metal1 19320 4998 19320 4998 0 _1151_
rlabel metal2 18538 4998 18538 4998 0 _1152_
rlabel metal1 20010 12614 20010 12614 0 _1153_
rlabel metal2 20470 16762 20470 16762 0 _1154_
rlabel metal1 20562 13294 20562 13294 0 _1155_
rlabel metal1 20056 12818 20056 12818 0 _1156_
rlabel metal1 19458 12954 19458 12954 0 _1157_
rlabel metal1 13570 18666 13570 18666 0 _1158_
rlabel metal1 13018 18870 13018 18870 0 _1159_
rlabel metal1 10948 18190 10948 18190 0 _1160_
rlabel via2 23322 19261 23322 19261 0 _1161_
rlabel metal1 22770 19380 22770 19380 0 _1162_
rlabel metal1 24518 19312 24518 19312 0 _1163_
rlabel metal1 24380 18938 24380 18938 0 _1164_
rlabel metal1 23598 19346 23598 19346 0 _1165_
rlabel metal2 20010 19720 20010 19720 0 _1166_
rlabel metal1 17296 11730 17296 11730 0 _1167_
rlabel metal2 21482 11679 21482 11679 0 _1168_
rlabel metal1 13662 17102 13662 17102 0 _1169_
rlabel via1 12208 17646 12208 17646 0 _1170_
rlabel metal1 11316 17850 11316 17850 0 _1171_
rlabel metal2 12834 18564 12834 18564 0 _1172_
rlabel metal1 22034 32470 22034 32470 0 _1173_
rlabel metal1 22816 32198 22816 32198 0 _1174_
rlabel metal3 19757 19108 19757 19108 0 _1175_
rlabel metal1 22172 18870 22172 18870 0 _1176_
rlabel metal1 17618 18734 17618 18734 0 _1177_
rlabel metal1 13478 18292 13478 18292 0 _1178_
rlabel metal1 12420 18666 12420 18666 0 _1179_
rlabel metal1 10626 18360 10626 18360 0 _1180_
rlabel metal2 13110 18564 13110 18564 0 _1181_
rlabel metal2 12558 16966 12558 16966 0 _1182_
rlabel metal1 5704 19278 5704 19278 0 _1183_
rlabel metal1 10442 17068 10442 17068 0 _1184_
rlabel metal2 11086 20468 11086 20468 0 _1185_
rlabel metal1 6762 18326 6762 18326 0 _1186_
rlabel metal1 8970 16490 8970 16490 0 _1187_
rlabel metal2 8418 18156 8418 18156 0 _1188_
rlabel metal2 5658 16082 5658 16082 0 _1189_
rlabel metal1 8142 15674 8142 15674 0 _1190_
rlabel metal2 8694 18700 8694 18700 0 _1191_
rlabel metal1 8372 18394 8372 18394 0 _1192_
rlabel metal1 8648 30158 8648 30158 0 _1193_
rlabel metal1 24702 12410 24702 12410 0 _1194_
rlabel metal1 20102 21964 20102 21964 0 _1195_
rlabel metal1 23736 13770 23736 13770 0 _1196_
rlabel metal1 23414 15130 23414 15130 0 _1197_
rlabel metal1 23000 20434 23000 20434 0 _1198_
rlabel metal1 24472 18394 24472 18394 0 _1199_
rlabel metal1 23966 20978 23966 20978 0 _1200_
rlabel metal1 23690 23086 23690 23086 0 _1201_
rlabel metal1 23920 22406 23920 22406 0 _1202_
rlabel metal1 24242 16762 24242 16762 0 _1203_
rlabel metal2 23690 21114 23690 21114 0 _1204_
rlabel metal2 24518 19346 24518 19346 0 _1205_
rlabel metal1 24518 20570 24518 20570 0 _1206_
rlabel metal1 24610 20842 24610 20842 0 _1207_
rlabel metal1 23414 20978 23414 20978 0 _1208_
rlabel metal1 23598 18598 23598 18598 0 _1209_
rlabel metal2 23138 19890 23138 19890 0 _1210_
rlabel metal2 19918 21522 19918 21522 0 _1211_
rlabel metal1 19734 21862 19734 21862 0 _1212_
rlabel metal1 19596 15538 19596 15538 0 _1213_
rlabel metal1 19550 15436 19550 15436 0 _1214_
rlabel metal2 16606 28730 16606 28730 0 _1215_
rlabel metal2 16882 25874 16882 25874 0 _1216_
rlabel metal1 17388 23290 17388 23290 0 _1217_
rlabel metal1 16238 28050 16238 28050 0 _1218_
rlabel metal1 18170 23154 18170 23154 0 _1219_
rlabel metal1 21482 23596 21482 23596 0 _1220_
rlabel metal2 20654 23970 20654 23970 0 _1221_
rlabel metal1 21068 24378 21068 24378 0 _1222_
rlabel metal1 21068 29138 21068 29138 0 _1223_
rlabel metal1 19826 24276 19826 24276 0 _1224_
rlabel metal1 21436 28186 21436 28186 0 _1225_
rlabel metal1 20746 28084 20746 28084 0 _1226_
rlabel metal1 13386 28016 13386 28016 0 _1227_
rlabel metal1 13064 28526 13064 28526 0 _1228_
rlabel metal1 14306 28050 14306 28050 0 _1229_
rlabel via2 22954 10693 22954 10693 0 _1230_
rlabel metal1 15410 21998 15410 21998 0 _1231_
rlabel metal1 17388 21658 17388 21658 0 _1232_
rlabel metal1 16146 21590 16146 21590 0 _1233_
rlabel metal2 13202 28628 13202 28628 0 _1234_
rlabel metal1 8648 28526 8648 28526 0 _1235_
rlabel metal2 9154 27914 9154 27914 0 _1236_
rlabel metal1 7958 20502 7958 20502 0 _1237_
rlabel metal1 7636 14790 7636 14790 0 _1238_
rlabel metal1 7268 9622 7268 9622 0 _1239_
rlabel metal1 13708 7990 13708 7990 0 _1240_
rlabel metal1 13248 21114 13248 21114 0 _1241_
rlabel metal1 13018 20808 13018 20808 0 _1242_
rlabel metal1 15456 14790 15456 14790 0 _1243_
rlabel metal2 14306 11084 14306 11084 0 _1244_
rlabel metal2 6854 14688 6854 14688 0 _1245_
rlabel metal1 7222 14518 7222 14518 0 _1246_
rlabel metal1 13432 13838 13432 13838 0 _1247_
rlabel metal2 14122 7990 14122 7990 0 _1248_
rlabel metal1 13616 9418 13616 9418 0 _1249_
rlabel metal1 15548 13974 15548 13974 0 _1250_
rlabel metal2 13938 14212 13938 14212 0 _1251_
rlabel metal1 12328 14382 12328 14382 0 _1252_
rlabel metal1 10672 14450 10672 14450 0 _1253_
rlabel via2 8694 14467 8694 14467 0 _1254_
rlabel metal1 10074 5814 10074 5814 0 _1255_
rlabel metal1 10580 14246 10580 14246 0 _1256_
rlabel metal2 8326 14144 8326 14144 0 _1257_
rlabel metal1 15318 22066 15318 22066 0 _1258_
rlabel metal1 14398 22610 14398 22610 0 _1259_
rlabel metal1 19366 32538 19366 32538 0 _1260_
rlabel metal1 19780 32266 19780 32266 0 _1261_
rlabel metal1 20010 21454 20010 21454 0 _1262_
rlabel metal2 15410 6630 15410 6630 0 _1263_
rlabel metal1 19780 21318 19780 21318 0 _1264_
rlabel metal1 18906 21624 18906 21624 0 _1265_
rlabel metal1 19872 21658 19872 21658 0 _1266_
rlabel metal1 18630 23732 18630 23732 0 _1267_
rlabel metal1 14674 22678 14674 22678 0 _1268_
rlabel metal1 19274 23698 19274 23698 0 _1269_
rlabel metal2 14674 22559 14674 22559 0 _1270_
rlabel metal1 12006 23494 12006 23494 0 _1271_
rlabel metal2 12558 21896 12558 21896 0 _1272_
rlabel metal1 20332 15062 20332 15062 0 _1273_
rlabel metal1 19872 15674 19872 15674 0 _1274_
rlabel metal1 14260 21998 14260 21998 0 _1275_
rlabel metal1 12788 22678 12788 22678 0 _1276_
rlabel metal1 5336 22610 5336 22610 0 _1277_
rlabel metal1 13294 23052 13294 23052 0 _1278_
rlabel metal1 12834 21998 12834 21998 0 _1279_
rlabel via1 9064 22610 9064 22610 0 _1280_
rlabel metal1 8878 23120 8878 23120 0 _1281_
rlabel metal1 8648 21522 8648 21522 0 _1282_
rlabel metal2 7866 22780 7866 22780 0 _1283_
rlabel metal2 9430 23137 9430 23137 0 _1284_
rlabel metal1 9430 22712 9430 22712 0 _1285_
rlabel metal2 2622 31994 2622 31994 0 _1286_
rlabel metal1 8740 14042 8740 14042 0 _1287_
rlabel metal1 7912 14042 7912 14042 0 _1288_
rlabel metal2 7130 7106 7130 7106 0 _1289_
rlabel metal1 8740 8942 8740 8942 0 _1290_
rlabel metal1 8510 9146 8510 9146 0 _1291_
rlabel metal1 10304 7854 10304 7854 0 _1292_
rlabel metal2 10718 24922 10718 24922 0 _1293_
rlabel metal1 9430 24072 9430 24072 0 _1294_
rlabel metal1 6440 24310 6440 24310 0 _1295_
rlabel metal2 4830 26928 4830 26928 0 _1296_
rlabel metal1 5336 17170 5336 17170 0 _1297_
rlabel metal1 5198 17102 5198 17102 0 _1298_
rlabel metal1 5014 17204 5014 17204 0 _1299_
rlabel metal1 4738 17034 4738 17034 0 _1300_
rlabel metal2 12466 28747 12466 28747 0 _1301_
rlabel metal1 4554 27438 4554 27438 0 _1302_
rlabel metal1 2438 20978 2438 20978 0 _1303_
rlabel metal1 6072 14790 6072 14790 0 _1304_
rlabel metal1 5612 22202 5612 22202 0 _1305_
rlabel metal1 5980 32878 5980 32878 0 _1306_
rlabel metal2 2070 19142 2070 19142 0 _1307_
rlabel metal1 7498 13804 7498 13804 0 _1308_
rlabel metal1 6900 13906 6900 13906 0 _1309_
rlabel metal2 6578 14348 6578 14348 0 _1310_
rlabel metal1 6348 13838 6348 13838 0 _1311_
rlabel metal2 6394 6494 6394 6494 0 _1312_
rlabel via1 7129 8942 7129 8942 0 _1313_
rlabel metal2 6394 9350 6394 9350 0 _1314_
rlabel metal2 9154 17884 9154 17884 0 _1315_
rlabel metal1 9154 17782 9154 17782 0 _1316_
rlabel metal1 6762 16422 6762 16422 0 _1317_
rlabel via2 7774 18411 7774 18411 0 _1318_
rlabel metal1 9108 28050 9108 28050 0 _1319_
rlabel metal1 7728 25330 7728 25330 0 _1320_
rlabel metal1 8326 24650 8326 24650 0 _1321_
rlabel metal1 9844 25262 9844 25262 0 _1322_
rlabel metal1 9154 25330 9154 25330 0 _1323_
rlabel metal1 8694 25398 8694 25398 0 _1324_
rlabel metal2 7866 18887 7866 18887 0 _1325_
rlabel metal1 7360 25942 7360 25942 0 _1326_
rlabel metal1 6532 16626 6532 16626 0 _1327_
rlabel metal1 5612 13362 5612 13362 0 _1328_
rlabel metal2 7406 15708 7406 15708 0 _1329_
rlabel metal1 6164 13294 6164 13294 0 _1330_
rlabel metal1 5796 13294 5796 13294 0 _1331_
rlabel metal2 6946 22916 6946 22916 0 _1332_
rlabel metal1 7038 22984 7038 22984 0 _1333_
rlabel metal1 6486 15062 6486 15062 0 _1334_
rlabel metal1 5842 13940 5842 13940 0 _1335_
rlabel via2 19274 19771 19274 19771 0 clk
rlabel metal3 19849 21964 19849 21964 0 clknet_0_clk
rlabel metal1 7774 7412 7774 7412 0 clknet_4_0_0_clk
rlabel via2 33534 9571 33534 9571 0 clknet_4_10_0_clk
rlabel metal1 32062 16694 32062 16694 0 clknet_4_11_0_clk
rlabel metal2 14122 32368 14122 32368 0 clknet_4_12_0_clk
rlabel metal1 16146 36210 16146 36210 0 clknet_4_13_0_clk
rlabel metal1 31510 32946 31510 32946 0 clknet_4_14_0_clk
rlabel metal2 23874 36992 23874 36992 0 clknet_4_15_0_clk
rlabel metal2 1426 11696 1426 11696 0 clknet_4_1_0_clk
rlabel metal1 14168 2482 14168 2482 0 clknet_4_2_0_clk
rlabel metal1 11408 2482 11408 2482 0 clknet_4_3_0_clk
rlabel metal2 1426 17918 1426 17918 0 clknet_4_4_0_clk
rlabel metal1 2622 25738 2622 25738 0 clknet_4_5_0_clk
rlabel metal1 5934 16082 5934 16082 0 clknet_4_6_0_clk
rlabel metal1 6394 35700 6394 35700 0 clknet_4_7_0_clk
rlabel metal1 21850 3060 21850 3060 0 clknet_4_8_0_clk
rlabel metal2 15042 20128 15042 20128 0 clknet_4_9_0_clk
rlabel metal2 36110 21335 36110 21335 0 dataBusIn[0]
rlabel metal2 36110 21913 36110 21913 0 dataBusIn[1]
rlabel metal2 36110 22559 36110 22559 0 dataBusIn[2]
rlabel metal1 29762 37230 29762 37230 0 dataBusIn[3]
rlabel metal1 29072 37230 29072 37230 0 dataBusIn[4]
rlabel metal2 35282 16575 35282 16575 0 dataBusIn[5]
rlabel metal2 36018 24667 36018 24667 0 dataBusIn[6]
rlabel metal2 36110 24021 36110 24021 0 dataBusIn[7]
rlabel metal2 15502 1520 15502 1520 0 dataBusOut[0]
rlabel metal2 14214 1520 14214 1520 0 dataBusOut[1]
rlabel metal1 13846 4488 13846 4488 0 dataBusOut[2]
rlabel metal2 11638 1418 11638 1418 0 dataBusOut[3]
rlabel metal2 12282 959 12282 959 0 dataBusOut[4]
rlabel metal2 9706 1231 9706 1231 0 dataBusOut[5]
rlabel metal2 10350 1690 10350 1690 0 dataBusOut[6]
rlabel metal2 12926 2234 12926 2234 0 dataBusOut[7]
rlabel metal2 20654 1520 20654 1520 0 dataBusSelect
rlabel metal1 1472 30158 1472 30158 0 gpio[0]
rlabel metal2 22218 36856 22218 36856 0 gpio[10]
rlabel metal1 24886 34646 24886 34646 0 gpio[11]
rlabel metal1 21850 36856 21850 36856 0 gpio[12]
rlabel metal2 21942 36652 21942 36652 0 gpio[13]
rlabel metal1 21390 36652 21390 36652 0 gpio[14]
rlabel metal1 24472 35666 24472 35666 0 gpio[15]
rlabel metal2 13570 1588 13570 1588 0 gpio[16]
rlabel metal2 14858 1690 14858 1690 0 gpio[17]
rlabel metal1 20194 3026 20194 3026 0 gpio[18]
rlabel metal2 21850 3196 21850 3196 0 gpio[19]
rlabel metal1 1564 29206 1564 29206 0 gpio[1]
rlabel metal2 15318 4250 15318 4250 0 gpio[20]
rlabel metal3 35420 15844 35420 15844 0 gpio[21]
rlabel metal2 21942 1588 21942 1588 0 gpio[22]
rlabel metal1 8050 2822 8050 2822 0 gpio[23]
rlabel metal2 21298 1792 21298 1792 0 gpio[24]
rlabel via2 1426 27965 1426 27965 0 gpio[2]
rlabel metal1 1472 28594 1472 28594 0 gpio[3]
rlabel metal2 3174 30260 3174 30260 0 gpio[4]
rlabel metal2 2438 31705 2438 31705 0 gpio[5]
rlabel metal1 1794 31382 1794 31382 0 gpio[6]
rlabel metal1 1426 32470 1426 32470 0 gpio[7]
rlabel metal2 21666 35088 21666 35088 0 gpio[8]
rlabel metal1 22586 36006 22586 36006 0 gpio[9]
rlabel metal1 36202 21658 36202 21658 0 net1
rlabel metal1 14076 2414 14076 2414 0 net10
rlabel metal1 35374 8942 35374 8942 0 net100
rlabel metal1 27968 11186 27968 11186 0 net101
rlabel metal1 33166 6732 33166 6732 0 net102
rlabel metal1 34822 11322 34822 11322 0 net103
rlabel metal1 23460 29002 23460 29002 0 net104
rlabel metal1 18676 15606 18676 15606 0 net105
rlabel metal1 15318 7786 15318 7786 0 net106
rlabel metal2 21390 14450 21390 14450 0 net107
rlabel metal2 17434 12988 17434 12988 0 net108
rlabel metal1 21574 5202 21574 5202 0 net109
rlabel metal2 13662 2587 13662 2587 0 net11
rlabel metal1 17894 25296 17894 25296 0 net110
rlabel metal1 20148 19278 20148 19278 0 net111
rlabel metal1 15732 7514 15732 7514 0 net112
rlabel metal1 17250 19856 17250 19856 0 net113
rlabel metal2 19366 14943 19366 14943 0 net114
rlabel metal1 13340 9690 13340 9690 0 net115
rlabel metal2 14674 6800 14674 6800 0 net116
rlabel metal1 20930 10676 20930 10676 0 net117
rlabel metal2 17986 17408 17986 17408 0 net118
rlabel metal1 17664 17238 17664 17238 0 net119
rlabel metal1 10764 2618 10764 2618 0 net12
rlabel metal1 14582 18734 14582 18734 0 net120
rlabel via1 21942 32402 21942 32402 0 net121
rlabel metal1 21390 30226 21390 30226 0 net122
rlabel metal2 17756 31892 17756 31892 0 net123
rlabel metal1 21344 24106 21344 24106 0 net124
rlabel metal2 21574 18445 21574 18445 0 net125
rlabel metal1 19780 32878 19780 32878 0 net126
rlabel metal1 10534 2414 10534 2414 0 net127
rlabel metal2 12558 2414 12558 2414 0 net128
rlabel metal1 19918 3128 19918 3128 0 net129
rlabel metal1 8786 2346 8786 2346 0 net13
rlabel metal2 9798 17714 9798 17714 0 net130
rlabel metal2 9706 17000 9706 17000 0 net131
rlabel metal2 18630 4063 18630 4063 0 net132
rlabel metal1 33587 16490 33587 16490 0 net133
rlabel metal1 2951 21590 2951 21590 0 net134
rlabel metal1 2744 28118 2744 28118 0 net135
rlabel metal1 17204 21114 17204 21114 0 net136
rlabel metal1 10449 32470 10449 32470 0 net137
rlabel metal1 16376 36006 16376 36006 0 net138
rlabel metal1 21673 36142 21673 36142 0 net139
rlabel metal1 8556 2414 8556 2414 0 net14
rlabel metal1 26135 33558 26135 33558 0 net140
rlabel metal1 22816 34646 22816 34646 0 net141
rlabel metal1 32752 33830 32752 33830 0 net142
rlabel metal1 32660 33966 32660 33966 0 net143
rlabel via2 17066 20893 17066 20893 0 net144
rlabel via1 13569 23698 13569 23698 0 net145
rlabel metal2 33810 28832 33810 28832 0 net146
rlabel metal2 21206 26639 21206 26639 0 net147
rlabel metal1 18032 2482 18032 2482 0 net148
rlabel metal1 14214 3706 14214 3706 0 net149
rlabel metal2 8142 5576 8142 5576 0 net15
rlabel metal1 27416 34578 27416 34578 0 net150
rlabel metal1 15640 20502 15640 20502 0 net151
rlabel metal1 14398 4624 14398 4624 0 net152
rlabel metal2 17342 3740 17342 3740 0 net153
rlabel metal1 13294 4692 13294 4692 0 net154
rlabel metal1 17710 3162 17710 3162 0 net155
rlabel metal2 18078 4318 18078 4318 0 net156
rlabel metal2 17526 3162 17526 3162 0 net157
rlabel metal1 2668 18258 2668 18258 0 net158
rlabel metal2 2346 16762 2346 16762 0 net159
rlabel metal1 8096 4590 8096 4590 0 net16
rlabel metal1 11086 19346 11086 19346 0 net160
rlabel metal1 6992 17306 6992 17306 0 net161
rlabel metal2 7590 15946 7590 15946 0 net162
rlabel metal1 2668 19346 2668 19346 0 net163
rlabel metal1 7406 18666 7406 18666 0 net164
rlabel metal2 3634 16320 3634 16320 0 net165
rlabel metal1 9982 18394 9982 18394 0 net166
rlabel metal1 6716 16490 6716 16490 0 net167
rlabel metal1 10258 5678 10258 5678 0 net168
rlabel metal1 24334 2550 24334 2550 0 net169
rlabel metal1 12880 2618 12880 2618 0 net17
rlabel metal2 9338 15878 9338 15878 0 net170
rlabel metal1 4416 15402 4416 15402 0 net171
rlabel metal1 11224 15402 11224 15402 0 net172
rlabel metal1 5152 16218 5152 16218 0 net173
rlabel metal1 10810 4012 10810 4012 0 net174
rlabel metal2 23414 32674 23414 32674 0 net175
rlabel metal1 12282 3094 12282 3094 0 net176
rlabel metal2 9982 4386 9982 4386 0 net177
rlabel metal2 14582 4556 14582 4556 0 net178
rlabel metal2 8326 3740 8326 3740 0 net179
rlabel metal1 20654 2822 20654 2822 0 net18
rlabel metal1 4416 14314 4416 14314 0 net180
rlabel metal2 16146 4318 16146 4318 0 net181
rlabel metal1 3864 13906 3864 13906 0 net182
rlabel metal1 11132 4658 11132 4658 0 net183
rlabel metal2 13110 20706 13110 20706 0 net184
rlabel metal2 8970 2924 8970 2924 0 net185
rlabel metal1 23690 27336 23690 27336 0 net186
rlabel metal2 25714 31994 25714 31994 0 net187
rlabel metal1 6900 21998 6900 21998 0 net188
rlabel metal1 4554 22202 4554 22202 0 net189
rlabel metal1 7774 32878 7774 32878 0 net19
rlabel metal1 10396 20842 10396 20842 0 net190
rlabel metal2 23506 33184 23506 33184 0 net191
rlabel metal2 2806 21114 2806 21114 0 net192
rlabel metal1 9844 20570 9844 20570 0 net193
rlabel metal1 7958 20570 7958 20570 0 net194
rlabel metal2 10350 22848 10350 22848 0 net195
rlabel metal2 4738 23120 4738 23120 0 net196
rlabel metal1 10534 13260 10534 13260 0 net197
rlabel metal1 3726 21930 3726 21930 0 net198
rlabel metal2 28566 33354 28566 33354 0 net199
rlabel metal1 13708 31722 13708 31722 0 net2
rlabel metal2 18262 33524 18262 33524 0 net20
rlabel metal1 18078 26996 18078 26996 0 net200
rlabel metal2 25438 33796 25438 33796 0 net201
rlabel metal2 5290 25500 5290 25500 0 net202
rlabel metal2 5290 24412 5290 24412 0 net203
rlabel metal1 32706 32946 32706 32946 0 net21
rlabel metal1 7176 33490 7176 33490 0 net22
rlabel metal1 10350 34000 10350 34000 0 net23
rlabel metal2 7682 33456 7682 33456 0 net24
rlabel metal1 12190 33422 12190 33422 0 net25
rlabel metal1 16330 36788 16330 36788 0 net26
rlabel metal1 8924 12954 8924 12954 0 net27
rlabel metal1 29164 25874 29164 25874 0 net28
rlabel metal1 7176 26962 7176 26962 0 net29
rlabel metal1 12972 21590 12972 21590 0 net3
rlabel metal2 9614 26894 9614 26894 0 net30
rlabel metal1 4554 11662 4554 11662 0 net31
rlabel metal2 10626 13022 10626 13022 0 net32
rlabel via1 28185 20842 28185 20842 0 net33
rlabel metal1 31602 15912 31602 15912 0 net34
rlabel metal1 32798 14994 32798 14994 0 net35
rlabel metal2 31878 17731 31878 17731 0 net36
rlabel metal1 29716 17646 29716 17646 0 net37
rlabel metal1 26220 26554 26220 26554 0 net38
rlabel metal1 27692 32878 27692 32878 0 net39
rlabel metal2 13478 29444 13478 29444 0 net4
rlabel viali 33536 30226 33536 30226 0 net40
rlabel metal1 24150 32878 24150 32878 0 net41
rlabel via2 28198 32453 28198 32453 0 net42
rlabel metal1 12466 28084 12466 28084 0 net43
rlabel metal1 8878 34034 8878 34034 0 net44
rlabel metal1 18124 33422 18124 33422 0 net45
rlabel metal1 12604 19346 12604 19346 0 net46
rlabel metal1 24058 28492 24058 28492 0 net47
rlabel metal1 19182 33456 19182 33456 0 net48
rlabel metal2 13248 4658 13248 4658 0 net49
rlabel metal2 29302 35020 29302 35020 0 net5
rlabel metal1 15502 20910 15502 20910 0 net50
rlabel metal2 21206 27812 21206 27812 0 net51
rlabel metal1 26266 28458 26266 28458 0 net52
rlabel metal2 16790 25738 16790 25738 0 net53
rlabel metal2 14812 12682 14812 12682 0 net54
rlabel metal2 19688 6766 19688 6766 0 net55
rlabel metal1 12926 17646 12926 17646 0 net56
rlabel metal2 20286 15385 20286 15385 0 net57
rlabel metal1 30130 30226 30130 30226 0 net58
rlabel metal1 28566 29172 28566 29172 0 net59
rlabel via2 35006 12155 35006 12155 0 net6
rlabel metal1 19688 19346 19688 19346 0 net60
rlabel metal1 16882 15402 16882 15402 0 net61
rlabel metal1 16698 13294 16698 13294 0 net62
rlabel metal2 14904 16082 14904 16082 0 net63
rlabel metal1 18630 25806 18630 25806 0 net64
rlabel metal1 18814 23698 18814 23698 0 net65
rlabel metal1 17112 17102 17112 17102 0 net66
rlabel metal2 15410 28356 15410 28356 0 net67
rlabel metal1 16146 20264 16146 20264 0 net68
rlabel metal1 18308 14926 18308 14926 0 net69
rlabel metal1 12742 29070 12742 29070 0 net7
rlabel metal1 18354 15572 18354 15572 0 net70
rlabel metal1 18944 12070 18944 12070 0 net71
rlabel metal1 21080 28458 21080 28458 0 net72
rlabel via3 17595 12852 17595 12852 0 net73
rlabel metal2 19366 7684 19366 7684 0 net74
rlabel metal1 25622 22542 25622 22542 0 net75
rlabel metal1 18492 14858 18492 14858 0 net76
rlabel metal2 32154 11118 32154 11118 0 net77
rlabel metal1 20424 28526 20424 28526 0 net78
rlabel metal1 35098 28560 35098 28560 0 net79
rlabel metal1 36064 24378 36064 24378 0 net8
rlabel metal1 28198 11152 28198 11152 0 net80
rlabel metal1 27278 13940 27278 13940 0 net81
rlabel metal1 17572 20502 17572 20502 0 net82
rlabel metal2 32706 27540 32706 27540 0 net83
rlabel metal2 17618 23664 17618 23664 0 net84
rlabel metal1 24334 10438 24334 10438 0 net85
rlabel metal1 17710 13260 17710 13260 0 net86
rlabel metal1 29624 9486 29624 9486 0 net87
rlabel metal1 21068 19822 21068 19822 0 net88
rlabel metal1 30176 7990 30176 7990 0 net89
rlabel metal1 35972 3706 35972 3706 0 net9
rlabel metal1 27554 10098 27554 10098 0 net90
rlabel metal1 33350 6766 33350 6766 0 net91
rlabel metal1 31924 8398 31924 8398 0 net92
rlabel metal2 30130 8160 30130 8160 0 net93
rlabel metal2 27554 10268 27554 10268 0 net94
rlabel metal1 33718 10166 33718 10166 0 net95
rlabel metal1 33718 10064 33718 10064 0 net96
rlabel metal1 28060 10642 28060 10642 0 net97
rlabel metal1 28152 5746 28152 5746 0 net98
rlabel metal1 35512 8806 35512 8806 0 net99
rlabel via2 36110 3485 36110 3485 0 nrst
rlabel metal1 16238 17204 16238 17204 0 top8227.PSRCurrentValue\[0\]
rlabel metal2 12742 5984 12742 5984 0 top8227.PSRCurrentValue\[1\]
rlabel metal1 14168 7854 14168 7854 0 top8227.PSRCurrentValue\[2\]
rlabel via2 9706 8483 9706 8483 0 top8227.PSRCurrentValue\[3\]
rlabel via2 13846 6307 13846 6307 0 top8227.PSRCurrentValue\[6\]
rlabel metal2 13570 5593 13570 5593 0 top8227.PSRCurrentValue\[7\]
rlabel metal1 13110 20026 13110 20026 0 top8227.branchBackward
rlabel metal1 14812 18394 14812 18394 0 top8227.branchForward
rlabel metal1 26358 32266 26358 32266 0 top8227.demux.isAddressing
rlabel via2 15870 4131 15870 4131 0 top8227.demux.nmi
rlabel metal1 20240 26758 20240 26758 0 top8227.demux.reset
rlabel metal1 17342 27574 17342 27574 0 top8227.demux.setInterruptFlag
rlabel metal1 27255 32742 27255 32742 0 top8227.demux.state_machine.currentAddress\[0\]
rlabel metal1 28290 34034 28290 34034 0 top8227.demux.state_machine.currentAddress\[10\]
rlabel metal1 24610 31824 24610 31824 0 top8227.demux.state_machine.currentAddress\[11\]
rlabel metal2 15870 32708 15870 32708 0 top8227.demux.state_machine.currentAddress\[12\]
rlabel metal2 29210 33660 29210 33660 0 top8227.demux.state_machine.currentAddress\[1\]
rlabel metal2 30038 32742 30038 32742 0 top8227.demux.state_machine.currentAddress\[2\]
rlabel metal1 22678 33626 22678 33626 0 top8227.demux.state_machine.currentAddress\[3\]
rlabel metal2 32338 32980 32338 32980 0 top8227.demux.state_machine.currentAddress\[4\]
rlabel metal1 20838 31280 20838 31280 0 top8227.demux.state_machine.currentAddress\[5\]
rlabel metal1 21482 29104 21482 29104 0 top8227.demux.state_machine.currentAddress\[6\]
rlabel metal1 18262 29138 18262 29138 0 top8227.demux.state_machine.currentAddress\[7\]
rlabel metal1 28060 33830 28060 33830 0 top8227.demux.state_machine.currentAddress\[8\]
rlabel metal1 26220 32334 26220 32334 0 top8227.demux.state_machine.currentAddress\[9\]
rlabel metal2 34822 11322 34822 11322 0 top8227.demux.state_machine.currentInstruction\[0\]
rlabel metal1 34454 8398 34454 8398 0 top8227.demux.state_machine.currentInstruction\[1\]
rlabel metal1 35006 9690 35006 9690 0 top8227.demux.state_machine.currentInstruction\[2\]
rlabel metal2 35512 9996 35512 9996 0 top8227.demux.state_machine.currentInstruction\[3\]
rlabel metal1 32338 16218 32338 16218 0 top8227.demux.state_machine.currentInstruction\[4\]
rlabel metal1 33994 16558 33994 16558 0 top8227.demux.state_machine.currentInstruction\[5\]
rlabel metal1 26105 29274 26105 29274 0 top8227.demux.state_machine.timeState\[0\]
rlabel metal1 20424 19414 20424 19414 0 top8227.demux.state_machine.timeState\[1\]
rlabel metal2 24058 4454 24058 4454 0 top8227.demux.state_machine.timeState\[2\]
rlabel metal1 25346 28186 25346 28186 0 top8227.demux.state_machine.timeState\[3\]
rlabel via3 21965 18020 21965 18020 0 top8227.demux.state_machine.timeState\[4\]
rlabel metal1 19734 23766 19734 23766 0 top8227.demux.state_machine.timeState\[5\]
rlabel via2 21022 29597 21022 29597 0 top8227.demux.state_machine.timeState\[6\]
rlabel metal2 15962 20706 15962 20706 0 top8227.freeCarry
rlabel metal1 15594 2482 15594 2482 0 top8227.instructionLoader.interruptInjector.interruptRequest
rlabel metal1 18354 4080 18354 4080 0 top8227.instructionLoader.interruptInjector.irqGenerated
rlabel metal1 18722 2618 18722 2618 0 top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
rlabel metal2 16514 2329 16514 2329 0 top8227.instructionLoader.interruptInjector.irqSync.nextQ2
rlabel metal2 14306 3774 14306 3774 0 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
rlabel metal1 15824 4250 15824 4250 0 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
rlabel metal1 13616 2618 13616 2618 0 top8227.instructionLoader.interruptInjector.nmiSync.in
rlabel metal2 13018 3332 13018 3332 0 top8227.instructionLoader.interruptInjector.nmiSync.nextQ2
rlabel metal2 19550 27370 19550 27370 0 top8227.instructionLoader.interruptInjector.resetDetected
rlabel metal1 9200 17306 9200 17306 0 top8227.internalDataflow.accRegToDB\[0\]
rlabel metal2 11178 23868 11178 23868 0 top8227.internalDataflow.accRegToDB\[1\]
rlabel metal1 3266 20978 3266 20978 0 top8227.internalDataflow.accRegToDB\[2\]
rlabel metal2 3174 24599 3174 24599 0 top8227.internalDataflow.accRegToDB\[3\]
rlabel metal1 3910 25670 3910 25670 0 top8227.internalDataflow.accRegToDB\[4\]
rlabel metal1 6210 24684 6210 24684 0 top8227.internalDataflow.accRegToDB\[5\]
rlabel metal2 2346 21386 2346 21386 0 top8227.internalDataflow.accRegToDB\[6\]
rlabel metal1 12742 26316 12742 26316 0 top8227.internalDataflow.accRegToDB\[7\]
rlabel metal1 14536 34102 14536 34102 0 top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
rlabel metal2 14674 34238 14674 34238 0 top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
rlabel metal1 12880 34714 12880 34714 0 top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
rlabel via2 14214 33507 14214 33507 0 top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
rlabel metal2 14766 35887 14766 35887 0 top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
rlabel metal1 15318 36346 15318 36346 0 top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
rlabel metal1 10672 28730 10672 28730 0 top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
rlabel metal2 13018 26690 13018 26690 0 top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
rlabel metal1 12880 31246 12880 31246 0 top8227.internalDataflow.addressLowBusModule.busInputs\[16\]
rlabel metal1 11730 25296 11730 25296 0 top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
rlabel metal2 8832 21828 8832 21828 0 top8227.internalDataflow.addressLowBusModule.busInputs\[18\]
rlabel metal1 7038 24038 7038 24038 0 top8227.internalDataflow.addressLowBusModule.busInputs\[19\]
rlabel metal1 5750 22644 5750 22644 0 top8227.internalDataflow.addressLowBusModule.busInputs\[20\]
rlabel metal1 7866 34034 7866 34034 0 top8227.internalDataflow.addressLowBusModule.busInputs\[21\]
rlabel metal2 6486 34289 6486 34289 0 top8227.internalDataflow.addressLowBusModule.busInputs\[22\]
rlabel metal1 12972 19278 12972 19278 0 top8227.internalDataflow.addressLowBusModule.busInputs\[23\]
rlabel metal3 11224 17340 11224 17340 0 top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
rlabel metal2 11960 21556 11960 21556 0 top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
rlabel metal1 3174 12308 3174 12308 0 top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
rlabel metal1 3680 17646 3680 17646 0 top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
rlabel metal1 3588 13770 3588 13770 0 top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
rlabel metal4 2668 19108 2668 19108 0 top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
rlabel via2 4646 20893 4646 20893 0 top8227.internalDataflow.addressLowBusModule.busInputs\[30\]
rlabel metal2 8602 15521 8602 15521 0 top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
rlabel metal1 10764 20434 10764 20434 0 top8227.internalDataflow.addressLowBusModule.busInputs\[32\]
rlabel metal1 10810 21488 10810 21488 0 top8227.internalDataflow.addressLowBusModule.busInputs\[33\]
rlabel metal2 5106 22338 5106 22338 0 top8227.internalDataflow.addressLowBusModule.busInputs\[34\]
rlabel metal2 5428 20366 5428 20366 0 top8227.internalDataflow.addressLowBusModule.busInputs\[35\]
rlabel metal1 4002 22066 4002 22066 0 top8227.internalDataflow.addressLowBusModule.busInputs\[36\]
rlabel metal1 7452 21318 7452 21318 0 top8227.internalDataflow.addressLowBusModule.busInputs\[37\]
rlabel metal1 4922 20944 4922 20944 0 top8227.internalDataflow.addressLowBusModule.busInputs\[38\]
rlabel metal1 8878 20978 8878 20978 0 top8227.internalDataflow.addressLowBusModule.busInputs\[39\]
rlabel metal2 11454 8092 11454 8092 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
rlabel metal1 10396 6222 10396 6222 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
rlabel metal1 12834 6970 12834 6970 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
rlabel metal1 10212 9010 10212 9010 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
rlabel metal1 9883 6970 9883 6970 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
rlabel metal1 9706 15538 9706 15538 0 top8227.internalDataflow.stackBusModule.busInputs\[32\]
rlabel metal2 11362 16762 11362 16762 0 top8227.internalDataflow.stackBusModule.busInputs\[33\]
rlabel metal1 5198 15606 5198 15606 0 top8227.internalDataflow.stackBusModule.busInputs\[34\]
rlabel metal1 4186 14518 4186 14518 0 top8227.internalDataflow.stackBusModule.busInputs\[35\]
rlabel metal2 3726 15674 3726 15674 0 top8227.internalDataflow.stackBusModule.busInputs\[36\]
rlabel metal1 6946 16558 6946 16558 0 top8227.internalDataflow.stackBusModule.busInputs\[37\]
rlabel metal1 5750 16014 5750 16014 0 top8227.internalDataflow.stackBusModule.busInputs\[38\]
rlabel metal1 8372 16218 8372 16218 0 top8227.internalDataflow.stackBusModule.busInputs\[39\]
rlabel metal2 10718 19108 10718 19108 0 top8227.internalDataflow.stackBusModule.busInputs\[40\]
rlabel metal1 11638 20026 11638 20026 0 top8227.internalDataflow.stackBusModule.busInputs\[41\]
rlabel metal2 3450 19516 3450 19516 0 top8227.internalDataflow.stackBusModule.busInputs\[42\]
rlabel via1 3542 18938 3542 18938 0 top8227.internalDataflow.stackBusModule.busInputs\[43\]
rlabel metal2 4370 16388 4370 16388 0 top8227.internalDataflow.stackBusModule.busInputs\[44\]
rlabel metal2 7130 18088 7130 18088 0 top8227.internalDataflow.stackBusModule.busInputs\[45\]
rlabel metal1 3128 17306 3128 17306 0 top8227.internalDataflow.stackBusModule.busInputs\[46\]
rlabel metal1 8142 19346 8142 19346 0 top8227.internalDataflow.stackBusModule.busInputs\[47\]
rlabel metal2 15042 4352 15042 4352 0 top8227.negEdgeDetector.q1
rlabel metal1 23506 2482 23506 2482 0 top8227.pulse_slower.currentEnableState\[0\]
rlabel metal1 24058 2482 24058 2482 0 top8227.pulse_slower.currentEnableState\[1\]
rlabel metal1 22034 3536 22034 3536 0 top8227.pulse_slower.nextEnableState\[0\]
rlabel metal1 25024 2618 25024 2618 0 top8227.pulse_slower.nextEnableState\[1\]
<< properties >>
string FIXED_BBOX 0 0 37582 39726
<< end >>

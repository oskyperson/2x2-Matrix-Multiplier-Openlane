VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO calculator_top
  CLASS BLOCK ;
  FOREIGN calculator_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 218.065 BY 228.785 ;
  PIN ColOut[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END ColOut[0]
  PIN ColOut[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END ColOut[1]
  PIN ColOut[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END ColOut[2]
  PIN ColOut[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END ColOut[3]
  PIN RowIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END RowIn[0]
  PIN RowIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END RowIn[1]
  PIN RowIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END RowIn[2]
  PIN RowIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END RowIn[3]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 217.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 212.760 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 212.760 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 217.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 212.760 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 212.760 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END clk
  PIN complete
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END complete
  PIN display_output[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 224.785 103.410 228.785 ;
    END
  END display_output[0]
  PIN display_output[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 149.640 218.065 150.240 ;
    END
  END display_output[10]
  PIN display_output[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 115.640 218.065 116.240 ;
    END
  END display_output[11]
  PIN display_output[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 146.240 218.065 146.840 ;
    END
  END display_output[12]
  PIN display_output[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 125.840 218.065 126.440 ;
    END
  END display_output[13]
  PIN display_output[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 142.840 218.065 143.440 ;
    END
  END display_output[14]
  PIN display_output[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 224.785 100.190 228.785 ;
    END
  END display_output[15]
  PIN display_output[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 224.785 106.630 228.785 ;
    END
  END display_output[1]
  PIN display_output[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 224.785 113.070 228.785 ;
    END
  END display_output[2]
  PIN display_output[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 224.785 119.510 228.785 ;
    END
  END display_output[3]
  PIN display_output[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 122.440 218.065 123.040 ;
    END
  END display_output[4]
  PIN display_output[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 139.440 218.065 140.040 ;
    END
  END display_output[5]
  PIN display_output[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 119.040 218.065 119.640 ;
    END
  END display_output[6]
  PIN display_output[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 136.040 218.065 136.640 ;
    END
  END display_output[7]
  PIN display_output[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 129.240 218.065 129.840 ;
    END
  END display_output[8]
  PIN display_output[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.065 132.640 218.065 133.240 ;
    END
  END display_output[9]
  PIN input_state_FPGA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END input_state_FPGA[0]
  PIN input_state_FPGA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END input_state_FPGA[1]
  PIN input_state_FPGA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END input_state_FPGA[2]
  PIN key_pressed
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END key_pressed
  PIN nRST
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 214.065 27.240 218.065 27.840 ;
    END
  END nRST
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 212.710 217.685 ;
      LAYER li1 ;
        RECT 5.520 10.795 212.520 217.685 ;
      LAYER met1 ;
        RECT 0.530 10.640 212.520 217.840 ;
      LAYER met2 ;
        RECT 0.550 224.505 99.630 225.490 ;
        RECT 100.470 224.505 102.850 225.490 ;
        RECT 103.690 224.505 106.070 225.490 ;
        RECT 106.910 224.505 112.510 225.490 ;
        RECT 113.350 224.505 118.950 225.490 ;
        RECT 119.790 224.505 211.500 225.490 ;
        RECT 0.550 4.280 211.500 224.505 ;
        RECT 0.550 4.000 57.770 4.280 ;
        RECT 58.610 4.000 211.500 4.280 ;
      LAYER met3 ;
        RECT 0.525 211.840 214.065 217.765 ;
        RECT 4.400 210.440 214.065 211.840 ;
        RECT 0.525 150.640 214.065 210.440 ;
        RECT 0.525 149.240 213.665 150.640 ;
        RECT 0.525 147.240 214.065 149.240 ;
        RECT 0.525 145.840 213.665 147.240 ;
        RECT 0.525 143.840 214.065 145.840 ;
        RECT 0.525 142.440 213.665 143.840 ;
        RECT 0.525 140.440 214.065 142.440 ;
        RECT 4.400 139.040 213.665 140.440 ;
        RECT 0.525 137.040 214.065 139.040 ;
        RECT 0.525 135.640 213.665 137.040 ;
        RECT 0.525 133.640 214.065 135.640 ;
        RECT 0.525 132.240 213.665 133.640 ;
        RECT 0.525 130.240 214.065 132.240 ;
        RECT 4.400 128.840 213.665 130.240 ;
        RECT 0.525 126.840 214.065 128.840 ;
        RECT 4.400 125.440 213.665 126.840 ;
        RECT 0.525 123.440 214.065 125.440 ;
        RECT 0.525 122.040 213.665 123.440 ;
        RECT 0.525 120.040 214.065 122.040 ;
        RECT 0.525 118.640 213.665 120.040 ;
        RECT 0.525 116.640 214.065 118.640 ;
        RECT 4.400 115.240 213.665 116.640 ;
        RECT 0.525 113.240 214.065 115.240 ;
        RECT 4.400 111.840 214.065 113.240 ;
        RECT 0.525 89.440 214.065 111.840 ;
        RECT 4.400 88.040 214.065 89.440 ;
        RECT 0.525 86.040 214.065 88.040 ;
        RECT 4.400 84.640 214.065 86.040 ;
        RECT 0.525 79.240 214.065 84.640 ;
        RECT 4.400 77.840 214.065 79.240 ;
        RECT 0.525 75.840 214.065 77.840 ;
        RECT 4.400 74.440 214.065 75.840 ;
        RECT 0.525 65.640 214.065 74.440 ;
        RECT 4.400 64.240 214.065 65.640 ;
        RECT 0.525 62.240 214.065 64.240 ;
        RECT 4.400 60.840 214.065 62.240 ;
        RECT 0.525 58.840 214.065 60.840 ;
        RECT 4.400 57.440 214.065 58.840 ;
        RECT 0.525 28.240 214.065 57.440 ;
        RECT 0.525 26.840 213.665 28.240 ;
        RECT 0.525 10.715 214.065 26.840 ;
      LAYER met4 ;
        RECT 85.855 54.575 174.240 194.305 ;
        RECT 176.640 54.575 177.540 194.305 ;
        RECT 179.940 54.575 201.185 194.305 ;
      LAYER met5 ;
        RECT 114.660 136.900 194.460 138.500 ;
  END
END calculator_top
END LIBRARY

